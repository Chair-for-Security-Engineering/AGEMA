/* modified netlist. Source: module Midori64 in file /Midori_round_based/AGEMA/Midori64.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module Midori64_GHPC_Pipeline_d1 (DataIn_s0, key_s0, clk, reset, enc_dec, key_s1, DataIn_s1, Fresh, DataOut_s0, done, DataOut_s1);
    input [63:0] DataIn_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input enc_dec ;
    input [127:0] key_s1 ;
    input [63:0] DataIn_s1 ;
    input [255:0] Fresh ;
    output [63:0] DataOut_s0 ;
    output done ;
    output [63:0] DataOut_s1 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3024 ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n12 ;
    wire controller_roundCounter_n11 ;
    wire controller_roundCounter_n10 ;
    wire controller_roundCounter_n9 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n7 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n3 ;
    wire controller_roundCounter_n2 ;
    wire controller_roundCounter_n1 ;
    wire controller_roundCounter_N10 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N8 ;
    wire controller_roundCounter_N7 ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_SelectedKey_0_ ;
    wire Midori_rounds_SelectedKey_1_ ;
    wire Midori_rounds_SelectedKey_2_ ;
    wire Midori_rounds_SelectedKey_3_ ;
    wire Midori_rounds_SelectedKey_4_ ;
    wire Midori_rounds_SelectedKey_5_ ;
    wire Midori_rounds_SelectedKey_6_ ;
    wire Midori_rounds_SelectedKey_7_ ;
    wire Midori_rounds_SelectedKey_8_ ;
    wire Midori_rounds_SelectedKey_9_ ;
    wire Midori_rounds_SelectedKey_10_ ;
    wire Midori_rounds_SelectedKey_11_ ;
    wire Midori_rounds_SelectedKey_12_ ;
    wire Midori_rounds_SelectedKey_13_ ;
    wire Midori_rounds_SelectedKey_14_ ;
    wire Midori_rounds_SelectedKey_15_ ;
    wire Midori_rounds_SelectedKey_16_ ;
    wire Midori_rounds_SelectedKey_17_ ;
    wire Midori_rounds_SelectedKey_18_ ;
    wire Midori_rounds_SelectedKey_19_ ;
    wire Midori_rounds_SelectedKey_20_ ;
    wire Midori_rounds_SelectedKey_21_ ;
    wire Midori_rounds_SelectedKey_22_ ;
    wire Midori_rounds_SelectedKey_23_ ;
    wire Midori_rounds_SelectedKey_24_ ;
    wire Midori_rounds_SelectedKey_25_ ;
    wire Midori_rounds_SelectedKey_26_ ;
    wire Midori_rounds_SelectedKey_27_ ;
    wire Midori_rounds_SelectedKey_28_ ;
    wire Midori_rounds_SelectedKey_29_ ;
    wire Midori_rounds_SelectedKey_30_ ;
    wire Midori_rounds_SelectedKey_31_ ;
    wire Midori_rounds_SelectedKey_32_ ;
    wire Midori_rounds_SelectedKey_33_ ;
    wire Midori_rounds_SelectedKey_34_ ;
    wire Midori_rounds_SelectedKey_35_ ;
    wire Midori_rounds_SelectedKey_36_ ;
    wire Midori_rounds_SelectedKey_37_ ;
    wire Midori_rounds_SelectedKey_38_ ;
    wire Midori_rounds_SelectedKey_39_ ;
    wire Midori_rounds_SelectedKey_40_ ;
    wire Midori_rounds_SelectedKey_41_ ;
    wire Midori_rounds_SelectedKey_42_ ;
    wire Midori_rounds_SelectedKey_43_ ;
    wire Midori_rounds_SelectedKey_44_ ;
    wire Midori_rounds_SelectedKey_45_ ;
    wire Midori_rounds_SelectedKey_46_ ;
    wire Midori_rounds_SelectedKey_47_ ;
    wire Midori_rounds_SelectedKey_48_ ;
    wire Midori_rounds_SelectedKey_49_ ;
    wire Midori_rounds_SelectedKey_50_ ;
    wire Midori_rounds_SelectedKey_51_ ;
    wire Midori_rounds_SelectedKey_52_ ;
    wire Midori_rounds_SelectedKey_53_ ;
    wire Midori_rounds_SelectedKey_54_ ;
    wire Midori_rounds_SelectedKey_55_ ;
    wire Midori_rounds_SelectedKey_56_ ;
    wire Midori_rounds_SelectedKey_57_ ;
    wire Midori_rounds_SelectedKey_58_ ;
    wire Midori_rounds_SelectedKey_59_ ;
    wire Midori_rounds_SelectedKey_60_ ;
    wire Midori_rounds_SelectedKey_61_ ;
    wire Midori_rounds_SelectedKey_62_ ;
    wire Midori_rounds_SelectedKey_63_ ;
    wire Midori_rounds_constant_MUX_n217 ;
    wire Midori_rounds_constant_MUX_n216 ;
    wire Midori_rounds_constant_MUX_n215 ;
    wire Midori_rounds_constant_MUX_n214 ;
    wire Midori_rounds_constant_MUX_n213 ;
    wire Midori_rounds_constant_MUX_n212 ;
    wire Midori_rounds_constant_MUX_n211 ;
    wire Midori_rounds_constant_MUX_n210 ;
    wire Midori_rounds_constant_MUX_n209 ;
    wire Midori_rounds_constant_MUX_n208 ;
    wire Midori_rounds_constant_MUX_n207 ;
    wire Midori_rounds_constant_MUX_n206 ;
    wire Midori_rounds_constant_MUX_n205 ;
    wire Midori_rounds_constant_MUX_n204 ;
    wire Midori_rounds_constant_MUX_n203 ;
    wire Midori_rounds_constant_MUX_n202 ;
    wire Midori_rounds_constant_MUX_n201 ;
    wire Midori_rounds_constant_MUX_n200 ;
    wire Midori_rounds_constant_MUX_n199 ;
    wire Midori_rounds_constant_MUX_n198 ;
    wire Midori_rounds_constant_MUX_n197 ;
    wire Midori_rounds_constant_MUX_n196 ;
    wire Midori_rounds_constant_MUX_n195 ;
    wire Midori_rounds_constant_MUX_n194 ;
    wire Midori_rounds_constant_MUX_n193 ;
    wire Midori_rounds_constant_MUX_n192 ;
    wire Midori_rounds_constant_MUX_n191 ;
    wire Midori_rounds_constant_MUX_n190 ;
    wire Midori_rounds_constant_MUX_n189 ;
    wire Midori_rounds_constant_MUX_n188 ;
    wire Midori_rounds_constant_MUX_n187 ;
    wire Midori_rounds_constant_MUX_n186 ;
    wire Midori_rounds_constant_MUX_n185 ;
    wire Midori_rounds_constant_MUX_n184 ;
    wire Midori_rounds_constant_MUX_n183 ;
    wire Midori_rounds_constant_MUX_n182 ;
    wire Midori_rounds_constant_MUX_n181 ;
    wire Midori_rounds_constant_MUX_n180 ;
    wire Midori_rounds_constant_MUX_n179 ;
    wire Midori_rounds_constant_MUX_n178 ;
    wire Midori_rounds_constant_MUX_n177 ;
    wire Midori_rounds_constant_MUX_n176 ;
    wire Midori_rounds_constant_MUX_n175 ;
    wire Midori_rounds_constant_MUX_n174 ;
    wire Midori_rounds_constant_MUX_n173 ;
    wire Midori_rounds_constant_MUX_n172 ;
    wire Midori_rounds_constant_MUX_n171 ;
    wire Midori_rounds_constant_MUX_n170 ;
    wire Midori_rounds_constant_MUX_n169 ;
    wire Midori_rounds_constant_MUX_n168 ;
    wire Midori_rounds_constant_MUX_n167 ;
    wire Midori_rounds_constant_MUX_n166 ;
    wire Midori_rounds_constant_MUX_n165 ;
    wire Midori_rounds_constant_MUX_n164 ;
    wire Midori_rounds_constant_MUX_n163 ;
    wire Midori_rounds_constant_MUX_n162 ;
    wire Midori_rounds_constant_MUX_n161 ;
    wire Midori_rounds_constant_MUX_n160 ;
    wire Midori_rounds_constant_MUX_n159 ;
    wire Midori_rounds_constant_MUX_n158 ;
    wire Midori_rounds_constant_MUX_n157 ;
    wire Midori_rounds_constant_MUX_n156 ;
    wire Midori_rounds_constant_MUX_n155 ;
    wire Midori_rounds_constant_MUX_n154 ;
    wire Midori_rounds_constant_MUX_n153 ;
    wire Midori_rounds_constant_MUX_n152 ;
    wire Midori_rounds_constant_MUX_n151 ;
    wire Midori_rounds_constant_MUX_n150 ;
    wire Midori_rounds_constant_MUX_n149 ;
    wire Midori_rounds_constant_MUX_n148 ;
    wire Midori_rounds_constant_MUX_n147 ;
    wire Midori_rounds_constant_MUX_n146 ;
    wire Midori_rounds_constant_MUX_n145 ;
    wire Midori_rounds_constant_MUX_n144 ;
    wire Midori_rounds_constant_MUX_n143 ;
    wire Midori_rounds_constant_MUX_n142 ;
    wire Midori_rounds_constant_MUX_n141 ;
    wire Midori_rounds_constant_MUX_n140 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n135 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_MUXInst_n11 ;
    wire Midori_rounds_MUXInst_n10 ;
    wire Midori_rounds_MUXInst_n9 ;
    wire Midori_rounds_MUXInst_n8 ;
    wire Midori_rounds_roundResult_Reg_SFF_0_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_1_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_2_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_3_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_4_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_5_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_6_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_7_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_8_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_9_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_10_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_11_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_12_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_13_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_14_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_15_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_16_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_17_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_18_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_19_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_20_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_21_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_22_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_23_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_24_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_25_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_26_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_27_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_28_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_29_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_30_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_31_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_32_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_33_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_34_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_35_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_36_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_37_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_38_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_39_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_40_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_41_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_42_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_43_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_44_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_45_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_46_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_47_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_48_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_49_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_50_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_51_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_52_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_53_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_54_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_55_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_56_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_57_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_58_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_59_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_60_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_61_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_62_DQ ;
    wire Midori_rounds_roundResult_Reg_SFF_63_DQ ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n4 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [15:0] Midori_rounds_round_Constant ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;

    /* cells in depth 0 */
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U64 ( .a ({key_s1[73], key_s0[73]}), .b ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1458, wk[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U63 ( .a ({key_s1[72], key_s0[72]}), .b ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1461, wk[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U62 ( .a ({key_s1[71], key_s0[71]}), .b ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1464, wk[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U61 ( .a ({key_s1[6], key_s0[6]}), .b ({key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1467, wk[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U60 ( .a ({key_s1[127], key_s0[127]}), .b ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1470, wk[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U59 ( .a ({key_s1[126], key_s0[126]}), .b ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1473, wk[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U58 ( .a ({key_s1[125], key_s0[125]}), .b ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1476, wk[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U57 ( .a ({key_s1[124], key_s0[124]}), .b ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1479, wk[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U56 ( .a ({key_s1[5], key_s0[5]}), .b ({key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1482, wk[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U55 ( .a ({key_s1[123], key_s0[123]}), .b ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1485, wk[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U54 ( .a ({key_s1[122], key_s0[122]}), .b ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1488, wk[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U53 ( .a ({key_s1[121], key_s0[121]}), .b ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1491, wk[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U52 ( .a ({key_s1[120], key_s0[120]}), .b ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1494, wk[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U51 ( .a ({key_s1[119], key_s0[119]}), .b ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1497, wk[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U50 ( .a ({key_s1[118], key_s0[118]}), .b ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1500, wk[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U49 ( .a ({key_s1[117], key_s0[117]}), .b ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1503, wk[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U48 ( .a ({key_s1[116], key_s0[116]}), .b ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1506, wk[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U47 ( .a ({key_s1[115], key_s0[115]}), .b ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1509, wk[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U46 ( .a ({key_s1[114], key_s0[114]}), .b ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1512, wk[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U45 ( .a ({key_s1[4], key_s0[4]}), .b ({key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1515, wk[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U44 ( .a ({key_s1[113], key_s0[113]}), .b ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1518, wk[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U43 ( .a ({key_s1[112], key_s0[112]}), .b ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1521, wk[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U42 ( .a ({key_s1[111], key_s0[111]}), .b ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1524, wk[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U41 ( .a ({key_s1[110], key_s0[110]}), .b ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1527, wk[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U40 ( .a ({key_s1[109], key_s0[109]}), .b ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1530, wk[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U39 ( .a ({key_s1[108], key_s0[108]}), .b ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1533, wk[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U38 ( .a ({key_s1[107], key_s0[107]}), .b ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1536, wk[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U37 ( .a ({key_s1[106], key_s0[106]}), .b ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1539, wk[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U36 ( .a ({key_s1[105], key_s0[105]}), .b ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1542, wk[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U35 ( .a ({key_s1[104], key_s0[104]}), .b ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1545, wk[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U34 ( .a ({key_s1[3], key_s0[3]}), .b ({key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1548, wk[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U33 ( .a ({key_s1[103], key_s0[103]}), .b ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1551, wk[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U32 ( .a ({key_s1[102], key_s0[102]}), .b ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1554, wk[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U31 ( .a ({key_s1[101], key_s0[101]}), .b ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1557, wk[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U30 ( .a ({key_s1[100], key_s0[100]}), .b ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1560, wk[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U29 ( .a ({key_s1[35], key_s0[35]}), .b ({key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_1563, wk[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U28 ( .a ({key_s1[34], key_s0[34]}), .b ({key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_1566, wk[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U27 ( .a ({key_s1[33], key_s0[33]}), .b ({key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_1569, wk[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U26 ( .a ({key_s1[32], key_s0[32]}), .b ({key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_1572, wk[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U25 ( .a ({key_s1[31], key_s0[31]}), .b ({key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_1575, wk[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U24 ( .a ({key_s1[30], key_s0[30]}), .b ({key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_1578, wk[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U23 ( .a ({key_s1[2], key_s0[2]}), .b ({key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1581, wk[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U22 ( .a ({key_s1[29], key_s0[29]}), .b ({key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_1584, wk[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U21 ( .a ({key_s1[28], key_s0[28]}), .b ({key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_1587, wk[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U20 ( .a ({key_s1[27], key_s0[27]}), .b ({key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_1590, wk[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U19 ( .a ({key_s1[26], key_s0[26]}), .b ({key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_1593, wk[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U18 ( .a ({key_s1[25], key_s0[25]}), .b ({key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_1596, wk[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U17 ( .a ({key_s1[24], key_s0[24]}), .b ({key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_1599, wk[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U16 ( .a ({key_s1[23], key_s0[23]}), .b ({key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_1602, wk[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U15 ( .a ({key_s1[22], key_s0[22]}), .b ({key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_1605, wk[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U14 ( .a ({key_s1[21], key_s0[21]}), .b ({key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_1608, wk[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U13 ( .a ({key_s1[20], key_s0[20]}), .b ({key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_1611, wk[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U12 ( .a ({key_s1[1], key_s0[1]}), .b ({key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1614, wk[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U11 ( .a ({key_s1[19], key_s0[19]}), .b ({key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_1617, wk[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U10 ( .a ({key_s1[18], key_s0[18]}), .b ({key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_1620, wk[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U9 ( .a ({key_s1[17], key_s0[17]}), .b ({key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_1623, wk[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U8 ( .a ({key_s1[16], key_s0[16]}), .b ({key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_1626, wk[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U7 ( .a ({key_s1[15], key_s0[15]}), .b ({key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_1629, wk[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U6 ( .a ({key_s1[14], key_s0[14]}), .b ({key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_1632, wk[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U5 ( .a ({key_s1[13], key_s0[13]}), .b ({key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_1635, wk[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U4 ( .a ({key_s1[12], key_s0[12]}), .b ({key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_1638, wk[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U3 ( .a ({key_s1[11], key_s0[11]}), .b ({key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_1641, wk[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U2 ( .a ({key_s1[10], key_s0[10]}), .b ({key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_1644, wk[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) keys_U1 ( .a ({key_s1[0], key_s0[0]}), .b ({key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_1647, wk[0]}) ) ;
    NOR2_X1 controller_U3 ( .A1 (controller_n2), .A2 (controller_n1), .ZN (new_AGEMA_signal_3024) ) ;
    NAND2_X1 controller_U2 ( .A1 (round_Signal[0]), .A2 (round_Signal[1]), .ZN (controller_n1) ) ;
    NAND2_X1 controller_U1 ( .A1 (round_Signal[2]), .A2 (round_Signal[3]), .ZN (controller_n2) ) ;
    INV_X1 controller_roundCounter_U14 ( .A (controller_roundCounter_n13), .ZN (controller_roundCounter_n2) ) ;
    MUX2_X1 controller_roundCounter_U13 ( .S (controller_roundCounter_n6), .A (controller_roundCounter_n12), .B (controller_roundCounter_n11), .Z (controller_roundCounter_n13) ) ;
    NOR2_X1 controller_roundCounter_U12 ( .A1 (reset), .A2 (controller_roundCounter_n10), .ZN (controller_roundCounter_N8) ) ;
    XNOR2_X1 controller_roundCounter_U11 ( .A (round_Signal[0]), .B (round_Signal[1]), .ZN (controller_roundCounter_n10) ) ;
    MUX2_X1 controller_roundCounter_U10 ( .S (round_Signal[3]), .A (controller_roundCounter_n9), .B (controller_roundCounter_n8), .Z (controller_roundCounter_N10) ) ;
    NAND2_X1 controller_roundCounter_U9 ( .A1 (controller_roundCounter_n12), .A2 (controller_roundCounter_n7), .ZN (controller_roundCounter_n8) ) ;
    NAND2_X1 controller_roundCounter_U8 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n3), .ZN (controller_roundCounter_n7) ) ;
    NOR2_X1 controller_roundCounter_U7 ( .A1 (controller_roundCounter_n5), .A2 (controller_roundCounter_N7), .ZN (controller_roundCounter_n12) ) ;
    NOR2_X1 controller_roundCounter_U6 ( .A1 (round_Signal[1]), .A2 (reset), .ZN (controller_roundCounter_n5) ) ;
    NOR2_X1 controller_roundCounter_U5 ( .A1 (controller_roundCounter_n6), .A2 (controller_roundCounter_n11), .ZN (controller_roundCounter_n9) ) ;
    NAND2_X1 controller_roundCounter_U4 ( .A1 (round_Signal[1]), .A2 (controller_roundCounter_n4), .ZN (controller_roundCounter_n11) ) ;
    NOR2_X1 controller_roundCounter_U3 ( .A1 (reset), .A2 (controller_roundCounter_n1), .ZN (controller_roundCounter_n4) ) ;
    NOR2_X1 controller_roundCounter_U2 ( .A1 (reset), .A2 (round_Signal[0]), .ZN (controller_roundCounter_N7) ) ;
    INV_X1 controller_roundCounter_U1 ( .A (reset), .ZN (controller_roundCounter_n3) ) ;
    INV_X1 controller_roundCounter_count_reg_0__U1 ( .A (round_Signal[0]), .ZN (controller_roundCounter_n1) ) ;
    INV_X1 controller_roundCounter_count_reg_2__U1 ( .A (round_Signal[2]), .ZN (controller_roundCounter_n6) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U64 ( .a ({new_AGEMA_signal_1458, wk[9]}), .b ({DataIn_s1[9], DataIn_s0[9]}), .c ({new_AGEMA_signal_1790, Midori_add_Result_Start[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U63 ( .a ({new_AGEMA_signal_1461, wk[8]}), .b ({DataIn_s1[8], DataIn_s0[8]}), .c ({new_AGEMA_signal_1792, Midori_add_Result_Start[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U62 ( .a ({new_AGEMA_signal_1464, wk[7]}), .b ({DataIn_s1[7], DataIn_s0[7]}), .c ({new_AGEMA_signal_1794, Midori_add_Result_Start[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U61 ( .a ({new_AGEMA_signal_1467, wk[6]}), .b ({DataIn_s1[6], DataIn_s0[6]}), .c ({new_AGEMA_signal_1796, Midori_add_Result_Start[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U60 ( .a ({new_AGEMA_signal_1470, wk[63]}), .b ({DataIn_s1[63], DataIn_s0[63]}), .c ({new_AGEMA_signal_1798, Midori_add_Result_Start[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U59 ( .a ({new_AGEMA_signal_1473, wk[62]}), .b ({DataIn_s1[62], DataIn_s0[62]}), .c ({new_AGEMA_signal_1800, Midori_add_Result_Start[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U58 ( .a ({new_AGEMA_signal_1476, wk[61]}), .b ({DataIn_s1[61], DataIn_s0[61]}), .c ({new_AGEMA_signal_1802, Midori_add_Result_Start[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U57 ( .a ({new_AGEMA_signal_1479, wk[60]}), .b ({DataIn_s1[60], DataIn_s0[60]}), .c ({new_AGEMA_signal_1804, Midori_add_Result_Start[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U56 ( .a ({new_AGEMA_signal_1482, wk[5]}), .b ({DataIn_s1[5], DataIn_s0[5]}), .c ({new_AGEMA_signal_1806, Midori_add_Result_Start[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U55 ( .a ({new_AGEMA_signal_1485, wk[59]}), .b ({DataIn_s1[59], DataIn_s0[59]}), .c ({new_AGEMA_signal_1808, Midori_add_Result_Start[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U54 ( .a ({new_AGEMA_signal_1488, wk[58]}), .b ({DataIn_s1[58], DataIn_s0[58]}), .c ({new_AGEMA_signal_1810, Midori_add_Result_Start[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U53 ( .a ({new_AGEMA_signal_1491, wk[57]}), .b ({DataIn_s1[57], DataIn_s0[57]}), .c ({new_AGEMA_signal_1812, Midori_add_Result_Start[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U52 ( .a ({new_AGEMA_signal_1494, wk[56]}), .b ({DataIn_s1[56], DataIn_s0[56]}), .c ({new_AGEMA_signal_1814, Midori_add_Result_Start[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U51 ( .a ({new_AGEMA_signal_1497, wk[55]}), .b ({DataIn_s1[55], DataIn_s0[55]}), .c ({new_AGEMA_signal_1816, Midori_add_Result_Start[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U50 ( .a ({new_AGEMA_signal_1500, wk[54]}), .b ({DataIn_s1[54], DataIn_s0[54]}), .c ({new_AGEMA_signal_1818, Midori_add_Result_Start[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U49 ( .a ({new_AGEMA_signal_1503, wk[53]}), .b ({DataIn_s1[53], DataIn_s0[53]}), .c ({new_AGEMA_signal_1820, Midori_add_Result_Start[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U48 ( .a ({new_AGEMA_signal_1506, wk[52]}), .b ({DataIn_s1[52], DataIn_s0[52]}), .c ({new_AGEMA_signal_1822, Midori_add_Result_Start[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U47 ( .a ({new_AGEMA_signal_1509, wk[51]}), .b ({DataIn_s1[51], DataIn_s0[51]}), .c ({new_AGEMA_signal_1824, Midori_add_Result_Start[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U46 ( .a ({new_AGEMA_signal_1512, wk[50]}), .b ({DataIn_s1[50], DataIn_s0[50]}), .c ({new_AGEMA_signal_1826, Midori_add_Result_Start[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U45 ( .a ({new_AGEMA_signal_1515, wk[4]}), .b ({DataIn_s1[4], DataIn_s0[4]}), .c ({new_AGEMA_signal_1828, Midori_add_Result_Start[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U44 ( .a ({new_AGEMA_signal_1518, wk[49]}), .b ({DataIn_s1[49], DataIn_s0[49]}), .c ({new_AGEMA_signal_1830, Midori_add_Result_Start[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U43 ( .a ({new_AGEMA_signal_1521, wk[48]}), .b ({DataIn_s1[48], DataIn_s0[48]}), .c ({new_AGEMA_signal_1832, Midori_add_Result_Start[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U42 ( .a ({new_AGEMA_signal_1524, wk[47]}), .b ({DataIn_s1[47], DataIn_s0[47]}), .c ({new_AGEMA_signal_1834, Midori_add_Result_Start[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U41 ( .a ({new_AGEMA_signal_1527, wk[46]}), .b ({DataIn_s1[46], DataIn_s0[46]}), .c ({new_AGEMA_signal_1836, Midori_add_Result_Start[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U40 ( .a ({new_AGEMA_signal_1530, wk[45]}), .b ({DataIn_s1[45], DataIn_s0[45]}), .c ({new_AGEMA_signal_1838, Midori_add_Result_Start[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U39 ( .a ({new_AGEMA_signal_1533, wk[44]}), .b ({DataIn_s1[44], DataIn_s0[44]}), .c ({new_AGEMA_signal_1840, Midori_add_Result_Start[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U38 ( .a ({new_AGEMA_signal_1536, wk[43]}), .b ({DataIn_s1[43], DataIn_s0[43]}), .c ({new_AGEMA_signal_1842, Midori_add_Result_Start[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U37 ( .a ({new_AGEMA_signal_1539, wk[42]}), .b ({DataIn_s1[42], DataIn_s0[42]}), .c ({new_AGEMA_signal_1844, Midori_add_Result_Start[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U36 ( .a ({new_AGEMA_signal_1542, wk[41]}), .b ({DataIn_s1[41], DataIn_s0[41]}), .c ({new_AGEMA_signal_1846, Midori_add_Result_Start[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U35 ( .a ({new_AGEMA_signal_1545, wk[40]}), .b ({DataIn_s1[40], DataIn_s0[40]}), .c ({new_AGEMA_signal_1848, Midori_add_Result_Start[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U34 ( .a ({new_AGEMA_signal_1548, wk[3]}), .b ({DataIn_s1[3], DataIn_s0[3]}), .c ({new_AGEMA_signal_1850, Midori_add_Result_Start[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U33 ( .a ({new_AGEMA_signal_1551, wk[39]}), .b ({DataIn_s1[39], DataIn_s0[39]}), .c ({new_AGEMA_signal_1852, Midori_add_Result_Start[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U32 ( .a ({new_AGEMA_signal_1554, wk[38]}), .b ({DataIn_s1[38], DataIn_s0[38]}), .c ({new_AGEMA_signal_1854, Midori_add_Result_Start[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U31 ( .a ({new_AGEMA_signal_1557, wk[37]}), .b ({DataIn_s1[37], DataIn_s0[37]}), .c ({new_AGEMA_signal_1856, Midori_add_Result_Start[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U30 ( .a ({new_AGEMA_signal_1560, wk[36]}), .b ({DataIn_s1[36], DataIn_s0[36]}), .c ({new_AGEMA_signal_1858, Midori_add_Result_Start[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U29 ( .a ({new_AGEMA_signal_1563, wk[35]}), .b ({DataIn_s1[35], DataIn_s0[35]}), .c ({new_AGEMA_signal_1860, Midori_add_Result_Start[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U28 ( .a ({new_AGEMA_signal_1566, wk[34]}), .b ({DataIn_s1[34], DataIn_s0[34]}), .c ({new_AGEMA_signal_1862, Midori_add_Result_Start[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U27 ( .a ({new_AGEMA_signal_1569, wk[33]}), .b ({DataIn_s1[33], DataIn_s0[33]}), .c ({new_AGEMA_signal_1864, Midori_add_Result_Start[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U26 ( .a ({new_AGEMA_signal_1572, wk[32]}), .b ({DataIn_s1[32], DataIn_s0[32]}), .c ({new_AGEMA_signal_1866, Midori_add_Result_Start[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U25 ( .a ({new_AGEMA_signal_1575, wk[31]}), .b ({DataIn_s1[31], DataIn_s0[31]}), .c ({new_AGEMA_signal_1868, Midori_add_Result_Start[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U24 ( .a ({new_AGEMA_signal_1578, wk[30]}), .b ({DataIn_s1[30], DataIn_s0[30]}), .c ({new_AGEMA_signal_1870, Midori_add_Result_Start[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U23 ( .a ({new_AGEMA_signal_1581, wk[2]}), .b ({DataIn_s1[2], DataIn_s0[2]}), .c ({new_AGEMA_signal_1872, Midori_add_Result_Start[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U22 ( .a ({new_AGEMA_signal_1584, wk[29]}), .b ({DataIn_s1[29], DataIn_s0[29]}), .c ({new_AGEMA_signal_1874, Midori_add_Result_Start[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U21 ( .a ({new_AGEMA_signal_1587, wk[28]}), .b ({DataIn_s1[28], DataIn_s0[28]}), .c ({new_AGEMA_signal_1876, Midori_add_Result_Start[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U20 ( .a ({new_AGEMA_signal_1590, wk[27]}), .b ({DataIn_s1[27], DataIn_s0[27]}), .c ({new_AGEMA_signal_1878, Midori_add_Result_Start[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U19 ( .a ({new_AGEMA_signal_1593, wk[26]}), .b ({DataIn_s1[26], DataIn_s0[26]}), .c ({new_AGEMA_signal_1880, Midori_add_Result_Start[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U18 ( .a ({new_AGEMA_signal_1596, wk[25]}), .b ({DataIn_s1[25], DataIn_s0[25]}), .c ({new_AGEMA_signal_1882, Midori_add_Result_Start[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U17 ( .a ({new_AGEMA_signal_1599, wk[24]}), .b ({DataIn_s1[24], DataIn_s0[24]}), .c ({new_AGEMA_signal_1884, Midori_add_Result_Start[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U16 ( .a ({new_AGEMA_signal_1602, wk[23]}), .b ({DataIn_s1[23], DataIn_s0[23]}), .c ({new_AGEMA_signal_1886, Midori_add_Result_Start[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U15 ( .a ({new_AGEMA_signal_1605, wk[22]}), .b ({DataIn_s1[22], DataIn_s0[22]}), .c ({new_AGEMA_signal_1888, Midori_add_Result_Start[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U14 ( .a ({new_AGEMA_signal_1608, wk[21]}), .b ({DataIn_s1[21], DataIn_s0[21]}), .c ({new_AGEMA_signal_1890, Midori_add_Result_Start[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U13 ( .a ({new_AGEMA_signal_1611, wk[20]}), .b ({DataIn_s1[20], DataIn_s0[20]}), .c ({new_AGEMA_signal_1892, Midori_add_Result_Start[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U12 ( .a ({new_AGEMA_signal_1614, wk[1]}), .b ({DataIn_s1[1], DataIn_s0[1]}), .c ({new_AGEMA_signal_1894, Midori_add_Result_Start[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U11 ( .a ({new_AGEMA_signal_1617, wk[19]}), .b ({DataIn_s1[19], DataIn_s0[19]}), .c ({new_AGEMA_signal_1896, Midori_add_Result_Start[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U10 ( .a ({new_AGEMA_signal_1620, wk[18]}), .b ({DataIn_s1[18], DataIn_s0[18]}), .c ({new_AGEMA_signal_1898, Midori_add_Result_Start[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U9 ( .a ({new_AGEMA_signal_1623, wk[17]}), .b ({DataIn_s1[17], DataIn_s0[17]}), .c ({new_AGEMA_signal_1900, Midori_add_Result_Start[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U8 ( .a ({new_AGEMA_signal_1626, wk[16]}), .b ({DataIn_s1[16], DataIn_s0[16]}), .c ({new_AGEMA_signal_1902, Midori_add_Result_Start[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U7 ( .a ({new_AGEMA_signal_1629, wk[15]}), .b ({DataIn_s1[15], DataIn_s0[15]}), .c ({new_AGEMA_signal_1904, Midori_add_Result_Start[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U6 ( .a ({new_AGEMA_signal_1632, wk[14]}), .b ({DataIn_s1[14], DataIn_s0[14]}), .c ({new_AGEMA_signal_1906, Midori_add_Result_Start[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U5 ( .a ({new_AGEMA_signal_1635, wk[13]}), .b ({DataIn_s1[13], DataIn_s0[13]}), .c ({new_AGEMA_signal_1908, Midori_add_Result_Start[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U4 ( .a ({new_AGEMA_signal_1638, wk[12]}), .b ({DataIn_s1[12], DataIn_s0[12]}), .c ({new_AGEMA_signal_1910, Midori_add_Result_Start[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U3 ( .a ({new_AGEMA_signal_1641, wk[11]}), .b ({DataIn_s1[11], DataIn_s0[11]}), .c ({new_AGEMA_signal_1912, Midori_add_Result_Start[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U2 ( .a ({new_AGEMA_signal_1644, wk[10]}), .b ({DataIn_s1[10], DataIn_s0[10]}), .c ({new_AGEMA_signal_1914, Midori_add_Result_Start[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U1 ( .a ({new_AGEMA_signal_1647, wk[0]}), .b ({DataIn_s1[0], DataIn_s0[0]}), .c ({new_AGEMA_signal_1916, Midori_add_Result_Start[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U78 ( .a ({new_AGEMA_signal_1653, Midori_rounds_SelectedKey_8_}), .b ({1'b0, Midori_rounds_round_Constant[2]}), .c ({new_AGEMA_signal_2441, Midori_rounds_n16}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U71 ( .a ({new_AGEMA_signal_2060, Midori_rounds_SelectedKey_60_}), .b ({1'b0, Midori_rounds_round_Constant[15]}), .c ({new_AGEMA_signal_2496, Midori_rounds_n15}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U65 ( .a ({new_AGEMA_signal_2056, Midori_rounds_SelectedKey_56_}), .b ({1'b0, Midori_rounds_round_Constant[14]}), .c ({new_AGEMA_signal_2497, Midori_rounds_n14}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U60 ( .a ({new_AGEMA_signal_2052, Midori_rounds_SelectedKey_52_}), .b ({1'b0, Midori_rounds_round_Constant[13]}), .c ({new_AGEMA_signal_2498, Midori_rounds_n13}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U56 ( .a ({new_AGEMA_signal_1652, Midori_rounds_SelectedKey_4_}), .b ({1'b0, Midori_rounds_round_Constant[1]}), .c ({new_AGEMA_signal_2499, Midori_rounds_n12}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U53 ( .a ({new_AGEMA_signal_2048, Midori_rounds_SelectedKey_48_}), .b ({1'b0, Midori_rounds_round_Constant[12]}), .c ({new_AGEMA_signal_2618, Midori_rounds_n11}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U48 ( .a ({new_AGEMA_signal_2044, Midori_rounds_SelectedKey_44_}), .b ({1'b0, Midori_rounds_round_Constant[11]}), .c ({new_AGEMA_signal_2460, Midori_rounds_n10}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U43 ( .a ({new_AGEMA_signal_2040, Midori_rounds_SelectedKey_40_}), .b ({1'b0, Midori_rounds_round_Constant[10]}), .c ({new_AGEMA_signal_2500, Midori_rounds_n9}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U37 ( .a ({new_AGEMA_signal_2036, Midori_rounds_SelectedKey_36_}), .b ({1'b0, Midori_rounds_round_Constant[9]}), .c ({new_AGEMA_signal_2468, Midori_rounds_n8}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U32 ( .a ({new_AGEMA_signal_2032, Midori_rounds_SelectedKey_32_}), .b ({1'b0, Midori_rounds_round_Constant[8]}), .c ({new_AGEMA_signal_2501, Midori_rounds_n7}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U26 ( .a ({new_AGEMA_signal_2028, Midori_rounds_SelectedKey_28_}), .b ({1'b0, Midori_rounds_round_Constant[7]}), .c ({new_AGEMA_signal_2564, Midori_rounds_n6}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U21 ( .a ({new_AGEMA_signal_2025, Midori_rounds_SelectedKey_24_}), .b ({1'b0, Midori_rounds_round_Constant[6]}), .c ({new_AGEMA_signal_2502, Midori_rounds_n5}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U16 ( .a ({new_AGEMA_signal_2021, Midori_rounds_SelectedKey_20_}), .b ({1'b0, Midori_rounds_round_Constant[5]}), .c ({new_AGEMA_signal_2482, Midori_rounds_n4}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U10 ( .a ({new_AGEMA_signal_2017, Midori_rounds_SelectedKey_16_}), .b ({1'b0, Midori_rounds_round_Constant[4]}), .c ({new_AGEMA_signal_2503, Midori_rounds_n3}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U5 ( .a ({new_AGEMA_signal_2016, Midori_rounds_SelectedKey_12_}), .b ({1'b0, Midori_rounds_round_Constant[3]}), .c ({new_AGEMA_signal_2504, Midori_rounds_n2}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U1 ( .a ({new_AGEMA_signal_1648, Midori_rounds_SelectedKey_0_}), .b ({1'b0, Midori_rounds_round_Constant[0]}), .c ({new_AGEMA_signal_2505, Midori_rounds_n1}) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U106 ( .A1 (Midori_rounds_constant_MUX_n217), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_round_Constant[9]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U105 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n214), .ZN (Midori_rounds_constant_MUX_n217) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U104 ( .A1 (Midori_rounds_constant_MUX_n213), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n214) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U103 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_round_Constant[8]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U102 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n208), .ZN (Midori_rounds_round_Constant[7]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U101 ( .A1 (Midori_rounds_round_Constant[11]), .A2 (Midori_rounds_constant_MUX_n207), .ZN (Midori_rounds_constant_MUX_n208) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U100 ( .A1 (Midori_rounds_constant_MUX_n206), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n207) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U99 ( .A1 (Midori_rounds_constant_MUX_n204), .A2 (Midori_rounds_constant_MUX_n203), .ZN (Midori_rounds_constant_MUX_n206) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U98 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n201), .ZN (Midori_rounds_round_Constant[6]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U97 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n199), .ZN (Midori_rounds_constant_MUX_n201) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U96 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n197), .ZN (Midori_rounds_round_Constant[5]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U95 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n196), .ZN (Midori_rounds_constant_MUX_n197) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U94 ( .A1 (Midori_rounds_constant_MUX_n195), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n196) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U93 ( .A1 (Midori_rounds_constant_MUX_n194), .A2 (Midori_rounds_constant_MUX_n195), .ZN (Midori_rounds_round_Constant[4]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U92 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n195) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U91 ( .A1 (Midori_rounds_constant_MUX_n191), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[3]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U90 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n189), .ZN (Midori_rounds_constant_MUX_n191) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U89 ( .A1 (Midori_rounds_constant_MUX_n188), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n189) ) ;
    INV_X1 Midori_rounds_constant_MUX_U88 ( .A (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n188) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U87 ( .A1 (Midori_rounds_constant_MUX_n215), .A2 (Midori_rounds_constant_MUX_n186), .ZN (Midori_rounds_round_Constant[2]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U86 ( .A1 (Midori_rounds_constant_MUX_n202), .A2 (Midori_rounds_constant_MUX_n185), .ZN (Midori_rounds_constant_MUX_n186) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U85 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n212), .ZN (Midori_rounds_constant_MUX_n202) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U84 ( .A1 (Midori_rounds_constant_MUX_n183), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n215) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U83 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n181), .ZN (Midori_rounds_round_Constant[1]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U82 ( .A1 (Midori_rounds_constant_MUX_n187), .A2 (Midori_rounds_constant_MUX_n180), .ZN (Midori_rounds_constant_MUX_n181) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U81 ( .A1 (Midori_rounds_constant_MUX_n212), .A2 (Midori_rounds_constant_MUX_n204), .ZN (Midori_rounds_constant_MUX_n180) ) ;
    INV_X1 Midori_rounds_constant_MUX_U80 ( .A (Midori_rounds_constant_MUX_n183), .ZN (Midori_rounds_constant_MUX_n204) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U79 ( .A1 (Midori_rounds_constant_MUX_n179), .A2 (Midori_rounds_constant_MUX_n178), .ZN (Midori_rounds_constant_MUX_n183) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U78 ( .A1 (Midori_rounds_constant_MUX_n177), .A2 (Midori_rounds_constant_MUX_n176), .ZN (Midori_rounds_constant_MUX_n178) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U77 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n175), .ZN (Midori_rounds_constant_MUX_n212) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U76 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n173), .Z (Midori_rounds_constant_MUX_n175) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U75 ( .A1 (Midori_rounds_constant_MUX_n172), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[15]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U74 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n172) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U73 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n194), .ZN (Midori_rounds_round_Constant[14]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U72 ( .A1 (Midori_rounds_constant_MUX_n169), .A2 (Midori_rounds_constant_MUX_n168), .ZN (Midori_rounds_constant_MUX_n194) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U71 ( .A1 (Midori_rounds_constant_MUX_n216), .A2 (Midori_rounds_constant_MUX_n205), .ZN (Midori_rounds_constant_MUX_n168) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U70 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n167), .ZN (Midori_rounds_constant_MUX_n205) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U69 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n167) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U68 ( .A1 (Midori_rounds_constant_MUX_n185), .A2 (Midori_rounds_constant_MUX_n164), .ZN (Midori_rounds_round_Constant[13]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U67 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n162), .ZN (Midori_rounds_constant_MUX_n164) ) ;
    INV_X1 Midori_rounds_constant_MUX_U66 ( .A (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n162) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U65 ( .A1 (Midori_rounds_constant_MUX_n161), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n185) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U64 ( .A1 (Midori_rounds_constant_MUX_n160), .A2 (Midori_rounds_constant_MUX_n190), .ZN (Midori_rounds_round_Constant[12]) ) ;
    INV_X1 Midori_rounds_constant_MUX_U63 ( .A (Midori_rounds_constant_MUX_n184), .ZN (Midori_rounds_constant_MUX_n190) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U62 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n159), .ZN (Midori_rounds_constant_MUX_n160) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U61 ( .A1 (Midori_rounds_constant_MUX_n211), .A2 (Midori_rounds_constant_MUX_n170), .ZN (Midori_rounds_constant_MUX_n159) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U60 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n169), .ZN (Midori_rounds_constant_MUX_n211) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U59 ( .A1 (Midori_rounds_constant_MUX_n198), .A2 (Midori_rounds_constant_MUX_n158), .ZN (Midori_rounds_constant_MUX_n169) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U58 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n157), .ZN (Midori_rounds_constant_MUX_n158) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U57 ( .A1 (Midori_rounds_constant_MUX_n165), .A2 (Midori_rounds_constant_MUX_n177), .ZN (Midori_rounds_constant_MUX_n157) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U56 ( .A1 (Midori_rounds_constant_MUX_n200), .A2 (Midori_rounds_constant_MUX_n156), .ZN (Midori_rounds_constant_MUX_n198) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U55 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n155), .ZN (Midori_rounds_constant_MUX_n156) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U54 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n176), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n155) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U53 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n154), .ZN (Midori_rounds_constant_MUX_n200) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U52 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n174), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n154) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U51 ( .A1 (Midori_rounds_constant_MUX_n199), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_round_Constant[11]) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U50 ( .A1 (Midori_rounds_constant_MUX_n170), .A2 (Midori_rounds_constant_MUX_n210), .ZN (Midori_rounds_constant_MUX_n199) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U49 ( .A1 (Midori_rounds_constant_MUX_n152), .A2 (Midori_rounds_constant_MUX_n151), .ZN (Midori_rounds_constant_MUX_n210) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U48 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n151) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U47 ( .A1 (Midori_rounds_constant_MUX_n150), .A2 (Midori_rounds_constant_MUX_n187), .ZN (Midori_rounds_constant_MUX_n170) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U46 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n149), .ZN (Midori_rounds_constant_MUX_n187) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U45 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n166), .Z (Midori_rounds_constant_MUX_n149) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U44 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (Midori_rounds_constant_MUX_n148), .ZN (Midori_rounds_constant_MUX_n150) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U43 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n148) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U42 ( .A1 (Midori_rounds_constant_MUX_n147), .A2 (Midori_rounds_constant_MUX_n171), .ZN (Midori_rounds_round_Constant[10]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U41 ( .A1 (Midori_rounds_constant_MUX_n146), .A2 (Midori_rounds_constant_MUX_n213), .ZN (Midori_rounds_constant_MUX_n171) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U40 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n145), .ZN (Midori_rounds_constant_MUX_n213) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U39 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n165), .B (Midori_rounds_constant_MUX_n177), .Z (Midori_rounds_constant_MUX_n145) ) ;
    INV_X1 Midori_rounds_constant_MUX_U38 ( .A (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_constant_MUX_n146) ) ;
    INV_X1 Midori_rounds_constant_MUX_U37 ( .A (Midori_rounds_constant_MUX_n193), .ZN (Midori_rounds_constant_MUX_n147) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U36 ( .A1 (Midori_rounds_constant_MUX_n182), .A2 (Midori_rounds_constant_MUX_n144), .ZN (Midori_rounds_round_Constant[0]) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U35 ( .A1 (Midori_rounds_constant_MUX_n203), .A2 (Midori_rounds_constant_MUX_n192), .ZN (Midori_rounds_constant_MUX_n144) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U34 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n143), .ZN (Midori_rounds_constant_MUX_n192) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U33 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n173), .B (Midori_rounds_constant_MUX_n174), .Z (Midori_rounds_constant_MUX_n143) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U32 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n174) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U31 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n173) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U30 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n139), .ZN (Midori_rounds_constant_MUX_n203) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U29 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n166), .B (Midori_rounds_constant_MUX_n176), .Z (Midori_rounds_constant_MUX_n139) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U28 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n152), .ZN (Midori_rounds_constant_MUX_n176) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U27 ( .A1 (round_Signal[3]), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n152) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U26 ( .A1 (Midori_rounds_constant_MUX_n138), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n166) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U25 ( .A1 (Midori_rounds_constant_MUX_n184), .A2 (Midori_rounds_constant_MUX_n137), .ZN (Midori_rounds_constant_MUX_n182) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U24 ( .A1 (Midori_rounds_constant_MUX_n209), .A2 (Midori_rounds_constant_MUX_n216), .ZN (Midori_rounds_constant_MUX_n137) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U23 ( .A1 (Midori_rounds_constant_MUX_n163), .A2 (Midori_rounds_constant_MUX_n136), .ZN (Midori_rounds_constant_MUX_n216) ) ;
    OR2_X1 Midori_rounds_constant_MUX_U22 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n142), .ZN (Midori_rounds_constant_MUX_n136) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U21 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n179), .ZN (Midori_rounds_constant_MUX_n163) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U20 ( .A1 (Midori_rounds_constant_MUX_n129), .A2 (round_Signal[2]), .ZN (Midori_rounds_constant_MUX_n179) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U19 ( .A1 (Midori_rounds_constant_MUX_n193), .A2 (Midori_rounds_constant_MUX_n161), .ZN (Midori_rounds_constant_MUX_n209) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U18 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n135), .ZN (Midori_rounds_constant_MUX_n161) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U17 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n177), .B (Midori_rounds_constant_MUX_n165), .Z (Midori_rounds_constant_MUX_n135) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U16 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n134), .ZN (Midori_rounds_constant_MUX_n165) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U15 ( .A1 (round_Signal[3]), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n134) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U14 ( .A1 (round_Signal[1]), .A2 (Midori_rounds_constant_MUX_n138), .ZN (Midori_rounds_constant_MUX_n177) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U13 ( .A1 (enc_dec), .A2 (Midori_rounds_constant_MUX_n133), .ZN (Midori_rounds_constant_MUX_n138) ) ;
    INV_X1 Midori_rounds_constant_MUX_U12 ( .A (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n133) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U11 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n132), .ZN (Midori_rounds_constant_MUX_n193) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U10 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n153), .B (Midori_rounds_constant_MUX_n131), .Z (Midori_rounds_constant_MUX_n132) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U9 ( .A1 (Midori_rounds_constant_MUX_n128), .A2 (Midori_rounds_constant_MUX_n130), .ZN (Midori_rounds_constant_MUX_n184) ) ;
    MUX2_X1 Midori_rounds_constant_MUX_U8 ( .S (round_Signal[2]), .A (Midori_rounds_constant_MUX_n131), .B (Midori_rounds_constant_MUX_n153), .Z (Midori_rounds_constant_MUX_n130) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U7 ( .A1 (Midori_rounds_constant_MUX_n140), .A2 (Midori_rounds_constant_MUX_n141), .ZN (Midori_rounds_constant_MUX_n153) ) ;
    INV_X1 Midori_rounds_constant_MUX_U6 ( .A (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n141) ) ;
    NOR2_X1 Midori_rounds_constant_MUX_U5 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n140) ) ;
    NAND2_X1 Midori_rounds_constant_MUX_U4 ( .A1 (Midori_rounds_constant_MUX_n142), .A2 (round_Signal[1]), .ZN (Midori_rounds_constant_MUX_n131) ) ;
    AND2_X1 Midori_rounds_constant_MUX_U3 ( .A1 (enc_dec), .A2 (round_Signal[3]), .ZN (Midori_rounds_constant_MUX_n142) ) ;
    INV_X1 Midori_rounds_constant_MUX_U2 ( .A (Midori_rounds_constant_MUX_n129), .ZN (Midori_rounds_constant_MUX_n128) ) ;
    INV_X1 Midori_rounds_constant_MUX_U1 ( .A (round_Signal[0]), .ZN (Midori_rounds_constant_MUX_n129) ) ;
    INV_X1 Midori_rounds_MUXInst_U4 ( .A (round_Signal[0]), .ZN (Midori_rounds_MUXInst_n11) ) ;
    INV_X1 Midori_rounds_MUXInst_U3 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n8) ) ;
    INV_X1 Midori_rounds_MUXInst_U2 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n9) ) ;
    INV_X1 Midori_rounds_MUXInst_U1 ( .A (Midori_rounds_MUXInst_n11), .ZN (Midori_rounds_MUXInst_n10) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_0_U1 ( .s (round_Signal[0]), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1648, Midori_rounds_SelectedKey_0_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_1_U1 ( .s (round_Signal[0]), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1649, Midori_rounds_SelectedKey_1_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_2_U1 ( .s (round_Signal[0]), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1650, Midori_rounds_SelectedKey_2_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_3_U1 ( .s (round_Signal[0]), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1651, Midori_rounds_SelectedKey_3_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_4_U1 ( .s (round_Signal[0]), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1652, Midori_rounds_SelectedKey_4_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_5_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_2013, Midori_rounds_SelectedKey_5_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_6_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_2014, Midori_rounds_SelectedKey_6_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_7_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_2015, Midori_rounds_SelectedKey_7_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_8_U1 ( .s (round_Signal[0]), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1653, Midori_rounds_SelectedKey_8_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_9_U1 ( .s (round_Signal[0]), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1654, Midori_rounds_SelectedKey_9_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_10_U1 ( .s (round_Signal[0]), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1655, Midori_rounds_SelectedKey_10_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_11_U1 ( .s (round_Signal[0]), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1656, Midori_rounds_SelectedKey_11_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_12_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_2016, Midori_rounds_SelectedKey_12_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_13_U1 ( .s (round_Signal[0]), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1657, Midori_rounds_SelectedKey_13_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_14_U1 ( .s (round_Signal[0]), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1658, Midori_rounds_SelectedKey_14_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_15_U1 ( .s (round_Signal[0]), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1659, Midori_rounds_SelectedKey_15_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_16_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_2017, Midori_rounds_SelectedKey_16_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_17_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_2018, Midori_rounds_SelectedKey_17_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_18_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_2019, Midori_rounds_SelectedKey_18_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_19_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_2020, Midori_rounds_SelectedKey_19_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_20_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_2021, Midori_rounds_SelectedKey_20_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_21_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_2022, Midori_rounds_SelectedKey_21_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_22_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_2023, Midori_rounds_SelectedKey_22_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_23_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_2024, Midori_rounds_SelectedKey_23_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_24_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_2025, Midori_rounds_SelectedKey_24_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_25_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_2026, Midori_rounds_SelectedKey_25_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_26_U1 ( .s (round_Signal[0]), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1660, Midori_rounds_SelectedKey_26_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_27_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_2027, Midori_rounds_SelectedKey_27_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_28_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_2028, Midori_rounds_SelectedKey_28_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_29_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_2029, Midori_rounds_SelectedKey_29_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_30_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_2030, Midori_rounds_SelectedKey_30_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_31_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_2031, Midori_rounds_SelectedKey_31_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_32_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2032, Midori_rounds_SelectedKey_32_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_33_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_2033, Midori_rounds_SelectedKey_33_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_34_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2034, Midori_rounds_SelectedKey_34_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_35_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2035, Midori_rounds_SelectedKey_35_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_36_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_2036, Midori_rounds_SelectedKey_36_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_37_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2037, Midori_rounds_SelectedKey_37_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_38_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2038, Midori_rounds_SelectedKey_38_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_39_U1 ( .s (Midori_rounds_MUXInst_n10), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_2039, Midori_rounds_SelectedKey_39_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_40_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2040, Midori_rounds_SelectedKey_40_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_41_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2041, Midori_rounds_SelectedKey_41_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_42_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2042, Midori_rounds_SelectedKey_42_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_43_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2043, Midori_rounds_SelectedKey_43_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_44_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2044, Midori_rounds_SelectedKey_44_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_45_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2045, Midori_rounds_SelectedKey_45_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_46_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2046, Midori_rounds_SelectedKey_46_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_47_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2047, Midori_rounds_SelectedKey_47_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_48_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2048, Midori_rounds_SelectedKey_48_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_49_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2049, Midori_rounds_SelectedKey_49_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_50_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2050, Midori_rounds_SelectedKey_50_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_51_U1 ( .s (Midori_rounds_MUXInst_n9), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2051, Midori_rounds_SelectedKey_51_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_52_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2052, Midori_rounds_SelectedKey_52_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_53_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_2053, Midori_rounds_SelectedKey_53_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_54_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_2054, Midori_rounds_SelectedKey_54_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_55_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2055, Midori_rounds_SelectedKey_55_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_56_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_2056, Midori_rounds_SelectedKey_56_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_57_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2057, Midori_rounds_SelectedKey_57_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_58_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2058, Midori_rounds_SelectedKey_58_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_59_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_2059, Midori_rounds_SelectedKey_59_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_60_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2060, Midori_rounds_SelectedKey_60_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_61_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2061, Midori_rounds_SelectedKey_61_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_62_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_2062, Midori_rounds_SelectedKey_62_}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_MUXInst_mux_inst_63_U1 ( .s (Midori_rounds_MUXInst_n8), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2063, Midori_rounds_SelectedKey_63_}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U4 ( .a ({new_AGEMA_signal_1661, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1666, Midori_rounds_sub_sBox_PRINCE_0_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U2 ( .a ({new_AGEMA_signal_1662, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1667, Midori_rounds_sub_sBox_PRINCE_0_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U1 ( .a ({new_AGEMA_signal_1664, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1668, Midori_rounds_sub_sBox_PRINCE_0_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .a ({new_AGEMA_signal_1669, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1674, Midori_rounds_sub_sBox_PRINCE_1_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U2 ( .a ({new_AGEMA_signal_1670, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1675, Midori_rounds_sub_sBox_PRINCE_1_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .a ({new_AGEMA_signal_1672, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1676, Midori_rounds_sub_sBox_PRINCE_1_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .a ({new_AGEMA_signal_1677, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1682, Midori_rounds_sub_sBox_PRINCE_2_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U2 ( .a ({new_AGEMA_signal_1678, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1683, Midori_rounds_sub_sBox_PRINCE_2_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .a ({new_AGEMA_signal_1680, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1684, Midori_rounds_sub_sBox_PRINCE_2_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .a ({new_AGEMA_signal_1685, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1690, Midori_rounds_sub_sBox_PRINCE_3_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U2 ( .a ({new_AGEMA_signal_1686, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1691, Midori_rounds_sub_sBox_PRINCE_3_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .a ({new_AGEMA_signal_1688, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1692, Midori_rounds_sub_sBox_PRINCE_3_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .a ({new_AGEMA_signal_1693, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1698, Midori_rounds_sub_sBox_PRINCE_4_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U2 ( .a ({new_AGEMA_signal_1694, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1699, Midori_rounds_sub_sBox_PRINCE_4_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .a ({new_AGEMA_signal_1696, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1700, Midori_rounds_sub_sBox_PRINCE_4_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .a ({new_AGEMA_signal_1701, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1706, Midori_rounds_sub_sBox_PRINCE_5_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U2 ( .a ({new_AGEMA_signal_1702, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1707, Midori_rounds_sub_sBox_PRINCE_5_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .a ({new_AGEMA_signal_1704, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1708, Midori_rounds_sub_sBox_PRINCE_5_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .a ({new_AGEMA_signal_1709, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1714, Midori_rounds_sub_sBox_PRINCE_6_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U2 ( .a ({new_AGEMA_signal_1710, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1715, Midori_rounds_sub_sBox_PRINCE_6_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .a ({new_AGEMA_signal_1712, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1716, Midori_rounds_sub_sBox_PRINCE_6_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U4 ( .a ({new_AGEMA_signal_1717, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1722, Midori_rounds_sub_sBox_PRINCE_7_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U2 ( .a ({new_AGEMA_signal_1718, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1723, Midori_rounds_sub_sBox_PRINCE_7_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U1 ( .a ({new_AGEMA_signal_1720, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1724, Midori_rounds_sub_sBox_PRINCE_7_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U4 ( .a ({new_AGEMA_signal_1725, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_1730, Midori_rounds_sub_sBox_PRINCE_8_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U2 ( .a ({new_AGEMA_signal_1726, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_1731, Midori_rounds_sub_sBox_PRINCE_8_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U1 ( .a ({new_AGEMA_signal_1728, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_1732, Midori_rounds_sub_sBox_PRINCE_8_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U4 ( .a ({new_AGEMA_signal_1733, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_1738, Midori_rounds_sub_sBox_PRINCE_9_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U2 ( .a ({new_AGEMA_signal_1734, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_1739, Midori_rounds_sub_sBox_PRINCE_9_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U1 ( .a ({new_AGEMA_signal_1736, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_1740, Midori_rounds_sub_sBox_PRINCE_9_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .a ({new_AGEMA_signal_1741, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_1746, Midori_rounds_sub_sBox_PRINCE_10_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U2 ( .a ({new_AGEMA_signal_1742, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_1747, Midori_rounds_sub_sBox_PRINCE_10_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .a ({new_AGEMA_signal_1744, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_1748, Midori_rounds_sub_sBox_PRINCE_10_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .a ({new_AGEMA_signal_1749, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_1754, Midori_rounds_sub_sBox_PRINCE_11_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U2 ( .a ({new_AGEMA_signal_1750, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_1755, Midori_rounds_sub_sBox_PRINCE_11_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .a ({new_AGEMA_signal_1752, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_1756, Midori_rounds_sub_sBox_PRINCE_11_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .a ({new_AGEMA_signal_1757, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_1762, Midori_rounds_sub_sBox_PRINCE_12_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U2 ( .a ({new_AGEMA_signal_1758, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_1763, Midori_rounds_sub_sBox_PRINCE_12_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .a ({new_AGEMA_signal_1760, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_1764, Midori_rounds_sub_sBox_PRINCE_12_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U4 ( .a ({new_AGEMA_signal_1765, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_1770, Midori_rounds_sub_sBox_PRINCE_13_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U2 ( .a ({new_AGEMA_signal_1766, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_1771, Midori_rounds_sub_sBox_PRINCE_13_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U1 ( .a ({new_AGEMA_signal_1768, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_1772, Midori_rounds_sub_sBox_PRINCE_13_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U4 ( .a ({new_AGEMA_signal_1773, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_1778, Midori_rounds_sub_sBox_PRINCE_14_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U2 ( .a ({new_AGEMA_signal_1774, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_1779, Midori_rounds_sub_sBox_PRINCE_14_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U1 ( .a ({new_AGEMA_signal_1776, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_1780, Midori_rounds_sub_sBox_PRINCE_14_n9}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .a ({new_AGEMA_signal_1781, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_1786, Midori_rounds_sub_sBox_PRINCE_15_n7}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U2 ( .a ({new_AGEMA_signal_1782, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_1787, Midori_rounds_sub_sBox_PRINCE_15_n8}) ) ;
    not_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .a ({new_AGEMA_signal_1784, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_1788, Midori_rounds_sub_sBox_PRINCE_15_n9}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_3024), .Q (new_AGEMA_signal_3025) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (clk), .D (Midori_rounds_roundReg_out[1]), .Q (new_AGEMA_signal_3096) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (clk), .D (new_AGEMA_signal_2064), .Q (new_AGEMA_signal_3098) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n9), .Q (new_AGEMA_signal_3100) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (clk), .D (new_AGEMA_signal_1668), .Q (new_AGEMA_signal_3102) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (clk), .D (Midori_rounds_roundReg_out[0]), .Q (new_AGEMA_signal_3104) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (clk), .D (new_AGEMA_signal_1661), .Q (new_AGEMA_signal_3106) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n7), .Q (new_AGEMA_signal_3108) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (clk), .D (new_AGEMA_signal_1666), .Q (new_AGEMA_signal_3110) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (clk), .D (Midori_rounds_roundReg_out[5]), .Q (new_AGEMA_signal_3112) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (clk), .D (new_AGEMA_signal_2069), .Q (new_AGEMA_signal_3114) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n9), .Q (new_AGEMA_signal_3116) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (clk), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_3118) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (clk), .D (Midori_rounds_roundReg_out[4]), .Q (new_AGEMA_signal_3120) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (clk), .D (new_AGEMA_signal_1669), .Q (new_AGEMA_signal_3122) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n7), .Q (new_AGEMA_signal_3124) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (clk), .D (new_AGEMA_signal_1674), .Q (new_AGEMA_signal_3126) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (clk), .D (Midori_rounds_roundReg_out[9]), .Q (new_AGEMA_signal_3128) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (clk), .D (new_AGEMA_signal_2074), .Q (new_AGEMA_signal_3130) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n9), .Q (new_AGEMA_signal_3132) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (clk), .D (new_AGEMA_signal_1684), .Q (new_AGEMA_signal_3134) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (clk), .D (Midori_rounds_roundReg_out[8]), .Q (new_AGEMA_signal_3136) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (clk), .D (new_AGEMA_signal_1677), .Q (new_AGEMA_signal_3138) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n7), .Q (new_AGEMA_signal_3140) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (clk), .D (new_AGEMA_signal_1682), .Q (new_AGEMA_signal_3142) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (clk), .D (Midori_rounds_roundReg_out[13]), .Q (new_AGEMA_signal_3144) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (clk), .D (new_AGEMA_signal_2079), .Q (new_AGEMA_signal_3146) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n9), .Q (new_AGEMA_signal_3148) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (clk), .D (new_AGEMA_signal_1692), .Q (new_AGEMA_signal_3150) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (clk), .D (Midori_rounds_roundReg_out[12]), .Q (new_AGEMA_signal_3152) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (clk), .D (new_AGEMA_signal_1685), .Q (new_AGEMA_signal_3154) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n7), .Q (new_AGEMA_signal_3156) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (clk), .D (new_AGEMA_signal_1690), .Q (new_AGEMA_signal_3158) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (clk), .D (Midori_rounds_roundReg_out[17]), .Q (new_AGEMA_signal_3160) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (clk), .D (new_AGEMA_signal_2084), .Q (new_AGEMA_signal_3162) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n9), .Q (new_AGEMA_signal_3164) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (clk), .D (new_AGEMA_signal_1700), .Q (new_AGEMA_signal_3166) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (clk), .D (Midori_rounds_roundReg_out[16]), .Q (new_AGEMA_signal_3168) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (clk), .D (new_AGEMA_signal_1693), .Q (new_AGEMA_signal_3170) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n7), .Q (new_AGEMA_signal_3172) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (clk), .D (new_AGEMA_signal_1698), .Q (new_AGEMA_signal_3174) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (clk), .D (Midori_rounds_roundReg_out[21]), .Q (new_AGEMA_signal_3176) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (clk), .D (new_AGEMA_signal_2089), .Q (new_AGEMA_signal_3178) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n9), .Q (new_AGEMA_signal_3180) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (clk), .D (new_AGEMA_signal_1708), .Q (new_AGEMA_signal_3182) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (clk), .D (Midori_rounds_roundReg_out[20]), .Q (new_AGEMA_signal_3184) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (clk), .D (new_AGEMA_signal_1701), .Q (new_AGEMA_signal_3186) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n7), .Q (new_AGEMA_signal_3188) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (clk), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_3190) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (clk), .D (Midori_rounds_roundReg_out[25]), .Q (new_AGEMA_signal_3192) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (clk), .D (new_AGEMA_signal_2094), .Q (new_AGEMA_signal_3194) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n9), .Q (new_AGEMA_signal_3196) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (clk), .D (new_AGEMA_signal_1716), .Q (new_AGEMA_signal_3198) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (clk), .D (Midori_rounds_roundReg_out[24]), .Q (new_AGEMA_signal_3200) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (clk), .D (new_AGEMA_signal_1709), .Q (new_AGEMA_signal_3202) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n7), .Q (new_AGEMA_signal_3204) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (clk), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_3206) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (clk), .D (Midori_rounds_roundReg_out[29]), .Q (new_AGEMA_signal_3208) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (clk), .D (new_AGEMA_signal_2099), .Q (new_AGEMA_signal_3210) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n9), .Q (new_AGEMA_signal_3212) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (clk), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_3214) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (clk), .D (Midori_rounds_roundReg_out[28]), .Q (new_AGEMA_signal_3216) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (clk), .D (new_AGEMA_signal_1717), .Q (new_AGEMA_signal_3218) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n7), .Q (new_AGEMA_signal_3220) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (clk), .D (new_AGEMA_signal_1722), .Q (new_AGEMA_signal_3222) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (clk), .D (Midori_rounds_roundReg_out[33]), .Q (new_AGEMA_signal_3224) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (clk), .D (new_AGEMA_signal_2104), .Q (new_AGEMA_signal_3226) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n9), .Q (new_AGEMA_signal_3228) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (clk), .D (new_AGEMA_signal_1732), .Q (new_AGEMA_signal_3230) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (clk), .D (Midori_rounds_roundReg_out[32]), .Q (new_AGEMA_signal_3232) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (clk), .D (new_AGEMA_signal_1725), .Q (new_AGEMA_signal_3234) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n7), .Q (new_AGEMA_signal_3236) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (clk), .D (new_AGEMA_signal_1730), .Q (new_AGEMA_signal_3238) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (clk), .D (Midori_rounds_roundReg_out[37]), .Q (new_AGEMA_signal_3240) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (clk), .D (new_AGEMA_signal_2109), .Q (new_AGEMA_signal_3242) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n9), .Q (new_AGEMA_signal_3244) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (clk), .D (new_AGEMA_signal_1740), .Q (new_AGEMA_signal_3246) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (clk), .D (Midori_rounds_roundReg_out[36]), .Q (new_AGEMA_signal_3248) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (clk), .D (new_AGEMA_signal_1733), .Q (new_AGEMA_signal_3250) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n7), .Q (new_AGEMA_signal_3252) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (clk), .D (new_AGEMA_signal_1738), .Q (new_AGEMA_signal_3254) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (clk), .D (Midori_rounds_roundReg_out[41]), .Q (new_AGEMA_signal_3256) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (clk), .D (new_AGEMA_signal_2114), .Q (new_AGEMA_signal_3258) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n9), .Q (new_AGEMA_signal_3260) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (clk), .D (new_AGEMA_signal_1748), .Q (new_AGEMA_signal_3262) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (clk), .D (Midori_rounds_roundReg_out[40]), .Q (new_AGEMA_signal_3264) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (clk), .D (new_AGEMA_signal_1741), .Q (new_AGEMA_signal_3266) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n7), .Q (new_AGEMA_signal_3268) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (clk), .D (new_AGEMA_signal_1746), .Q (new_AGEMA_signal_3270) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (clk), .D (Midori_rounds_roundReg_out[45]), .Q (new_AGEMA_signal_3272) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (clk), .D (new_AGEMA_signal_2119), .Q (new_AGEMA_signal_3274) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n9), .Q (new_AGEMA_signal_3276) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (clk), .D (new_AGEMA_signal_1756), .Q (new_AGEMA_signal_3278) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (clk), .D (Midori_rounds_roundReg_out[44]), .Q (new_AGEMA_signal_3280) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (clk), .D (new_AGEMA_signal_1749), .Q (new_AGEMA_signal_3282) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n7), .Q (new_AGEMA_signal_3284) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (clk), .D (new_AGEMA_signal_1754), .Q (new_AGEMA_signal_3286) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (clk), .D (Midori_rounds_roundReg_out[49]), .Q (new_AGEMA_signal_3288) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (clk), .D (new_AGEMA_signal_2124), .Q (new_AGEMA_signal_3290) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n9), .Q (new_AGEMA_signal_3292) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (clk), .D (new_AGEMA_signal_1764), .Q (new_AGEMA_signal_3294) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (clk), .D (Midori_rounds_roundReg_out[48]), .Q (new_AGEMA_signal_3296) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (clk), .D (new_AGEMA_signal_1757), .Q (new_AGEMA_signal_3298) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n7), .Q (new_AGEMA_signal_3300) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (clk), .D (new_AGEMA_signal_1762), .Q (new_AGEMA_signal_3302) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (clk), .D (Midori_rounds_roundReg_out[53]), .Q (new_AGEMA_signal_3304) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (clk), .D (new_AGEMA_signal_2129), .Q (new_AGEMA_signal_3306) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n9), .Q (new_AGEMA_signal_3308) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (clk), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_3310) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (clk), .D (Midori_rounds_roundReg_out[52]), .Q (new_AGEMA_signal_3312) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (clk), .D (new_AGEMA_signal_1765), .Q (new_AGEMA_signal_3314) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n7), .Q (new_AGEMA_signal_3316) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (clk), .D (new_AGEMA_signal_1770), .Q (new_AGEMA_signal_3318) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (clk), .D (Midori_rounds_roundReg_out[57]), .Q (new_AGEMA_signal_3320) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (clk), .D (new_AGEMA_signal_2134), .Q (new_AGEMA_signal_3322) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n9), .Q (new_AGEMA_signal_3324) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (clk), .D (new_AGEMA_signal_1780), .Q (new_AGEMA_signal_3326) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (clk), .D (Midori_rounds_roundReg_out[56]), .Q (new_AGEMA_signal_3328) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (clk), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_3330) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n7), .Q (new_AGEMA_signal_3332) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (clk), .D (new_AGEMA_signal_1778), .Q (new_AGEMA_signal_3334) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (clk), .D (Midori_rounds_roundReg_out[61]), .Q (new_AGEMA_signal_3336) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (clk), .D (new_AGEMA_signal_2139), .Q (new_AGEMA_signal_3338) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n9), .Q (new_AGEMA_signal_3340) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (clk), .D (new_AGEMA_signal_1788), .Q (new_AGEMA_signal_3342) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (clk), .D (Midori_rounds_roundReg_out[60]), .Q (new_AGEMA_signal_3344) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (clk), .D (new_AGEMA_signal_1781), .Q (new_AGEMA_signal_3346) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n7), .Q (new_AGEMA_signal_3348) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (clk), .D (new_AGEMA_signal_1786), .Q (new_AGEMA_signal_3350) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (clk), .D (wk[9]), .Q (new_AGEMA_signal_3352) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (clk), .D (new_AGEMA_signal_1458), .Q (new_AGEMA_signal_3358) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (clk), .D (wk[7]), .Q (new_AGEMA_signal_3364) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (clk), .D (new_AGEMA_signal_1464), .Q (new_AGEMA_signal_3370) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (clk), .D (wk[63]), .Q (new_AGEMA_signal_3376) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (clk), .D (new_AGEMA_signal_1470), .Q (new_AGEMA_signal_3382) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (clk), .D (wk[61]), .Q (new_AGEMA_signal_3388) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (clk), .D (new_AGEMA_signal_1476), .Q (new_AGEMA_signal_3394) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (clk), .D (wk[5]), .Q (new_AGEMA_signal_3400) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (clk), .D (new_AGEMA_signal_1482), .Q (new_AGEMA_signal_3406) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (clk), .D (wk[59]), .Q (new_AGEMA_signal_3412) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (clk), .D (new_AGEMA_signal_1485), .Q (new_AGEMA_signal_3418) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (clk), .D (wk[57]), .Q (new_AGEMA_signal_3424) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_3430) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (clk), .D (wk[55]), .Q (new_AGEMA_signal_3436) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (clk), .D (new_AGEMA_signal_1497), .Q (new_AGEMA_signal_3442) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (clk), .D (wk[53]), .Q (new_AGEMA_signal_3448) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_3454) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (clk), .D (wk[51]), .Q (new_AGEMA_signal_3460) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_3466) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (clk), .D (wk[49]), .Q (new_AGEMA_signal_3472) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (clk), .D (new_AGEMA_signal_1518), .Q (new_AGEMA_signal_3478) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (clk), .D (wk[47]), .Q (new_AGEMA_signal_3484) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (clk), .D (new_AGEMA_signal_1524), .Q (new_AGEMA_signal_3490) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (clk), .D (wk[45]), .Q (new_AGEMA_signal_3496) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (clk), .D (new_AGEMA_signal_1530), .Q (new_AGEMA_signal_3502) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (clk), .D (wk[43]), .Q (new_AGEMA_signal_3508) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (clk), .D (new_AGEMA_signal_1536), .Q (new_AGEMA_signal_3514) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (clk), .D (wk[41]), .Q (new_AGEMA_signal_3520) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (clk), .D (new_AGEMA_signal_1542), .Q (new_AGEMA_signal_3526) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (clk), .D (wk[3]), .Q (new_AGEMA_signal_3532) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (clk), .D (new_AGEMA_signal_1548), .Q (new_AGEMA_signal_3538) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (clk), .D (wk[39]), .Q (new_AGEMA_signal_3544) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (clk), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_3550) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (clk), .D (wk[37]), .Q (new_AGEMA_signal_3556) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (clk), .D (new_AGEMA_signal_1557), .Q (new_AGEMA_signal_3562) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (clk), .D (wk[35]), .Q (new_AGEMA_signal_3568) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (clk), .D (new_AGEMA_signal_1563), .Q (new_AGEMA_signal_3574) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (clk), .D (wk[33]), .Q (new_AGEMA_signal_3580) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (clk), .D (new_AGEMA_signal_1569), .Q (new_AGEMA_signal_3586) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (clk), .D (wk[31]), .Q (new_AGEMA_signal_3592) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (clk), .D (new_AGEMA_signal_1575), .Q (new_AGEMA_signal_3598) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (clk), .D (wk[29]), .Q (new_AGEMA_signal_3604) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (clk), .D (new_AGEMA_signal_1584), .Q (new_AGEMA_signal_3610) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (clk), .D (wk[27]), .Q (new_AGEMA_signal_3616) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (clk), .D (new_AGEMA_signal_1590), .Q (new_AGEMA_signal_3622) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (clk), .D (wk[25]), .Q (new_AGEMA_signal_3628) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (clk), .D (new_AGEMA_signal_1596), .Q (new_AGEMA_signal_3634) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (clk), .D (wk[23]), .Q (new_AGEMA_signal_3640) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (clk), .D (new_AGEMA_signal_1602), .Q (new_AGEMA_signal_3646) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (clk), .D (wk[21]), .Q (new_AGEMA_signal_3652) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (clk), .D (new_AGEMA_signal_1608), .Q (new_AGEMA_signal_3658) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (clk), .D (wk[1]), .Q (new_AGEMA_signal_3664) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (clk), .D (new_AGEMA_signal_1614), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (clk), .D (wk[19]), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (clk), .D (new_AGEMA_signal_1617), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (clk), .D (wk[17]), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (clk), .D (new_AGEMA_signal_1623), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (clk), .D (wk[15]), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (clk), .D (new_AGEMA_signal_1629), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (clk), .D (wk[13]), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (clk), .D (new_AGEMA_signal_1635), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (clk), .D (wk[11]), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (clk), .D (new_AGEMA_signal_1641), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (clk), .D (Midori_rounds_SelectedKey_9_), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (clk), .D (new_AGEMA_signal_1654), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (clk), .D (Midori_rounds_SelectedKey_7_), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (clk), .D (new_AGEMA_signal_2015), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (clk), .D (Midori_rounds_SelectedKey_63_), .Q (new_AGEMA_signal_3760) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (clk), .D (new_AGEMA_signal_2063), .Q (new_AGEMA_signal_3766) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (clk), .D (Midori_rounds_SelectedKey_61_), .Q (new_AGEMA_signal_3772) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (clk), .D (new_AGEMA_signal_2061), .Q (new_AGEMA_signal_3778) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (clk), .D (Midori_rounds_SelectedKey_5_), .Q (new_AGEMA_signal_3784) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (clk), .D (new_AGEMA_signal_2013), .Q (new_AGEMA_signal_3790) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (clk), .D (Midori_rounds_SelectedKey_59_), .Q (new_AGEMA_signal_3796) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (clk), .D (new_AGEMA_signal_2059), .Q (new_AGEMA_signal_3802) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (clk), .D (Midori_rounds_SelectedKey_57_), .Q (new_AGEMA_signal_3808) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (clk), .D (new_AGEMA_signal_2057), .Q (new_AGEMA_signal_3814) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (clk), .D (Midori_rounds_SelectedKey_55_), .Q (new_AGEMA_signal_3820) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (clk), .D (new_AGEMA_signal_2055), .Q (new_AGEMA_signal_3826) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (clk), .D (Midori_rounds_SelectedKey_53_), .Q (new_AGEMA_signal_3832) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_2053), .Q (new_AGEMA_signal_3838) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (clk), .D (Midori_rounds_SelectedKey_51_), .Q (new_AGEMA_signal_3844) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_2051), .Q (new_AGEMA_signal_3850) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (clk), .D (Midori_rounds_SelectedKey_49_), .Q (new_AGEMA_signal_3856) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (new_AGEMA_signal_2049), .Q (new_AGEMA_signal_3862) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (clk), .D (Midori_rounds_SelectedKey_47_), .Q (new_AGEMA_signal_3868) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (clk), .D (new_AGEMA_signal_2047), .Q (new_AGEMA_signal_3874) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (clk), .D (Midori_rounds_SelectedKey_45_), .Q (new_AGEMA_signal_3880) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (clk), .D (new_AGEMA_signal_2045), .Q (new_AGEMA_signal_3886) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (clk), .D (Midori_rounds_SelectedKey_43_), .Q (new_AGEMA_signal_3892) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (clk), .D (new_AGEMA_signal_2043), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (clk), .D (Midori_rounds_SelectedKey_41_), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (clk), .D (new_AGEMA_signal_2041), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (clk), .D (Midori_rounds_SelectedKey_3_), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (clk), .D (new_AGEMA_signal_1651), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (clk), .D (Midori_rounds_SelectedKey_39_), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (clk), .D (new_AGEMA_signal_2039), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (clk), .D (Midori_rounds_SelectedKey_37_), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (clk), .D (new_AGEMA_signal_2037), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (clk), .D (Midori_rounds_SelectedKey_35_), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (clk), .D (new_AGEMA_signal_2035), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (clk), .D (Midori_rounds_SelectedKey_33_), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (clk), .D (new_AGEMA_signal_2033), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (clk), .D (Midori_rounds_SelectedKey_31_), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (clk), .D (new_AGEMA_signal_2031), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (clk), .D (Midori_rounds_SelectedKey_29_), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (clk), .D (new_AGEMA_signal_2029), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (clk), .D (Midori_rounds_SelectedKey_27_), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (clk), .D (new_AGEMA_signal_2027), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (clk), .D (Midori_rounds_SelectedKey_25_), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (clk), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (clk), .D (Midori_rounds_SelectedKey_23_), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (clk), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (clk), .D (Midori_rounds_SelectedKey_21_), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (clk), .D (new_AGEMA_signal_2022), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (clk), .D (Midori_rounds_SelectedKey_1_), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (clk), .D (new_AGEMA_signal_1649), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (clk), .D (Midori_rounds_SelectedKey_19_), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (clk), .D (new_AGEMA_signal_2020), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (clk), .D (Midori_rounds_SelectedKey_17_), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (clk), .D (new_AGEMA_signal_2018), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (clk), .D (Midori_rounds_SelectedKey_15_), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (clk), .D (new_AGEMA_signal_1659), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (clk), .D (Midori_rounds_SelectedKey_13_), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (clk), .D (new_AGEMA_signal_1657), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (clk), .D (Midori_rounds_SelectedKey_11_), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (clk), .D (new_AGEMA_signal_1656), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (clk), .D (Midori_add_Result_Start[1]), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_1894), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (clk), .D (Midori_add_Result_Start[3]), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_1850), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (clk), .D (Midori_add_Result_Start[5]), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_1806), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (clk), .D (Midori_add_Result_Start[7]), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_1794), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (clk), .D (Midori_add_Result_Start[9]), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_1790), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (clk), .D (Midori_add_Result_Start[11]), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (clk), .D (Midori_add_Result_Start[13]), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (clk), .D (Midori_add_Result_Start[15]), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_1904), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (clk), .D (Midori_add_Result_Start[17]), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_1900), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (clk), .D (Midori_add_Result_Start[19]), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (clk), .D (Midori_add_Result_Start[21]), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_1890), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (clk), .D (Midori_add_Result_Start[23]), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_1886), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (clk), .D (Midori_add_Result_Start[25]), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (clk), .D (Midori_add_Result_Start[27]), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_1878), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (clk), .D (Midori_add_Result_Start[29]), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_1874), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (clk), .D (Midori_add_Result_Start[31]), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_1868), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (clk), .D (Midori_add_Result_Start[33]), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_1864), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (clk), .D (Midori_add_Result_Start[35]), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_1860), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (clk), .D (Midori_add_Result_Start[37]), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (clk), .D (Midori_add_Result_Start[39]), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (clk), .D (Midori_add_Result_Start[41]), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_4372) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (clk), .D (Midori_add_Result_Start[43]), .Q (new_AGEMA_signal_4378) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_1842), .Q (new_AGEMA_signal_4384) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (clk), .D (Midori_add_Result_Start[45]), .Q (new_AGEMA_signal_4390) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_4396) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (clk), .D (Midori_add_Result_Start[47]), .Q (new_AGEMA_signal_4402) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_1834), .Q (new_AGEMA_signal_4408) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (clk), .D (Midori_add_Result_Start[49]), .Q (new_AGEMA_signal_4414) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_1830), .Q (new_AGEMA_signal_4420) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (clk), .D (Midori_add_Result_Start[51]), .Q (new_AGEMA_signal_4426) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_1824), .Q (new_AGEMA_signal_4432) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (clk), .D (Midori_add_Result_Start[53]), .Q (new_AGEMA_signal_4438) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_4444) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (clk), .D (Midori_add_Result_Start[55]), .Q (new_AGEMA_signal_4450) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_1816), .Q (new_AGEMA_signal_4456) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (clk), .D (Midori_add_Result_Start[57]), .Q (new_AGEMA_signal_4462) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_1812), .Q (new_AGEMA_signal_4468) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (clk), .D (Midori_add_Result_Start[59]), .Q (new_AGEMA_signal_4474) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_1808), .Q (new_AGEMA_signal_4480) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (clk), .D (Midori_add_Result_Start[61]), .Q (new_AGEMA_signal_4486) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_4492) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (clk), .D (Midori_add_Result_Start[63]), .Q (new_AGEMA_signal_4498) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_1798), .Q (new_AGEMA_signal_4504) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C (clk), .D (enc_dec), .Q (new_AGEMA_signal_4702) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C (clk), .D (wk[8]), .Q (new_AGEMA_signal_4708) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_1461), .Q (new_AGEMA_signal_4716) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C (clk), .D (wk[6]), .Q (new_AGEMA_signal_4724) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_1467), .Q (new_AGEMA_signal_4732) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C (clk), .D (wk[62]), .Q (new_AGEMA_signal_4740) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_1473), .Q (new_AGEMA_signal_4748) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C (clk), .D (wk[60]), .Q (new_AGEMA_signal_4756) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_1479), .Q (new_AGEMA_signal_4764) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C (clk), .D (wk[58]), .Q (new_AGEMA_signal_4772) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_1488), .Q (new_AGEMA_signal_4780) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C (clk), .D (wk[56]), .Q (new_AGEMA_signal_4788) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_1494), .Q (new_AGEMA_signal_4796) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C (clk), .D (wk[54]), .Q (new_AGEMA_signal_4804) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_1500), .Q (new_AGEMA_signal_4812) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C (clk), .D (wk[52]), .Q (new_AGEMA_signal_4820) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_1506), .Q (new_AGEMA_signal_4828) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C (clk), .D (wk[50]), .Q (new_AGEMA_signal_4836) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_4844) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C (clk), .D (wk[4]), .Q (new_AGEMA_signal_4852) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_1515), .Q (new_AGEMA_signal_4860) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C (clk), .D (wk[48]), .Q (new_AGEMA_signal_4868) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_1521), .Q (new_AGEMA_signal_4876) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C (clk), .D (wk[46]), .Q (new_AGEMA_signal_4884) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_1527), .Q (new_AGEMA_signal_4892) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C (clk), .D (wk[44]), .Q (new_AGEMA_signal_4900) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_1533), .Q (new_AGEMA_signal_4908) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C (clk), .D (wk[42]), .Q (new_AGEMA_signal_4916) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_1539), .Q (new_AGEMA_signal_4924) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C (clk), .D (wk[40]), .Q (new_AGEMA_signal_4932) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_1545), .Q (new_AGEMA_signal_4940) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C (clk), .D (wk[38]), .Q (new_AGEMA_signal_4948) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_1554), .Q (new_AGEMA_signal_4956) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C (clk), .D (wk[36]), .Q (new_AGEMA_signal_4964) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_1560), .Q (new_AGEMA_signal_4972) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C (clk), .D (wk[34]), .Q (new_AGEMA_signal_4980) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_1566), .Q (new_AGEMA_signal_4988) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C (clk), .D (wk[32]), .Q (new_AGEMA_signal_4996) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_1572), .Q (new_AGEMA_signal_5004) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C (clk), .D (wk[30]), .Q (new_AGEMA_signal_5012) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_1578), .Q (new_AGEMA_signal_5020) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C (clk), .D (wk[2]), .Q (new_AGEMA_signal_5028) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_1581), .Q (new_AGEMA_signal_5036) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C (clk), .D (wk[28]), .Q (new_AGEMA_signal_5044) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_1587), .Q (new_AGEMA_signal_5052) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C (clk), .D (wk[26]), .Q (new_AGEMA_signal_5060) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_1593), .Q (new_AGEMA_signal_5068) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C (clk), .D (wk[24]), .Q (new_AGEMA_signal_5076) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_1599), .Q (new_AGEMA_signal_5084) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C (clk), .D (wk[22]), .Q (new_AGEMA_signal_5092) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_1605), .Q (new_AGEMA_signal_5100) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C (clk), .D (wk[20]), .Q (new_AGEMA_signal_5108) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_1611), .Q (new_AGEMA_signal_5116) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C (clk), .D (wk[18]), .Q (new_AGEMA_signal_5124) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_1620), .Q (new_AGEMA_signal_5132) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C (clk), .D (wk[16]), .Q (new_AGEMA_signal_5140) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_1626), .Q (new_AGEMA_signal_5148) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C (clk), .D (wk[14]), .Q (new_AGEMA_signal_5156) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_1632), .Q (new_AGEMA_signal_5164) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C (clk), .D (wk[12]), .Q (new_AGEMA_signal_5172) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_1638), .Q (new_AGEMA_signal_5180) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C (clk), .D (wk[10]), .Q (new_AGEMA_signal_5188) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_1644), .Q (new_AGEMA_signal_5196) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C (clk), .D (wk[0]), .Q (new_AGEMA_signal_5204) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_1647), .Q (new_AGEMA_signal_5212) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C (clk), .D (Midori_rounds_n16), .Q (new_AGEMA_signal_5220) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_5228) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C (clk), .D (Midori_rounds_SelectedKey_6_), .Q (new_AGEMA_signal_5236) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_2014), .Q (new_AGEMA_signal_5244) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C (clk), .D (Midori_rounds_SelectedKey_62_), .Q (new_AGEMA_signal_5252) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_2062), .Q (new_AGEMA_signal_5260) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C (clk), .D (Midori_rounds_n15), .Q (new_AGEMA_signal_5268) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_5276) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C (clk), .D (Midori_rounds_SelectedKey_58_), .Q (new_AGEMA_signal_5284) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_2058), .Q (new_AGEMA_signal_5292) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C (clk), .D (Midori_rounds_n14), .Q (new_AGEMA_signal_5300) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_2497), .Q (new_AGEMA_signal_5308) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C (clk), .D (Midori_rounds_SelectedKey_54_), .Q (new_AGEMA_signal_5316) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_2054), .Q (new_AGEMA_signal_5324) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C (clk), .D (Midori_rounds_n13), .Q (new_AGEMA_signal_5332) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_2498), .Q (new_AGEMA_signal_5340) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C (clk), .D (Midori_rounds_SelectedKey_50_), .Q (new_AGEMA_signal_5348) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_2050), .Q (new_AGEMA_signal_5356) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C (clk), .D (Midori_rounds_n12), .Q (new_AGEMA_signal_5364) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_2499), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C (clk), .D (Midori_rounds_n11), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_5388) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C (clk), .D (Midori_rounds_SelectedKey_46_), .Q (new_AGEMA_signal_5396) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_2046), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C (clk), .D (Midori_rounds_n10), .Q (new_AGEMA_signal_5412) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_2460), .Q (new_AGEMA_signal_5420) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C (clk), .D (Midori_rounds_SelectedKey_42_), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_2042), .Q (new_AGEMA_signal_5436) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C (clk), .D (Midori_rounds_n9), .Q (new_AGEMA_signal_5444) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_2500), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C (clk), .D (Midori_rounds_SelectedKey_38_), .Q (new_AGEMA_signal_5460) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_2038), .Q (new_AGEMA_signal_5468) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C (clk), .D (Midori_rounds_n8), .Q (new_AGEMA_signal_5476) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_5484) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C (clk), .D (Midori_rounds_SelectedKey_34_), .Q (new_AGEMA_signal_5492) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_2034), .Q (new_AGEMA_signal_5500) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C (clk), .D (Midori_rounds_n7), .Q (new_AGEMA_signal_5508) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_2501), .Q (new_AGEMA_signal_5516) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C (clk), .D (Midori_rounds_SelectedKey_30_), .Q (new_AGEMA_signal_5524) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_2030), .Q (new_AGEMA_signal_5532) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C (clk), .D (Midori_rounds_SelectedKey_2_), .Q (new_AGEMA_signal_5540) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_1650), .Q (new_AGEMA_signal_5548) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C (clk), .D (Midori_rounds_n6), .Q (new_AGEMA_signal_5556) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_2564), .Q (new_AGEMA_signal_5564) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C (clk), .D (Midori_rounds_SelectedKey_26_), .Q (new_AGEMA_signal_5572) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_1660), .Q (new_AGEMA_signal_5580) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C (clk), .D (Midori_rounds_n5), .Q (new_AGEMA_signal_5588) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_2502), .Q (new_AGEMA_signal_5596) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C (clk), .D (Midori_rounds_SelectedKey_22_), .Q (new_AGEMA_signal_5604) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_2023), .Q (new_AGEMA_signal_5612) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C (clk), .D (Midori_rounds_n4), .Q (new_AGEMA_signal_5620) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_2482), .Q (new_AGEMA_signal_5628) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C (clk), .D (Midori_rounds_SelectedKey_18_), .Q (new_AGEMA_signal_5636) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_2019), .Q (new_AGEMA_signal_5644) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C (clk), .D (Midori_rounds_n3), .Q (new_AGEMA_signal_5652) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_2503), .Q (new_AGEMA_signal_5660) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C (clk), .D (Midori_rounds_SelectedKey_14_), .Q (new_AGEMA_signal_5668) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_5676) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C (clk), .D (Midori_rounds_n2), .Q (new_AGEMA_signal_5684) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_2504), .Q (new_AGEMA_signal_5692) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C (clk), .D (Midori_rounds_SelectedKey_10_), .Q (new_AGEMA_signal_5700) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_1655), .Q (new_AGEMA_signal_5708) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C (clk), .D (Midori_rounds_n1), .Q (new_AGEMA_signal_5716) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_2505), .Q (new_AGEMA_signal_5724) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C (clk), .D (Midori_add_Result_Start[0]), .Q (new_AGEMA_signal_5734) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C (clk), .D (new_AGEMA_signal_1916), .Q (new_AGEMA_signal_5742) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C (clk), .D (Midori_add_Result_Start[2]), .Q (new_AGEMA_signal_5750) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C (clk), .D (new_AGEMA_signal_1872), .Q (new_AGEMA_signal_5758) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C (clk), .D (Midori_add_Result_Start[4]), .Q (new_AGEMA_signal_5766) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C (clk), .D (new_AGEMA_signal_1828), .Q (new_AGEMA_signal_5774) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C (clk), .D (Midori_add_Result_Start[6]), .Q (new_AGEMA_signal_5782) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C (clk), .D (new_AGEMA_signal_1796), .Q (new_AGEMA_signal_5790) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C (clk), .D (Midori_add_Result_Start[8]), .Q (new_AGEMA_signal_5798) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C (clk), .D (new_AGEMA_signal_1792), .Q (new_AGEMA_signal_5806) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C (clk), .D (Midori_add_Result_Start[10]), .Q (new_AGEMA_signal_5814) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C (clk), .D (new_AGEMA_signal_1914), .Q (new_AGEMA_signal_5822) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C (clk), .D (Midori_add_Result_Start[12]), .Q (new_AGEMA_signal_5830) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_5838) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C (clk), .D (Midori_add_Result_Start[14]), .Q (new_AGEMA_signal_5846) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C (clk), .D (new_AGEMA_signal_1906), .Q (new_AGEMA_signal_5854) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C (clk), .D (Midori_add_Result_Start[16]), .Q (new_AGEMA_signal_5862) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C (clk), .D (new_AGEMA_signal_1902), .Q (new_AGEMA_signal_5870) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C (clk), .D (Midori_add_Result_Start[18]), .Q (new_AGEMA_signal_5878) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_5886) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C (clk), .D (Midori_add_Result_Start[20]), .Q (new_AGEMA_signal_5894) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_5902) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C (clk), .D (Midori_add_Result_Start[22]), .Q (new_AGEMA_signal_5910) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_1888), .Q (new_AGEMA_signal_5918) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C (clk), .D (Midori_add_Result_Start[24]), .Q (new_AGEMA_signal_5926) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C (clk), .D (new_AGEMA_signal_1884), .Q (new_AGEMA_signal_5934) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C (clk), .D (Midori_add_Result_Start[26]), .Q (new_AGEMA_signal_5942) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C (clk), .D (new_AGEMA_signal_1880), .Q (new_AGEMA_signal_5950) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C (clk), .D (Midori_add_Result_Start[28]), .Q (new_AGEMA_signal_5958) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_1876), .Q (new_AGEMA_signal_5966) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C (clk), .D (Midori_add_Result_Start[30]), .Q (new_AGEMA_signal_5974) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_1870), .Q (new_AGEMA_signal_5982) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C (clk), .D (Midori_add_Result_Start[32]), .Q (new_AGEMA_signal_5990) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C (clk), .D (new_AGEMA_signal_1866), .Q (new_AGEMA_signal_5998) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C (clk), .D (Midori_add_Result_Start[34]), .Q (new_AGEMA_signal_6006) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_1862), .Q (new_AGEMA_signal_6014) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C (clk), .D (Midori_add_Result_Start[36]), .Q (new_AGEMA_signal_6022) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_6030) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C (clk), .D (Midori_add_Result_Start[38]), .Q (new_AGEMA_signal_6038) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_6046) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C (clk), .D (Midori_add_Result_Start[40]), .Q (new_AGEMA_signal_6054) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C (clk), .D (new_AGEMA_signal_1848), .Q (new_AGEMA_signal_6062) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C (clk), .D (Midori_add_Result_Start[42]), .Q (new_AGEMA_signal_6070) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_6078) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C (clk), .D (Midori_add_Result_Start[44]), .Q (new_AGEMA_signal_6086) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C (clk), .D (new_AGEMA_signal_1840), .Q (new_AGEMA_signal_6094) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C (clk), .D (Midori_add_Result_Start[46]), .Q (new_AGEMA_signal_6102) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C (clk), .D (new_AGEMA_signal_1836), .Q (new_AGEMA_signal_6110) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C (clk), .D (Midori_add_Result_Start[48]), .Q (new_AGEMA_signal_6118) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_6126) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C (clk), .D (Midori_add_Result_Start[50]), .Q (new_AGEMA_signal_6134) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C (clk), .D (new_AGEMA_signal_1826), .Q (new_AGEMA_signal_6142) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C (clk), .D (Midori_add_Result_Start[52]), .Q (new_AGEMA_signal_6150) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C (clk), .D (new_AGEMA_signal_1822), .Q (new_AGEMA_signal_6158) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C (clk), .D (Midori_add_Result_Start[54]), .Q (new_AGEMA_signal_6166) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C (clk), .D (new_AGEMA_signal_1818), .Q (new_AGEMA_signal_6174) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C (clk), .D (Midori_add_Result_Start[56]), .Q (new_AGEMA_signal_6182) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C (clk), .D (new_AGEMA_signal_1814), .Q (new_AGEMA_signal_6190) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C (clk), .D (Midori_add_Result_Start[58]), .Q (new_AGEMA_signal_6198) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C (clk), .D (new_AGEMA_signal_1810), .Q (new_AGEMA_signal_6206) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C (clk), .D (Midori_add_Result_Start[60]), .Q (new_AGEMA_signal_6214) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C (clk), .D (new_AGEMA_signal_1804), .Q (new_AGEMA_signal_6222) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C (clk), .D (Midori_add_Result_Start[62]), .Q (new_AGEMA_signal_6230) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C (clk), .D (new_AGEMA_signal_1800), .Q (new_AGEMA_signal_6238) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C (clk), .D (controller_roundCounter_N7), .Q (new_AGEMA_signal_6440) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C (clk), .D (controller_roundCounter_N8), .Q (new_AGEMA_signal_6448) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C (clk), .D (controller_roundCounter_n2), .Q (new_AGEMA_signal_6456) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C (clk), .D (controller_roundCounter_N10), .Q (new_AGEMA_signal_6464) ) ;

    /* cells in depth 2 */
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .a ({new_AGEMA_signal_1661, Midori_rounds_roundReg_out[0]}), .b ({new_AGEMA_signal_1662, Midori_rounds_roundReg_out[3]}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_1663, Midori_rounds_sub_sBox_PRINCE_0_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .a ({new_AGEMA_signal_1667, Midori_rounds_sub_sBox_PRINCE_0_n8}), .b ({new_AGEMA_signal_1666, Midori_rounds_sub_sBox_PRINCE_0_n7}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_1918, Midori_rounds_sub_sBox_PRINCE_0_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .a ({new_AGEMA_signal_1662, Midori_rounds_roundReg_out[3]}), .b ({new_AGEMA_signal_1668, Midori_rounds_sub_sBox_PRINCE_0_n9}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_1919, Midori_rounds_sub_sBox_PRINCE_0_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .a ({new_AGEMA_signal_1664, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1667, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_1920, Midori_rounds_sub_sBox_PRINCE_0_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .a ({new_AGEMA_signal_1664, Midori_rounds_roundReg_out[2]}), .b ({new_AGEMA_signal_1662, Midori_rounds_roundReg_out[3]}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_1665, Midori_rounds_sub_sBox_PRINCE_0_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .a ({new_AGEMA_signal_1668, Midori_rounds_sub_sBox_PRINCE_0_n9}), .b ({new_AGEMA_signal_1667, Midori_rounds_sub_sBox_PRINCE_0_n8}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_0_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .a ({new_AGEMA_signal_1669, Midori_rounds_roundReg_out[4]}), .b ({new_AGEMA_signal_1670, Midori_rounds_roundReg_out[7]}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_1671, Midori_rounds_sub_sBox_PRINCE_1_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .a ({new_AGEMA_signal_1675, Midori_rounds_sub_sBox_PRINCE_1_n8}), .b ({new_AGEMA_signal_1674, Midori_rounds_sub_sBox_PRINCE_1_n7}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_1924, Midori_rounds_sub_sBox_PRINCE_1_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .a ({new_AGEMA_signal_1670, Midori_rounds_roundReg_out[7]}), .b ({new_AGEMA_signal_1676, Midori_rounds_sub_sBox_PRINCE_1_n9}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_1925, Midori_rounds_sub_sBox_PRINCE_1_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .a ({new_AGEMA_signal_1672, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1675, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_1926, Midori_rounds_sub_sBox_PRINCE_1_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U5 ( .a ({new_AGEMA_signal_1672, Midori_rounds_roundReg_out[6]}), .b ({new_AGEMA_signal_1670, Midori_rounds_roundReg_out[7]}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_1673, Midori_rounds_sub_sBox_PRINCE_1_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U3 ( .a ({new_AGEMA_signal_1676, Midori_rounds_sub_sBox_PRINCE_1_n9}), .b ({new_AGEMA_signal_1675, Midori_rounds_sub_sBox_PRINCE_1_n8}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_1_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .a ({new_AGEMA_signal_1677, Midori_rounds_roundReg_out[8]}), .b ({new_AGEMA_signal_1678, Midori_rounds_roundReg_out[11]}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_1679, Midori_rounds_sub_sBox_PRINCE_2_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .a ({new_AGEMA_signal_1683, Midori_rounds_sub_sBox_PRINCE_2_n8}), .b ({new_AGEMA_signal_1682, Midori_rounds_sub_sBox_PRINCE_2_n7}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_1930, Midori_rounds_sub_sBox_PRINCE_2_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .a ({new_AGEMA_signal_1678, Midori_rounds_roundReg_out[11]}), .b ({new_AGEMA_signal_1684, Midori_rounds_sub_sBox_PRINCE_2_n9}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_1931, Midori_rounds_sub_sBox_PRINCE_2_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .a ({new_AGEMA_signal_1680, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1683, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_1932, Midori_rounds_sub_sBox_PRINCE_2_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U5 ( .a ({new_AGEMA_signal_1680, Midori_rounds_roundReg_out[10]}), .b ({new_AGEMA_signal_1678, Midori_rounds_roundReg_out[11]}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_1681, Midori_rounds_sub_sBox_PRINCE_2_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U3 ( .a ({new_AGEMA_signal_1684, Midori_rounds_sub_sBox_PRINCE_2_n9}), .b ({new_AGEMA_signal_1683, Midori_rounds_sub_sBox_PRINCE_2_n8}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_2_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .a ({new_AGEMA_signal_1685, Midori_rounds_roundReg_out[12]}), .b ({new_AGEMA_signal_1686, Midori_rounds_roundReg_out[15]}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_1687, Midori_rounds_sub_sBox_PRINCE_3_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .a ({new_AGEMA_signal_1691, Midori_rounds_sub_sBox_PRINCE_3_n8}), .b ({new_AGEMA_signal_1690, Midori_rounds_sub_sBox_PRINCE_3_n7}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_1936, Midori_rounds_sub_sBox_PRINCE_3_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .a ({new_AGEMA_signal_1686, Midori_rounds_roundReg_out[15]}), .b ({new_AGEMA_signal_1692, Midori_rounds_sub_sBox_PRINCE_3_n9}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_1937, Midori_rounds_sub_sBox_PRINCE_3_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .a ({new_AGEMA_signal_1688, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1691, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_1938, Midori_rounds_sub_sBox_PRINCE_3_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U5 ( .a ({new_AGEMA_signal_1688, Midori_rounds_roundReg_out[14]}), .b ({new_AGEMA_signal_1686, Midori_rounds_roundReg_out[15]}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_1689, Midori_rounds_sub_sBox_PRINCE_3_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U3 ( .a ({new_AGEMA_signal_1692, Midori_rounds_sub_sBox_PRINCE_3_n9}), .b ({new_AGEMA_signal_1691, Midori_rounds_sub_sBox_PRINCE_3_n8}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_3_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .a ({new_AGEMA_signal_1693, Midori_rounds_roundReg_out[16]}), .b ({new_AGEMA_signal_1694, Midori_rounds_roundReg_out[19]}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_1695, Midori_rounds_sub_sBox_PRINCE_4_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .a ({new_AGEMA_signal_1699, Midori_rounds_sub_sBox_PRINCE_4_n8}), .b ({new_AGEMA_signal_1698, Midori_rounds_sub_sBox_PRINCE_4_n7}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_1942, Midori_rounds_sub_sBox_PRINCE_4_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .a ({new_AGEMA_signal_1694, Midori_rounds_roundReg_out[19]}), .b ({new_AGEMA_signal_1700, Midori_rounds_sub_sBox_PRINCE_4_n9}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_1943, Midori_rounds_sub_sBox_PRINCE_4_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .a ({new_AGEMA_signal_1696, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1699, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_1944, Midori_rounds_sub_sBox_PRINCE_4_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U5 ( .a ({new_AGEMA_signal_1696, Midori_rounds_roundReg_out[18]}), .b ({new_AGEMA_signal_1694, Midori_rounds_roundReg_out[19]}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_1697, Midori_rounds_sub_sBox_PRINCE_4_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U3 ( .a ({new_AGEMA_signal_1700, Midori_rounds_sub_sBox_PRINCE_4_n9}), .b ({new_AGEMA_signal_1699, Midori_rounds_sub_sBox_PRINCE_4_n8}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_1946, Midori_rounds_sub_sBox_PRINCE_4_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .a ({new_AGEMA_signal_1701, Midori_rounds_roundReg_out[20]}), .b ({new_AGEMA_signal_1702, Midori_rounds_roundReg_out[23]}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_1703, Midori_rounds_sub_sBox_PRINCE_5_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .a ({new_AGEMA_signal_1707, Midori_rounds_sub_sBox_PRINCE_5_n8}), .b ({new_AGEMA_signal_1706, Midori_rounds_sub_sBox_PRINCE_5_n7}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_1948, Midori_rounds_sub_sBox_PRINCE_5_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .a ({new_AGEMA_signal_1702, Midori_rounds_roundReg_out[23]}), .b ({new_AGEMA_signal_1708, Midori_rounds_sub_sBox_PRINCE_5_n9}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_1949, Midori_rounds_sub_sBox_PRINCE_5_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .a ({new_AGEMA_signal_1704, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1707, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_1950, Midori_rounds_sub_sBox_PRINCE_5_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U5 ( .a ({new_AGEMA_signal_1704, Midori_rounds_roundReg_out[22]}), .b ({new_AGEMA_signal_1702, Midori_rounds_roundReg_out[23]}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_1705, Midori_rounds_sub_sBox_PRINCE_5_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U3 ( .a ({new_AGEMA_signal_1708, Midori_rounds_sub_sBox_PRINCE_5_n9}), .b ({new_AGEMA_signal_1707, Midori_rounds_sub_sBox_PRINCE_5_n8}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_1952, Midori_rounds_sub_sBox_PRINCE_5_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .a ({new_AGEMA_signal_1709, Midori_rounds_roundReg_out[24]}), .b ({new_AGEMA_signal_1710, Midori_rounds_roundReg_out[27]}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_1711, Midori_rounds_sub_sBox_PRINCE_6_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .a ({new_AGEMA_signal_1715, Midori_rounds_sub_sBox_PRINCE_6_n8}), .b ({new_AGEMA_signal_1714, Midori_rounds_sub_sBox_PRINCE_6_n7}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_1954, Midori_rounds_sub_sBox_PRINCE_6_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .a ({new_AGEMA_signal_1710, Midori_rounds_roundReg_out[27]}), .b ({new_AGEMA_signal_1716, Midori_rounds_sub_sBox_PRINCE_6_n9}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_1955, Midori_rounds_sub_sBox_PRINCE_6_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .a ({new_AGEMA_signal_1712, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1715, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_1956, Midori_rounds_sub_sBox_PRINCE_6_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U5 ( .a ({new_AGEMA_signal_1712, Midori_rounds_roundReg_out[26]}), .b ({new_AGEMA_signal_1710, Midori_rounds_roundReg_out[27]}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_1713, Midori_rounds_sub_sBox_PRINCE_6_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U3 ( .a ({new_AGEMA_signal_1716, Midori_rounds_sub_sBox_PRINCE_6_n9}), .b ({new_AGEMA_signal_1715, Midori_rounds_sub_sBox_PRINCE_6_n8}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_6_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .a ({new_AGEMA_signal_1717, Midori_rounds_roundReg_out[28]}), .b ({new_AGEMA_signal_1718, Midori_rounds_roundReg_out[31]}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_1719, Midori_rounds_sub_sBox_PRINCE_7_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .a ({new_AGEMA_signal_1723, Midori_rounds_sub_sBox_PRINCE_7_n8}), .b ({new_AGEMA_signal_1722, Midori_rounds_sub_sBox_PRINCE_7_n7}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_1960, Midori_rounds_sub_sBox_PRINCE_7_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .a ({new_AGEMA_signal_1718, Midori_rounds_roundReg_out[31]}), .b ({new_AGEMA_signal_1724, Midori_rounds_sub_sBox_PRINCE_7_n9}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_1961, Midori_rounds_sub_sBox_PRINCE_7_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .a ({new_AGEMA_signal_1720, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1723, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_1962, Midori_rounds_sub_sBox_PRINCE_7_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .a ({new_AGEMA_signal_1720, Midori_rounds_roundReg_out[30]}), .b ({new_AGEMA_signal_1718, Midori_rounds_roundReg_out[31]}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_1721, Midori_rounds_sub_sBox_PRINCE_7_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .a ({new_AGEMA_signal_1724, Midori_rounds_sub_sBox_PRINCE_7_n9}), .b ({new_AGEMA_signal_1723, Midori_rounds_sub_sBox_PRINCE_7_n8}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_1964, Midori_rounds_sub_sBox_PRINCE_7_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .a ({new_AGEMA_signal_1725, Midori_rounds_roundReg_out[32]}), .b ({new_AGEMA_signal_1726, Midori_rounds_roundReg_out[35]}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_1727, Midori_rounds_sub_sBox_PRINCE_8_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .a ({new_AGEMA_signal_1731, Midori_rounds_sub_sBox_PRINCE_8_n8}), .b ({new_AGEMA_signal_1730, Midori_rounds_sub_sBox_PRINCE_8_n7}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_1966, Midori_rounds_sub_sBox_PRINCE_8_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .a ({new_AGEMA_signal_1726, Midori_rounds_roundReg_out[35]}), .b ({new_AGEMA_signal_1732, Midori_rounds_sub_sBox_PRINCE_8_n9}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_1967, Midori_rounds_sub_sBox_PRINCE_8_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .a ({new_AGEMA_signal_1728, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_1731, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_1968, Midori_rounds_sub_sBox_PRINCE_8_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .a ({new_AGEMA_signal_1728, Midori_rounds_roundReg_out[34]}), .b ({new_AGEMA_signal_1726, Midori_rounds_roundReg_out[35]}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_1729, Midori_rounds_sub_sBox_PRINCE_8_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .a ({new_AGEMA_signal_1732, Midori_rounds_sub_sBox_PRINCE_8_n9}), .b ({new_AGEMA_signal_1731, Midori_rounds_sub_sBox_PRINCE_8_n8}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_8_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .a ({new_AGEMA_signal_1733, Midori_rounds_roundReg_out[36]}), .b ({new_AGEMA_signal_1734, Midori_rounds_roundReg_out[39]}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_1735, Midori_rounds_sub_sBox_PRINCE_9_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .a ({new_AGEMA_signal_1739, Midori_rounds_sub_sBox_PRINCE_9_n8}), .b ({new_AGEMA_signal_1738, Midori_rounds_sub_sBox_PRINCE_9_n7}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_1972, Midori_rounds_sub_sBox_PRINCE_9_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .a ({new_AGEMA_signal_1734, Midori_rounds_roundReg_out[39]}), .b ({new_AGEMA_signal_1740, Midori_rounds_sub_sBox_PRINCE_9_n9}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_1973, Midori_rounds_sub_sBox_PRINCE_9_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .a ({new_AGEMA_signal_1736, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_1739, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_1974, Midori_rounds_sub_sBox_PRINCE_9_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .a ({new_AGEMA_signal_1736, Midori_rounds_roundReg_out[38]}), .b ({new_AGEMA_signal_1734, Midori_rounds_roundReg_out[39]}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_1737, Midori_rounds_sub_sBox_PRINCE_9_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .a ({new_AGEMA_signal_1740, Midori_rounds_sub_sBox_PRINCE_9_n9}), .b ({new_AGEMA_signal_1739, Midori_rounds_sub_sBox_PRINCE_9_n8}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_9_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .a ({new_AGEMA_signal_1741, Midori_rounds_roundReg_out[40]}), .b ({new_AGEMA_signal_1742, Midori_rounds_roundReg_out[43]}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_1743, Midori_rounds_sub_sBox_PRINCE_10_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .a ({new_AGEMA_signal_1747, Midori_rounds_sub_sBox_PRINCE_10_n8}), .b ({new_AGEMA_signal_1746, Midori_rounds_sub_sBox_PRINCE_10_n7}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_1978, Midori_rounds_sub_sBox_PRINCE_10_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .a ({new_AGEMA_signal_1742, Midori_rounds_roundReg_out[43]}), .b ({new_AGEMA_signal_1748, Midori_rounds_sub_sBox_PRINCE_10_n9}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_1979, Midori_rounds_sub_sBox_PRINCE_10_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .a ({new_AGEMA_signal_1744, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_1747, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_1980, Midori_rounds_sub_sBox_PRINCE_10_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U5 ( .a ({new_AGEMA_signal_1744, Midori_rounds_roundReg_out[42]}), .b ({new_AGEMA_signal_1742, Midori_rounds_roundReg_out[43]}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_1745, Midori_rounds_sub_sBox_PRINCE_10_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U3 ( .a ({new_AGEMA_signal_1748, Midori_rounds_sub_sBox_PRINCE_10_n9}), .b ({new_AGEMA_signal_1747, Midori_rounds_sub_sBox_PRINCE_10_n8}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_10_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .a ({new_AGEMA_signal_1749, Midori_rounds_roundReg_out[44]}), .b ({new_AGEMA_signal_1750, Midori_rounds_roundReg_out[47]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_1751, Midori_rounds_sub_sBox_PRINCE_11_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .a ({new_AGEMA_signal_1755, Midori_rounds_sub_sBox_PRINCE_11_n8}), .b ({new_AGEMA_signal_1754, Midori_rounds_sub_sBox_PRINCE_11_n7}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_1984, Midori_rounds_sub_sBox_PRINCE_11_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .a ({new_AGEMA_signal_1750, Midori_rounds_roundReg_out[47]}), .b ({new_AGEMA_signal_1756, Midori_rounds_sub_sBox_PRINCE_11_n9}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_1985, Midori_rounds_sub_sBox_PRINCE_11_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .a ({new_AGEMA_signal_1752, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_1755, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_1986, Midori_rounds_sub_sBox_PRINCE_11_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U5 ( .a ({new_AGEMA_signal_1752, Midori_rounds_roundReg_out[46]}), .b ({new_AGEMA_signal_1750, Midori_rounds_roundReg_out[47]}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_1753, Midori_rounds_sub_sBox_PRINCE_11_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U3 ( .a ({new_AGEMA_signal_1756, Midori_rounds_sub_sBox_PRINCE_11_n9}), .b ({new_AGEMA_signal_1755, Midori_rounds_sub_sBox_PRINCE_11_n8}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_11_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .a ({new_AGEMA_signal_1757, Midori_rounds_roundReg_out[48]}), .b ({new_AGEMA_signal_1758, Midori_rounds_roundReg_out[51]}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_1759, Midori_rounds_sub_sBox_PRINCE_12_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .a ({new_AGEMA_signal_1763, Midori_rounds_sub_sBox_PRINCE_12_n8}), .b ({new_AGEMA_signal_1762, Midori_rounds_sub_sBox_PRINCE_12_n7}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_1990, Midori_rounds_sub_sBox_PRINCE_12_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .a ({new_AGEMA_signal_1758, Midori_rounds_roundReg_out[51]}), .b ({new_AGEMA_signal_1764, Midori_rounds_sub_sBox_PRINCE_12_n9}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_1991, Midori_rounds_sub_sBox_PRINCE_12_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .a ({new_AGEMA_signal_1760, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_1763, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_1992, Midori_rounds_sub_sBox_PRINCE_12_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U5 ( .a ({new_AGEMA_signal_1760, Midori_rounds_roundReg_out[50]}), .b ({new_AGEMA_signal_1758, Midori_rounds_roundReg_out[51]}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_1761, Midori_rounds_sub_sBox_PRINCE_12_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U3 ( .a ({new_AGEMA_signal_1764, Midori_rounds_sub_sBox_PRINCE_12_n9}), .b ({new_AGEMA_signal_1763, Midori_rounds_sub_sBox_PRINCE_12_n8}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_1994, Midori_rounds_sub_sBox_PRINCE_12_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .a ({new_AGEMA_signal_1765, Midori_rounds_roundReg_out[52]}), .b ({new_AGEMA_signal_1766, Midori_rounds_roundReg_out[55]}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_1767, Midori_rounds_sub_sBox_PRINCE_13_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .a ({new_AGEMA_signal_1771, Midori_rounds_sub_sBox_PRINCE_13_n8}), .b ({new_AGEMA_signal_1770, Midori_rounds_sub_sBox_PRINCE_13_n7}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_1996, Midori_rounds_sub_sBox_PRINCE_13_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .a ({new_AGEMA_signal_1766, Midori_rounds_roundReg_out[55]}), .b ({new_AGEMA_signal_1772, Midori_rounds_sub_sBox_PRINCE_13_n9}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_1997, Midori_rounds_sub_sBox_PRINCE_13_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .a ({new_AGEMA_signal_1768, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_1771, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_1998, Midori_rounds_sub_sBox_PRINCE_13_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .a ({new_AGEMA_signal_1768, Midori_rounds_roundReg_out[54]}), .b ({new_AGEMA_signal_1766, Midori_rounds_roundReg_out[55]}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_1769, Midori_rounds_sub_sBox_PRINCE_13_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .a ({new_AGEMA_signal_1772, Midori_rounds_sub_sBox_PRINCE_13_n9}), .b ({new_AGEMA_signal_1771, Midori_rounds_sub_sBox_PRINCE_13_n8}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_2000, Midori_rounds_sub_sBox_PRINCE_13_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .a ({new_AGEMA_signal_1773, Midori_rounds_roundReg_out[56]}), .b ({new_AGEMA_signal_1774, Midori_rounds_roundReg_out[59]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_1775, Midori_rounds_sub_sBox_PRINCE_14_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .a ({new_AGEMA_signal_1779, Midori_rounds_sub_sBox_PRINCE_14_n8}), .b ({new_AGEMA_signal_1778, Midori_rounds_sub_sBox_PRINCE_14_n7}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_2002, Midori_rounds_sub_sBox_PRINCE_14_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .a ({new_AGEMA_signal_1774, Midori_rounds_roundReg_out[59]}), .b ({new_AGEMA_signal_1780, Midori_rounds_sub_sBox_PRINCE_14_n9}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_2003, Midori_rounds_sub_sBox_PRINCE_14_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .a ({new_AGEMA_signal_1776, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_1779, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_2004, Midori_rounds_sub_sBox_PRINCE_14_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .a ({new_AGEMA_signal_1776, Midori_rounds_roundReg_out[58]}), .b ({new_AGEMA_signal_1774, Midori_rounds_roundReg_out[59]}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_1777, Midori_rounds_sub_sBox_PRINCE_14_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .a ({new_AGEMA_signal_1780, Midori_rounds_sub_sBox_PRINCE_14_n9}), .b ({new_AGEMA_signal_1779, Midori_rounds_sub_sBox_PRINCE_14_n8}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_14_n13}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .a ({new_AGEMA_signal_1781, Midori_rounds_roundReg_out[60]}), .b ({new_AGEMA_signal_1782, Midori_rounds_roundReg_out[63]}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_1783, Midori_rounds_sub_sBox_PRINCE_15_n10}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .a ({new_AGEMA_signal_1787, Midori_rounds_sub_sBox_PRINCE_15_n8}), .b ({new_AGEMA_signal_1786, Midori_rounds_sub_sBox_PRINCE_15_n7}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_2008, Midori_rounds_sub_sBox_PRINCE_15_n15}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .a ({new_AGEMA_signal_1782, Midori_rounds_roundReg_out[63]}), .b ({new_AGEMA_signal_1788, Midori_rounds_sub_sBox_PRINCE_15_n9}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_2009, Midori_rounds_sub_sBox_PRINCE_15_n4}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .a ({new_AGEMA_signal_1784, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_1787, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_2010, Midori_rounds_sub_sBox_PRINCE_15_n6}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U5 ( .a ({new_AGEMA_signal_1784, Midori_rounds_roundReg_out[62]}), .b ({new_AGEMA_signal_1782, Midori_rounds_roundReg_out[63]}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_1785, Midori_rounds_sub_sBox_PRINCE_15_n1}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U3 ( .a ({new_AGEMA_signal_1788, Midori_rounds_sub_sBox_PRINCE_15_n9}), .b ({new_AGEMA_signal_1787, Midori_rounds_sub_sBox_PRINCE_15_n8}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_2012, Midori_rounds_sub_sBox_PRINCE_15_n13}) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_3025), .Q (new_AGEMA_signal_3026) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (clk), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_3097) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (clk), .D (new_AGEMA_signal_3098), .Q (new_AGEMA_signal_3099) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (clk), .D (new_AGEMA_signal_3100), .Q (new_AGEMA_signal_3101) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (clk), .D (new_AGEMA_signal_3102), .Q (new_AGEMA_signal_3103) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (clk), .D (new_AGEMA_signal_3104), .Q (new_AGEMA_signal_3105) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (clk), .D (new_AGEMA_signal_3106), .Q (new_AGEMA_signal_3107) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_3109) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (clk), .D (new_AGEMA_signal_3110), .Q (new_AGEMA_signal_3111) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (clk), .D (new_AGEMA_signal_3112), .Q (new_AGEMA_signal_3113) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (clk), .D (new_AGEMA_signal_3114), .Q (new_AGEMA_signal_3115) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (clk), .D (new_AGEMA_signal_3116), .Q (new_AGEMA_signal_3117) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (clk), .D (new_AGEMA_signal_3118), .Q (new_AGEMA_signal_3119) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (clk), .D (new_AGEMA_signal_3120), .Q (new_AGEMA_signal_3121) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (clk), .D (new_AGEMA_signal_3122), .Q (new_AGEMA_signal_3123) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (clk), .D (new_AGEMA_signal_3124), .Q (new_AGEMA_signal_3125) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (clk), .D (new_AGEMA_signal_3126), .Q (new_AGEMA_signal_3127) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (clk), .D (new_AGEMA_signal_3128), .Q (new_AGEMA_signal_3129) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (clk), .D (new_AGEMA_signal_3130), .Q (new_AGEMA_signal_3131) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (clk), .D (new_AGEMA_signal_3132), .Q (new_AGEMA_signal_3133) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (clk), .D (new_AGEMA_signal_3134), .Q (new_AGEMA_signal_3135) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (clk), .D (new_AGEMA_signal_3136), .Q (new_AGEMA_signal_3137) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (clk), .D (new_AGEMA_signal_3138), .Q (new_AGEMA_signal_3139) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (clk), .D (new_AGEMA_signal_3140), .Q (new_AGEMA_signal_3141) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (clk), .D (new_AGEMA_signal_3142), .Q (new_AGEMA_signal_3143) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (clk), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_3145) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (clk), .D (new_AGEMA_signal_3146), .Q (new_AGEMA_signal_3147) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (clk), .D (new_AGEMA_signal_3148), .Q (new_AGEMA_signal_3149) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (clk), .D (new_AGEMA_signal_3150), .Q (new_AGEMA_signal_3151) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (clk), .D (new_AGEMA_signal_3152), .Q (new_AGEMA_signal_3153) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (clk), .D (new_AGEMA_signal_3154), .Q (new_AGEMA_signal_3155) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (clk), .D (new_AGEMA_signal_3156), .Q (new_AGEMA_signal_3157) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (clk), .D (new_AGEMA_signal_3158), .Q (new_AGEMA_signal_3159) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (clk), .D (new_AGEMA_signal_3160), .Q (new_AGEMA_signal_3161) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (clk), .D (new_AGEMA_signal_3162), .Q (new_AGEMA_signal_3163) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (clk), .D (new_AGEMA_signal_3164), .Q (new_AGEMA_signal_3165) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (clk), .D (new_AGEMA_signal_3166), .Q (new_AGEMA_signal_3167) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (clk), .D (new_AGEMA_signal_3168), .Q (new_AGEMA_signal_3169) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (clk), .D (new_AGEMA_signal_3170), .Q (new_AGEMA_signal_3171) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (clk), .D (new_AGEMA_signal_3172), .Q (new_AGEMA_signal_3173) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (clk), .D (new_AGEMA_signal_3174), .Q (new_AGEMA_signal_3175) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (clk), .D (new_AGEMA_signal_3176), .Q (new_AGEMA_signal_3177) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (clk), .D (new_AGEMA_signal_3178), .Q (new_AGEMA_signal_3179) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (clk), .D (new_AGEMA_signal_3180), .Q (new_AGEMA_signal_3181) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (clk), .D (new_AGEMA_signal_3182), .Q (new_AGEMA_signal_3183) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (clk), .D (new_AGEMA_signal_3184), .Q (new_AGEMA_signal_3185) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (clk), .D (new_AGEMA_signal_3186), .Q (new_AGEMA_signal_3187) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (clk), .D (new_AGEMA_signal_3188), .Q (new_AGEMA_signal_3189) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (clk), .D (new_AGEMA_signal_3190), .Q (new_AGEMA_signal_3191) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (clk), .D (new_AGEMA_signal_3192), .Q (new_AGEMA_signal_3193) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (clk), .D (new_AGEMA_signal_3194), .Q (new_AGEMA_signal_3195) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (clk), .D (new_AGEMA_signal_3196), .Q (new_AGEMA_signal_3197) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (clk), .D (new_AGEMA_signal_3198), .Q (new_AGEMA_signal_3199) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (clk), .D (new_AGEMA_signal_3200), .Q (new_AGEMA_signal_3201) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (clk), .D (new_AGEMA_signal_3202), .Q (new_AGEMA_signal_3203) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (clk), .D (new_AGEMA_signal_3204), .Q (new_AGEMA_signal_3205) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (clk), .D (new_AGEMA_signal_3206), .Q (new_AGEMA_signal_3207) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (clk), .D (new_AGEMA_signal_3208), .Q (new_AGEMA_signal_3209) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (clk), .D (new_AGEMA_signal_3210), .Q (new_AGEMA_signal_3211) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (clk), .D (new_AGEMA_signal_3212), .Q (new_AGEMA_signal_3213) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (clk), .D (new_AGEMA_signal_3214), .Q (new_AGEMA_signal_3215) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (clk), .D (new_AGEMA_signal_3216), .Q (new_AGEMA_signal_3217) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (clk), .D (new_AGEMA_signal_3218), .Q (new_AGEMA_signal_3219) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (clk), .D (new_AGEMA_signal_3220), .Q (new_AGEMA_signal_3221) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (clk), .D (new_AGEMA_signal_3222), .Q (new_AGEMA_signal_3223) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (clk), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_3225) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (clk), .D (new_AGEMA_signal_3226), .Q (new_AGEMA_signal_3227) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (clk), .D (new_AGEMA_signal_3228), .Q (new_AGEMA_signal_3229) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (clk), .D (new_AGEMA_signal_3230), .Q (new_AGEMA_signal_3231) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (clk), .D (new_AGEMA_signal_3232), .Q (new_AGEMA_signal_3233) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (clk), .D (new_AGEMA_signal_3234), .Q (new_AGEMA_signal_3235) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (clk), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_3237) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (clk), .D (new_AGEMA_signal_3238), .Q (new_AGEMA_signal_3239) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (clk), .D (new_AGEMA_signal_3240), .Q (new_AGEMA_signal_3241) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (clk), .D (new_AGEMA_signal_3242), .Q (new_AGEMA_signal_3243) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (clk), .D (new_AGEMA_signal_3244), .Q (new_AGEMA_signal_3245) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (clk), .D (new_AGEMA_signal_3246), .Q (new_AGEMA_signal_3247) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (clk), .D (new_AGEMA_signal_3248), .Q (new_AGEMA_signal_3249) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (clk), .D (new_AGEMA_signal_3250), .Q (new_AGEMA_signal_3251) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (clk), .D (new_AGEMA_signal_3252), .Q (new_AGEMA_signal_3253) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (clk), .D (new_AGEMA_signal_3254), .Q (new_AGEMA_signal_3255) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (clk), .D (new_AGEMA_signal_3256), .Q (new_AGEMA_signal_3257) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (clk), .D (new_AGEMA_signal_3258), .Q (new_AGEMA_signal_3259) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (clk), .D (new_AGEMA_signal_3260), .Q (new_AGEMA_signal_3261) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (clk), .D (new_AGEMA_signal_3262), .Q (new_AGEMA_signal_3263) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (clk), .D (new_AGEMA_signal_3264), .Q (new_AGEMA_signal_3265) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (clk), .D (new_AGEMA_signal_3266), .Q (new_AGEMA_signal_3267) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (clk), .D (new_AGEMA_signal_3268), .Q (new_AGEMA_signal_3269) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (clk), .D (new_AGEMA_signal_3270), .Q (new_AGEMA_signal_3271) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (clk), .D (new_AGEMA_signal_3272), .Q (new_AGEMA_signal_3273) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (clk), .D (new_AGEMA_signal_3274), .Q (new_AGEMA_signal_3275) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (clk), .D (new_AGEMA_signal_3276), .Q (new_AGEMA_signal_3277) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (clk), .D (new_AGEMA_signal_3278), .Q (new_AGEMA_signal_3279) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (clk), .D (new_AGEMA_signal_3280), .Q (new_AGEMA_signal_3281) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (clk), .D (new_AGEMA_signal_3282), .Q (new_AGEMA_signal_3283) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (clk), .D (new_AGEMA_signal_3284), .Q (new_AGEMA_signal_3285) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (clk), .D (new_AGEMA_signal_3286), .Q (new_AGEMA_signal_3287) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (clk), .D (new_AGEMA_signal_3288), .Q (new_AGEMA_signal_3289) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (clk), .D (new_AGEMA_signal_3290), .Q (new_AGEMA_signal_3291) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (clk), .D (new_AGEMA_signal_3292), .Q (new_AGEMA_signal_3293) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (clk), .D (new_AGEMA_signal_3294), .Q (new_AGEMA_signal_3295) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (clk), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_3297) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (clk), .D (new_AGEMA_signal_3298), .Q (new_AGEMA_signal_3299) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (clk), .D (new_AGEMA_signal_3300), .Q (new_AGEMA_signal_3301) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (clk), .D (new_AGEMA_signal_3302), .Q (new_AGEMA_signal_3303) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (clk), .D (new_AGEMA_signal_3304), .Q (new_AGEMA_signal_3305) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (clk), .D (new_AGEMA_signal_3306), .Q (new_AGEMA_signal_3307) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (clk), .D (new_AGEMA_signal_3308), .Q (new_AGEMA_signal_3309) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (clk), .D (new_AGEMA_signal_3310), .Q (new_AGEMA_signal_3311) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (clk), .D (new_AGEMA_signal_3312), .Q (new_AGEMA_signal_3313) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (clk), .D (new_AGEMA_signal_3314), .Q (new_AGEMA_signal_3315) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (clk), .D (new_AGEMA_signal_3316), .Q (new_AGEMA_signal_3317) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (clk), .D (new_AGEMA_signal_3318), .Q (new_AGEMA_signal_3319) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (clk), .D (new_AGEMA_signal_3320), .Q (new_AGEMA_signal_3321) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (clk), .D (new_AGEMA_signal_3322), .Q (new_AGEMA_signal_3323) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (clk), .D (new_AGEMA_signal_3324), .Q (new_AGEMA_signal_3325) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (clk), .D (new_AGEMA_signal_3326), .Q (new_AGEMA_signal_3327) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (clk), .D (new_AGEMA_signal_3328), .Q (new_AGEMA_signal_3329) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (clk), .D (new_AGEMA_signal_3330), .Q (new_AGEMA_signal_3331) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (clk), .D (new_AGEMA_signal_3332), .Q (new_AGEMA_signal_3333) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (clk), .D (new_AGEMA_signal_3334), .Q (new_AGEMA_signal_3335) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (clk), .D (new_AGEMA_signal_3336), .Q (new_AGEMA_signal_3337) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (clk), .D (new_AGEMA_signal_3338), .Q (new_AGEMA_signal_3339) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (clk), .D (new_AGEMA_signal_3340), .Q (new_AGEMA_signal_3341) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (clk), .D (new_AGEMA_signal_3342), .Q (new_AGEMA_signal_3343) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (clk), .D (new_AGEMA_signal_3344), .Q (new_AGEMA_signal_3345) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (clk), .D (new_AGEMA_signal_3346), .Q (new_AGEMA_signal_3347) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (clk), .D (new_AGEMA_signal_3348), .Q (new_AGEMA_signal_3349) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (clk), .D (new_AGEMA_signal_3350), .Q (new_AGEMA_signal_3351) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (clk), .D (new_AGEMA_signal_3352), .Q (new_AGEMA_signal_3353) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (clk), .D (new_AGEMA_signal_3358), .Q (new_AGEMA_signal_3359) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (clk), .D (new_AGEMA_signal_3364), .Q (new_AGEMA_signal_3365) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (clk), .D (new_AGEMA_signal_3370), .Q (new_AGEMA_signal_3371) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (clk), .D (new_AGEMA_signal_3376), .Q (new_AGEMA_signal_3377) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (clk), .D (new_AGEMA_signal_3382), .Q (new_AGEMA_signal_3383) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (clk), .D (new_AGEMA_signal_3388), .Q (new_AGEMA_signal_3389) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (clk), .D (new_AGEMA_signal_3394), .Q (new_AGEMA_signal_3395) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (clk), .D (new_AGEMA_signal_3400), .Q (new_AGEMA_signal_3401) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (clk), .D (new_AGEMA_signal_3406), .Q (new_AGEMA_signal_3407) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (clk), .D (new_AGEMA_signal_3412), .Q (new_AGEMA_signal_3413) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (clk), .D (new_AGEMA_signal_3418), .Q (new_AGEMA_signal_3419) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (clk), .D (new_AGEMA_signal_3424), .Q (new_AGEMA_signal_3425) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (clk), .D (new_AGEMA_signal_3430), .Q (new_AGEMA_signal_3431) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (clk), .D (new_AGEMA_signal_3436), .Q (new_AGEMA_signal_3437) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (clk), .D (new_AGEMA_signal_3442), .Q (new_AGEMA_signal_3443) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (clk), .D (new_AGEMA_signal_3448), .Q (new_AGEMA_signal_3449) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (clk), .D (new_AGEMA_signal_3454), .Q (new_AGEMA_signal_3455) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (clk), .D (new_AGEMA_signal_3460), .Q (new_AGEMA_signal_3461) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (clk), .D (new_AGEMA_signal_3466), .Q (new_AGEMA_signal_3467) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (clk), .D (new_AGEMA_signal_3472), .Q (new_AGEMA_signal_3473) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (clk), .D (new_AGEMA_signal_3478), .Q (new_AGEMA_signal_3479) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (clk), .D (new_AGEMA_signal_3484), .Q (new_AGEMA_signal_3485) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (clk), .D (new_AGEMA_signal_3490), .Q (new_AGEMA_signal_3491) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (clk), .D (new_AGEMA_signal_3496), .Q (new_AGEMA_signal_3497) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (clk), .D (new_AGEMA_signal_3502), .Q (new_AGEMA_signal_3503) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (clk), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_3509) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (clk), .D (new_AGEMA_signal_3514), .Q (new_AGEMA_signal_3515) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (clk), .D (new_AGEMA_signal_3520), .Q (new_AGEMA_signal_3521) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (clk), .D (new_AGEMA_signal_3526), .Q (new_AGEMA_signal_3527) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (clk), .D (new_AGEMA_signal_3532), .Q (new_AGEMA_signal_3533) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (clk), .D (new_AGEMA_signal_3538), .Q (new_AGEMA_signal_3539) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (clk), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_3545) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (clk), .D (new_AGEMA_signal_3550), .Q (new_AGEMA_signal_3551) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (clk), .D (new_AGEMA_signal_3556), .Q (new_AGEMA_signal_3557) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (clk), .D (new_AGEMA_signal_3562), .Q (new_AGEMA_signal_3563) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (clk), .D (new_AGEMA_signal_3568), .Q (new_AGEMA_signal_3569) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (clk), .D (new_AGEMA_signal_3574), .Q (new_AGEMA_signal_3575) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (clk), .D (new_AGEMA_signal_3580), .Q (new_AGEMA_signal_3581) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (clk), .D (new_AGEMA_signal_3586), .Q (new_AGEMA_signal_3587) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (clk), .D (new_AGEMA_signal_3592), .Q (new_AGEMA_signal_3593) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (clk), .D (new_AGEMA_signal_3598), .Q (new_AGEMA_signal_3599) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (clk), .D (new_AGEMA_signal_3604), .Q (new_AGEMA_signal_3605) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (clk), .D (new_AGEMA_signal_3610), .Q (new_AGEMA_signal_3611) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (clk), .D (new_AGEMA_signal_3616), .Q (new_AGEMA_signal_3617) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (clk), .D (new_AGEMA_signal_3622), .Q (new_AGEMA_signal_3623) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (clk), .D (new_AGEMA_signal_3628), .Q (new_AGEMA_signal_3629) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (clk), .D (new_AGEMA_signal_3634), .Q (new_AGEMA_signal_3635) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (clk), .D (new_AGEMA_signal_3640), .Q (new_AGEMA_signal_3641) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (clk), .D (new_AGEMA_signal_3646), .Q (new_AGEMA_signal_3647) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (clk), .D (new_AGEMA_signal_3652), .Q (new_AGEMA_signal_3653) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (clk), .D (new_AGEMA_signal_3658), .Q (new_AGEMA_signal_3659) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (clk), .D (new_AGEMA_signal_3664), .Q (new_AGEMA_signal_3665) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (clk), .D (new_AGEMA_signal_3670), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (clk), .D (new_AGEMA_signal_3676), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (clk), .D (new_AGEMA_signal_3682), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (clk), .D (new_AGEMA_signal_3688), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (clk), .D (new_AGEMA_signal_3694), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (clk), .D (new_AGEMA_signal_3700), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (clk), .D (new_AGEMA_signal_3706), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (clk), .D (new_AGEMA_signal_3712), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (clk), .D (new_AGEMA_signal_3718), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (clk), .D (new_AGEMA_signal_3724), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (clk), .D (new_AGEMA_signal_3730), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (clk), .D (new_AGEMA_signal_3736), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (clk), .D (new_AGEMA_signal_3742), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (clk), .D (new_AGEMA_signal_3748), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (clk), .D (new_AGEMA_signal_3754), .Q (new_AGEMA_signal_3755) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (clk), .D (new_AGEMA_signal_3760), .Q (new_AGEMA_signal_3761) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_3766), .Q (new_AGEMA_signal_3767) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_3772), .Q (new_AGEMA_signal_3773) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_3778), .Q (new_AGEMA_signal_3779) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_3784), .Q (new_AGEMA_signal_3785) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_3790), .Q (new_AGEMA_signal_3791) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_3796), .Q (new_AGEMA_signal_3797) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_3802), .Q (new_AGEMA_signal_3803) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_3808), .Q (new_AGEMA_signal_3809) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_3814), .Q (new_AGEMA_signal_3815) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_3820), .Q (new_AGEMA_signal_3821) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_3826), .Q (new_AGEMA_signal_3827) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_3832), .Q (new_AGEMA_signal_3833) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_3839) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_3844), .Q (new_AGEMA_signal_3845) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_3850), .Q (new_AGEMA_signal_3851) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_3856), .Q (new_AGEMA_signal_3857) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_3863) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_3868), .Q (new_AGEMA_signal_3869) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_3874), .Q (new_AGEMA_signal_3875) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_3880), .Q (new_AGEMA_signal_3881) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_3887) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_3892), .Q (new_AGEMA_signal_3893) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_3898), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_3904), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_3922), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_3940), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_3964), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_3970), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_4006), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_4018), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_4024), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_4036), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_4042), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_4054), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_4060), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_4066), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_4072), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_4078), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_4084), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_4090), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_4096), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_4102), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_4108), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_4114), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_4120), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_4132), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_4138), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_4144), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_4156), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_4162), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_4168), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_4174), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_4186), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_4192), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_4204), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_4210), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_4216), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_4222), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_4234), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_4240), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_4246), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_4252), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_4258), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_4264), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_4270), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_4276), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_4282), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_4288), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_4306), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_4330), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_4354), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_4372), .Q (new_AGEMA_signal_4373) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_4378), .Q (new_AGEMA_signal_4379) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_4384), .Q (new_AGEMA_signal_4385) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_4390), .Q (new_AGEMA_signal_4391) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_4396), .Q (new_AGEMA_signal_4397) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_4402), .Q (new_AGEMA_signal_4403) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_4408), .Q (new_AGEMA_signal_4409) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_4414), .Q (new_AGEMA_signal_4415) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_4420), .Q (new_AGEMA_signal_4421) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_4426), .Q (new_AGEMA_signal_4427) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_4432), .Q (new_AGEMA_signal_4433) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_4438), .Q (new_AGEMA_signal_4439) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_4444), .Q (new_AGEMA_signal_4445) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_4450), .Q (new_AGEMA_signal_4451) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_4456), .Q (new_AGEMA_signal_4457) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_4462), .Q (new_AGEMA_signal_4463) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_4468), .Q (new_AGEMA_signal_4469) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_4474), .Q (new_AGEMA_signal_4475) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_4480), .Q (new_AGEMA_signal_4481) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_4486), .Q (new_AGEMA_signal_4487) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_4492), .Q (new_AGEMA_signal_4493) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_4498), .Q (new_AGEMA_signal_4499) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_4504), .Q (new_AGEMA_signal_4505) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_4703) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_4709) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_4717) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_4740), .Q (new_AGEMA_signal_4741) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_4836), .Q (new_AGEMA_signal_4837) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_4861) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_4884), .Q (new_AGEMA_signal_4885) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_4893) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_4901) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_4908), .Q (new_AGEMA_signal_4909) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_4917) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_4925) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_4932), .Q (new_AGEMA_signal_4933) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_4940), .Q (new_AGEMA_signal_4941) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_4949) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_4956), .Q (new_AGEMA_signal_4957) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_4964), .Q (new_AGEMA_signal_4965) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_4973) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_4980), .Q (new_AGEMA_signal_4981) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_4988), .Q (new_AGEMA_signal_4989) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_4997) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_5005) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_5012), .Q (new_AGEMA_signal_5013) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_5021) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_5028), .Q (new_AGEMA_signal_5029) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_5036), .Q (new_AGEMA_signal_5037) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_5045) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_5052), .Q (new_AGEMA_signal_5053) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_5060), .Q (new_AGEMA_signal_5061) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_5069) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_5077) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_5084), .Q (new_AGEMA_signal_5085) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_5093) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_5100), .Q (new_AGEMA_signal_5101) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_5108), .Q (new_AGEMA_signal_5109) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_5117) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_5124), .Q (new_AGEMA_signal_5125) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_5132), .Q (new_AGEMA_signal_5133) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_5141) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_5149) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_5156), .Q (new_AGEMA_signal_5157) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_5165) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_5172), .Q (new_AGEMA_signal_5173) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_5180), .Q (new_AGEMA_signal_5181) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_5189) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_5197) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_5204), .Q (new_AGEMA_signal_5205) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_5213) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_5221) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_5228), .Q (new_AGEMA_signal_5229) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_5237) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_5244), .Q (new_AGEMA_signal_5245) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_5252), .Q (new_AGEMA_signal_5253) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_5261) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_5269) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_5276), .Q (new_AGEMA_signal_5277) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_5285) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_5293) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_5300), .Q (new_AGEMA_signal_5301) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_5309) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_5316), .Q (new_AGEMA_signal_5317) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_5324), .Q (new_AGEMA_signal_5325) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_5332), .Q (new_AGEMA_signal_5333) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_5341) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_5348), .Q (new_AGEMA_signal_5349) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_5357) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_5365) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_5389) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_5396), .Q (new_AGEMA_signal_5397) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_5413) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_5421) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_5735) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_5743) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_5751) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_5759) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_5767) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_5775) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_5783) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_5807) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_5831) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_5855) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_5879) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_5903) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_5927) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_5951) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_5975) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_5999) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_6023) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_6047) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_6071) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_6095) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_6119) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_6143) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_6166), .Q (new_AGEMA_signal_6167) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_6191) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_6215) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_6238), .Q (new_AGEMA_signal_6239) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_6441) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_6449) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_6465) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_3026), .Q (new_AGEMA_signal_3027) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (clk), .D (new_AGEMA_signal_3353), .Q (new_AGEMA_signal_3354) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (clk), .D (new_AGEMA_signal_3359), .Q (new_AGEMA_signal_3360) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (clk), .D (new_AGEMA_signal_3365), .Q (new_AGEMA_signal_3366) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (clk), .D (new_AGEMA_signal_3371), .Q (new_AGEMA_signal_3372) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (clk), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_3378) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (clk), .D (new_AGEMA_signal_3383), .Q (new_AGEMA_signal_3384) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (clk), .D (new_AGEMA_signal_3389), .Q (new_AGEMA_signal_3390) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (clk), .D (new_AGEMA_signal_3395), .Q (new_AGEMA_signal_3396) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (clk), .D (new_AGEMA_signal_3401), .Q (new_AGEMA_signal_3402) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (clk), .D (new_AGEMA_signal_3407), .Q (new_AGEMA_signal_3408) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (clk), .D (new_AGEMA_signal_3413), .Q (new_AGEMA_signal_3414) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (clk), .D (new_AGEMA_signal_3419), .Q (new_AGEMA_signal_3420) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (clk), .D (new_AGEMA_signal_3425), .Q (new_AGEMA_signal_3426) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (clk), .D (new_AGEMA_signal_3431), .Q (new_AGEMA_signal_3432) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (clk), .D (new_AGEMA_signal_3437), .Q (new_AGEMA_signal_3438) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (clk), .D (new_AGEMA_signal_3443), .Q (new_AGEMA_signal_3444) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (clk), .D (new_AGEMA_signal_3449), .Q (new_AGEMA_signal_3450) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (clk), .D (new_AGEMA_signal_3455), .Q (new_AGEMA_signal_3456) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (clk), .D (new_AGEMA_signal_3461), .Q (new_AGEMA_signal_3462) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (clk), .D (new_AGEMA_signal_3467), .Q (new_AGEMA_signal_3468) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (clk), .D (new_AGEMA_signal_3473), .Q (new_AGEMA_signal_3474) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (clk), .D (new_AGEMA_signal_3479), .Q (new_AGEMA_signal_3480) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (clk), .D (new_AGEMA_signal_3485), .Q (new_AGEMA_signal_3486) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (clk), .D (new_AGEMA_signal_3491), .Q (new_AGEMA_signal_3492) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (clk), .D (new_AGEMA_signal_3497), .Q (new_AGEMA_signal_3498) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (clk), .D (new_AGEMA_signal_3503), .Q (new_AGEMA_signal_3504) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (clk), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_3510) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (clk), .D (new_AGEMA_signal_3515), .Q (new_AGEMA_signal_3516) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (clk), .D (new_AGEMA_signal_3521), .Q (new_AGEMA_signal_3522) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (clk), .D (new_AGEMA_signal_3527), .Q (new_AGEMA_signal_3528) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (clk), .D (new_AGEMA_signal_3533), .Q (new_AGEMA_signal_3534) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (clk), .D (new_AGEMA_signal_3539), .Q (new_AGEMA_signal_3540) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (clk), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_3546) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (clk), .D (new_AGEMA_signal_3551), .Q (new_AGEMA_signal_3552) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (clk), .D (new_AGEMA_signal_3557), .Q (new_AGEMA_signal_3558) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (clk), .D (new_AGEMA_signal_3563), .Q (new_AGEMA_signal_3564) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (clk), .D (new_AGEMA_signal_3569), .Q (new_AGEMA_signal_3570) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (clk), .D (new_AGEMA_signal_3575), .Q (new_AGEMA_signal_3576) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (clk), .D (new_AGEMA_signal_3581), .Q (new_AGEMA_signal_3582) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (clk), .D (new_AGEMA_signal_3587), .Q (new_AGEMA_signal_3588) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (clk), .D (new_AGEMA_signal_3593), .Q (new_AGEMA_signal_3594) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (clk), .D (new_AGEMA_signal_3599), .Q (new_AGEMA_signal_3600) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (clk), .D (new_AGEMA_signal_3605), .Q (new_AGEMA_signal_3606) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (clk), .D (new_AGEMA_signal_3611), .Q (new_AGEMA_signal_3612) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (clk), .D (new_AGEMA_signal_3617), .Q (new_AGEMA_signal_3618) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (clk), .D (new_AGEMA_signal_3623), .Q (new_AGEMA_signal_3624) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (clk), .D (new_AGEMA_signal_3629), .Q (new_AGEMA_signal_3630) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (clk), .D (new_AGEMA_signal_3635), .Q (new_AGEMA_signal_3636) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (clk), .D (new_AGEMA_signal_3641), .Q (new_AGEMA_signal_3642) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (clk), .D (new_AGEMA_signal_3647), .Q (new_AGEMA_signal_3648) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (clk), .D (new_AGEMA_signal_3653), .Q (new_AGEMA_signal_3654) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (clk), .D (new_AGEMA_signal_3659), .Q (new_AGEMA_signal_3660) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (clk), .D (new_AGEMA_signal_3665), .Q (new_AGEMA_signal_3666) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (clk), .D (new_AGEMA_signal_3671), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (clk), .D (new_AGEMA_signal_3677), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (clk), .D (new_AGEMA_signal_3683), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (clk), .D (new_AGEMA_signal_3689), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (clk), .D (new_AGEMA_signal_3695), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (clk), .D (new_AGEMA_signal_3701), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (clk), .D (new_AGEMA_signal_3707), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (clk), .D (new_AGEMA_signal_3713), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (clk), .D (new_AGEMA_signal_3719), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (clk), .D (new_AGEMA_signal_3725), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (clk), .D (new_AGEMA_signal_3731), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (clk), .D (new_AGEMA_signal_3737), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (clk), .D (new_AGEMA_signal_3743), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (clk), .D (new_AGEMA_signal_3749), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (clk), .D (new_AGEMA_signal_3755), .Q (new_AGEMA_signal_3756) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (clk), .D (new_AGEMA_signal_3761), .Q (new_AGEMA_signal_3762) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (clk), .D (new_AGEMA_signal_3767), .Q (new_AGEMA_signal_3768) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (clk), .D (new_AGEMA_signal_3773), .Q (new_AGEMA_signal_3774) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (clk), .D (new_AGEMA_signal_3779), .Q (new_AGEMA_signal_3780) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (clk), .D (new_AGEMA_signal_3785), .Q (new_AGEMA_signal_3786) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (clk), .D (new_AGEMA_signal_3791), .Q (new_AGEMA_signal_3792) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (clk), .D (new_AGEMA_signal_3797), .Q (new_AGEMA_signal_3798) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (clk), .D (new_AGEMA_signal_3803), .Q (new_AGEMA_signal_3804) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (clk), .D (new_AGEMA_signal_3809), .Q (new_AGEMA_signal_3810) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (clk), .D (new_AGEMA_signal_3815), .Q (new_AGEMA_signal_3816) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (clk), .D (new_AGEMA_signal_3821), .Q (new_AGEMA_signal_3822) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (clk), .D (new_AGEMA_signal_3827), .Q (new_AGEMA_signal_3828) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_3833), .Q (new_AGEMA_signal_3834) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (clk), .D (new_AGEMA_signal_3839), .Q (new_AGEMA_signal_3840) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_3845), .Q (new_AGEMA_signal_3846) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (clk), .D (new_AGEMA_signal_3851), .Q (new_AGEMA_signal_3852) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_3857), .Q (new_AGEMA_signal_3858) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_3863), .Q (new_AGEMA_signal_3864) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (clk), .D (new_AGEMA_signal_3869), .Q (new_AGEMA_signal_3870) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_3875), .Q (new_AGEMA_signal_3876) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (clk), .D (new_AGEMA_signal_3881), .Q (new_AGEMA_signal_3882) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_3887), .Q (new_AGEMA_signal_3888) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (clk), .D (new_AGEMA_signal_3893), .Q (new_AGEMA_signal_3894) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_3899), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (clk), .D (new_AGEMA_signal_3905), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_3911), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (clk), .D (new_AGEMA_signal_3917), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_3923), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (clk), .D (new_AGEMA_signal_3929), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_3935), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (clk), .D (new_AGEMA_signal_3941), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_3947), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (clk), .D (new_AGEMA_signal_3953), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_3959), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (clk), .D (new_AGEMA_signal_3965), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_3971), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (clk), .D (new_AGEMA_signal_3977), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_3983), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (clk), .D (new_AGEMA_signal_3989), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_3995), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (clk), .D (new_AGEMA_signal_4001), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_4007), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (clk), .D (new_AGEMA_signal_4013), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_4019), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (clk), .D (new_AGEMA_signal_4025), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_4031), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (clk), .D (new_AGEMA_signal_4037), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_4043), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (clk), .D (new_AGEMA_signal_4049), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_4055), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (clk), .D (new_AGEMA_signal_4061), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_4067), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (clk), .D (new_AGEMA_signal_4073), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_4079), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (clk), .D (new_AGEMA_signal_4085), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_4091), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (clk), .D (new_AGEMA_signal_4097), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_4103), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (clk), .D (new_AGEMA_signal_4109), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_4115), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (clk), .D (new_AGEMA_signal_4121), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (clk), .D (new_AGEMA_signal_4127), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (clk), .D (new_AGEMA_signal_4133), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (clk), .D (new_AGEMA_signal_4139), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (clk), .D (new_AGEMA_signal_4145), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (clk), .D (new_AGEMA_signal_4151), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (clk), .D (new_AGEMA_signal_4157), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (clk), .D (new_AGEMA_signal_4163), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (clk), .D (new_AGEMA_signal_4169), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (clk), .D (new_AGEMA_signal_4175), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (clk), .D (new_AGEMA_signal_4181), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (clk), .D (new_AGEMA_signal_4187), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (clk), .D (new_AGEMA_signal_4193), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (clk), .D (new_AGEMA_signal_4199), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (clk), .D (new_AGEMA_signal_4205), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (clk), .D (new_AGEMA_signal_4211), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (clk), .D (new_AGEMA_signal_4217), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (clk), .D (new_AGEMA_signal_4223), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (clk), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (clk), .D (new_AGEMA_signal_4235), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (clk), .D (new_AGEMA_signal_4241), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (clk), .D (new_AGEMA_signal_4247), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (clk), .D (new_AGEMA_signal_4253), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (clk), .D (new_AGEMA_signal_4259), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (clk), .D (new_AGEMA_signal_4265), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (clk), .D (new_AGEMA_signal_4271), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (clk), .D (new_AGEMA_signal_4277), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (clk), .D (new_AGEMA_signal_4283), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (clk), .D (new_AGEMA_signal_4289), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (clk), .D (new_AGEMA_signal_4295), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (clk), .D (new_AGEMA_signal_4301), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (clk), .D (new_AGEMA_signal_4307), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (clk), .D (new_AGEMA_signal_4313), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (clk), .D (new_AGEMA_signal_4319), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (clk), .D (new_AGEMA_signal_4325), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (clk), .D (new_AGEMA_signal_4331), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (clk), .D (new_AGEMA_signal_4337), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (clk), .D (new_AGEMA_signal_4343), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (clk), .D (new_AGEMA_signal_4349), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (clk), .D (new_AGEMA_signal_4355), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (clk), .D (new_AGEMA_signal_4361), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (clk), .D (new_AGEMA_signal_4367), .Q (new_AGEMA_signal_4368) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (clk), .D (new_AGEMA_signal_4373), .Q (new_AGEMA_signal_4374) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (clk), .D (new_AGEMA_signal_4379), .Q (new_AGEMA_signal_4380) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (clk), .D (new_AGEMA_signal_4385), .Q (new_AGEMA_signal_4386) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (clk), .D (new_AGEMA_signal_4391), .Q (new_AGEMA_signal_4392) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (clk), .D (new_AGEMA_signal_4397), .Q (new_AGEMA_signal_4398) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (clk), .D (new_AGEMA_signal_4403), .Q (new_AGEMA_signal_4404) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (clk), .D (new_AGEMA_signal_4409), .Q (new_AGEMA_signal_4410) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (clk), .D (new_AGEMA_signal_4415), .Q (new_AGEMA_signal_4416) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (clk), .D (new_AGEMA_signal_4421), .Q (new_AGEMA_signal_4422) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (clk), .D (new_AGEMA_signal_4427), .Q (new_AGEMA_signal_4428) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (clk), .D (new_AGEMA_signal_4433), .Q (new_AGEMA_signal_4434) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (clk), .D (new_AGEMA_signal_4439), .Q (new_AGEMA_signal_4440) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (clk), .D (new_AGEMA_signal_4445), .Q (new_AGEMA_signal_4446) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (clk), .D (new_AGEMA_signal_4451), .Q (new_AGEMA_signal_4452) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (clk), .D (new_AGEMA_signal_4457), .Q (new_AGEMA_signal_4458) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (clk), .D (new_AGEMA_signal_4463), .Q (new_AGEMA_signal_4464) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (clk), .D (new_AGEMA_signal_4469), .Q (new_AGEMA_signal_4470) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (clk), .D (new_AGEMA_signal_4475), .Q (new_AGEMA_signal_4476) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (clk), .D (new_AGEMA_signal_4481), .Q (new_AGEMA_signal_4482) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (clk), .D (new_AGEMA_signal_4487), .Q (new_AGEMA_signal_4488) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (clk), .D (new_AGEMA_signal_4493), .Q (new_AGEMA_signal_4494) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (clk), .D (new_AGEMA_signal_4499), .Q (new_AGEMA_signal_4500) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (clk), .D (new_AGEMA_signal_4505), .Q (new_AGEMA_signal_4506) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n15), .Q (new_AGEMA_signal_4510) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (clk), .D (new_AGEMA_signal_1918), .Q (new_AGEMA_signal_4512) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_4514) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_3099), .Q (new_AGEMA_signal_4516) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n6), .Q (new_AGEMA_signal_4518) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_1920), .Q (new_AGEMA_signal_4520) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n15), .Q (new_AGEMA_signal_4522) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (clk), .D (new_AGEMA_signal_1924), .Q (new_AGEMA_signal_4524) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_3113), .Q (new_AGEMA_signal_4526) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_3115), .Q (new_AGEMA_signal_4528) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n6), .Q (new_AGEMA_signal_4530) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_1926), .Q (new_AGEMA_signal_4532) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n15), .Q (new_AGEMA_signal_4534) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (clk), .D (new_AGEMA_signal_1930), .Q (new_AGEMA_signal_4536) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_3129), .Q (new_AGEMA_signal_4538) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_3131), .Q (new_AGEMA_signal_4540) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n6), .Q (new_AGEMA_signal_4542) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_1932), .Q (new_AGEMA_signal_4544) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n15), .Q (new_AGEMA_signal_4546) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (clk), .D (new_AGEMA_signal_1936), .Q (new_AGEMA_signal_4548) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_3145), .Q (new_AGEMA_signal_4550) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_3147), .Q (new_AGEMA_signal_4552) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n6), .Q (new_AGEMA_signal_4554) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_1938), .Q (new_AGEMA_signal_4556) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n15), .Q (new_AGEMA_signal_4558) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_1942), .Q (new_AGEMA_signal_4560) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (new_AGEMA_signal_3161), .Q (new_AGEMA_signal_4562) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_3163), .Q (new_AGEMA_signal_4564) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n6), .Q (new_AGEMA_signal_4566) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_1944), .Q (new_AGEMA_signal_4568) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n15), .Q (new_AGEMA_signal_4570) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_1948), .Q (new_AGEMA_signal_4572) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_3177), .Q (new_AGEMA_signal_4574) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_3179), .Q (new_AGEMA_signal_4576) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n6), .Q (new_AGEMA_signal_4578) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_1950), .Q (new_AGEMA_signal_4580) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n15), .Q (new_AGEMA_signal_4582) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_1954), .Q (new_AGEMA_signal_4584) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_3193), .Q (new_AGEMA_signal_4586) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_3195), .Q (new_AGEMA_signal_4588) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n6), .Q (new_AGEMA_signal_4590) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_1956), .Q (new_AGEMA_signal_4592) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n15), .Q (new_AGEMA_signal_4594) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_1960), .Q (new_AGEMA_signal_4596) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_3209), .Q (new_AGEMA_signal_4598) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_3211), .Q (new_AGEMA_signal_4600) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n6), .Q (new_AGEMA_signal_4602) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_1962), .Q (new_AGEMA_signal_4604) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n15), .Q (new_AGEMA_signal_4606) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_1966), .Q (new_AGEMA_signal_4608) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_3225), .Q (new_AGEMA_signal_4610) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_3227), .Q (new_AGEMA_signal_4612) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n6), .Q (new_AGEMA_signal_4614) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_1968), .Q (new_AGEMA_signal_4616) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n15), .Q (new_AGEMA_signal_4618) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_1972), .Q (new_AGEMA_signal_4620) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_3241), .Q (new_AGEMA_signal_4622) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_3243), .Q (new_AGEMA_signal_4624) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n6), .Q (new_AGEMA_signal_4626) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_1974), .Q (new_AGEMA_signal_4628) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n15), .Q (new_AGEMA_signal_4630) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_1978), .Q (new_AGEMA_signal_4632) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_3257), .Q (new_AGEMA_signal_4634) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_3259), .Q (new_AGEMA_signal_4636) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n6), .Q (new_AGEMA_signal_4638) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_1980), .Q (new_AGEMA_signal_4640) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n15), .Q (new_AGEMA_signal_4642) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_1984), .Q (new_AGEMA_signal_4644) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_3273), .Q (new_AGEMA_signal_4646) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_3275), .Q (new_AGEMA_signal_4648) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n6), .Q (new_AGEMA_signal_4650) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_1986), .Q (new_AGEMA_signal_4652) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n15), .Q (new_AGEMA_signal_4654) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_1990), .Q (new_AGEMA_signal_4656) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C (clk), .D (new_AGEMA_signal_3289), .Q (new_AGEMA_signal_4658) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_3291), .Q (new_AGEMA_signal_4660) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n6), .Q (new_AGEMA_signal_4662) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_1992), .Q (new_AGEMA_signal_4664) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n15), .Q (new_AGEMA_signal_4666) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_1996), .Q (new_AGEMA_signal_4668) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_3305), .Q (new_AGEMA_signal_4670) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_3307), .Q (new_AGEMA_signal_4672) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n6), .Q (new_AGEMA_signal_4674) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_1998), .Q (new_AGEMA_signal_4676) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n15), .Q (new_AGEMA_signal_4678) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_2002), .Q (new_AGEMA_signal_4680) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C (clk), .D (new_AGEMA_signal_3321), .Q (new_AGEMA_signal_4682) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_3323), .Q (new_AGEMA_signal_4684) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n6), .Q (new_AGEMA_signal_4686) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_2004), .Q (new_AGEMA_signal_4688) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n15), .Q (new_AGEMA_signal_4690) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_4692) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_3337), .Q (new_AGEMA_signal_4694) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_3339), .Q (new_AGEMA_signal_4696) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n6), .Q (new_AGEMA_signal_4698) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_2010), .Q (new_AGEMA_signal_4700) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_4704) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_4709), .Q (new_AGEMA_signal_4710) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_4717), .Q (new_AGEMA_signal_4718) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_4725), .Q (new_AGEMA_signal_4726) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_4733), .Q (new_AGEMA_signal_4734) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_4741), .Q (new_AGEMA_signal_4742) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_4749), .Q (new_AGEMA_signal_4750) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_4757), .Q (new_AGEMA_signal_4758) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_4765), .Q (new_AGEMA_signal_4766) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_4773), .Q (new_AGEMA_signal_4774) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_4781), .Q (new_AGEMA_signal_4782) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_4789), .Q (new_AGEMA_signal_4790) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_4797), .Q (new_AGEMA_signal_4798) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_4805), .Q (new_AGEMA_signal_4806) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_4813), .Q (new_AGEMA_signal_4814) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_4821), .Q (new_AGEMA_signal_4822) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_4829), .Q (new_AGEMA_signal_4830) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_4837), .Q (new_AGEMA_signal_4838) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_4845), .Q (new_AGEMA_signal_4846) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C (clk), .D (new_AGEMA_signal_4853), .Q (new_AGEMA_signal_4854) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C (clk), .D (new_AGEMA_signal_4861), .Q (new_AGEMA_signal_4862) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C (clk), .D (new_AGEMA_signal_4869), .Q (new_AGEMA_signal_4870) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C (clk), .D (new_AGEMA_signal_4877), .Q (new_AGEMA_signal_4878) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C (clk), .D (new_AGEMA_signal_4885), .Q (new_AGEMA_signal_4886) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C (clk), .D (new_AGEMA_signal_4893), .Q (new_AGEMA_signal_4894) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C (clk), .D (new_AGEMA_signal_4901), .Q (new_AGEMA_signal_4902) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C (clk), .D (new_AGEMA_signal_4909), .Q (new_AGEMA_signal_4910) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C (clk), .D (new_AGEMA_signal_4917), .Q (new_AGEMA_signal_4918) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C (clk), .D (new_AGEMA_signal_4925), .Q (new_AGEMA_signal_4926) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C (clk), .D (new_AGEMA_signal_4933), .Q (new_AGEMA_signal_4934) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C (clk), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_4942) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C (clk), .D (new_AGEMA_signal_4949), .Q (new_AGEMA_signal_4950) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C (clk), .D (new_AGEMA_signal_4957), .Q (new_AGEMA_signal_4958) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C (clk), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_4966) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C (clk), .D (new_AGEMA_signal_4973), .Q (new_AGEMA_signal_4974) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C (clk), .D (new_AGEMA_signal_4981), .Q (new_AGEMA_signal_4982) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C (clk), .D (new_AGEMA_signal_4989), .Q (new_AGEMA_signal_4990) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C (clk), .D (new_AGEMA_signal_4997), .Q (new_AGEMA_signal_4998) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C (clk), .D (new_AGEMA_signal_5005), .Q (new_AGEMA_signal_5006) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_5014) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C (clk), .D (new_AGEMA_signal_5021), .Q (new_AGEMA_signal_5022) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C (clk), .D (new_AGEMA_signal_5029), .Q (new_AGEMA_signal_5030) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C (clk), .D (new_AGEMA_signal_5037), .Q (new_AGEMA_signal_5038) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C (clk), .D (new_AGEMA_signal_5045), .Q (new_AGEMA_signal_5046) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C (clk), .D (new_AGEMA_signal_5053), .Q (new_AGEMA_signal_5054) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C (clk), .D (new_AGEMA_signal_5061), .Q (new_AGEMA_signal_5062) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C (clk), .D (new_AGEMA_signal_5069), .Q (new_AGEMA_signal_5070) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C (clk), .D (new_AGEMA_signal_5077), .Q (new_AGEMA_signal_5078) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_5086) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C (clk), .D (new_AGEMA_signal_5093), .Q (new_AGEMA_signal_5094) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C (clk), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_5102) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C (clk), .D (new_AGEMA_signal_5109), .Q (new_AGEMA_signal_5110) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C (clk), .D (new_AGEMA_signal_5117), .Q (new_AGEMA_signal_5118) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C (clk), .D (new_AGEMA_signal_5125), .Q (new_AGEMA_signal_5126) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_5134) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C (clk), .D (new_AGEMA_signal_5141), .Q (new_AGEMA_signal_5142) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C (clk), .D (new_AGEMA_signal_5149), .Q (new_AGEMA_signal_5150) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_5158) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C (clk), .D (new_AGEMA_signal_5165), .Q (new_AGEMA_signal_5166) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_5174) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C (clk), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_5182) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C (clk), .D (new_AGEMA_signal_5189), .Q (new_AGEMA_signal_5190) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C (clk), .D (new_AGEMA_signal_5197), .Q (new_AGEMA_signal_5198) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_5206) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C (clk), .D (new_AGEMA_signal_5213), .Q (new_AGEMA_signal_5214) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C (clk), .D (new_AGEMA_signal_5221), .Q (new_AGEMA_signal_5222) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_5230) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C (clk), .D (new_AGEMA_signal_5237), .Q (new_AGEMA_signal_5238) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C (clk), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_5246) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C (clk), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_5254) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C (clk), .D (new_AGEMA_signal_5261), .Q (new_AGEMA_signal_5262) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C (clk), .D (new_AGEMA_signal_5269), .Q (new_AGEMA_signal_5270) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C (clk), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_5278) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C (clk), .D (new_AGEMA_signal_5285), .Q (new_AGEMA_signal_5286) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C (clk), .D (new_AGEMA_signal_5293), .Q (new_AGEMA_signal_5294) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C (clk), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_5302) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C (clk), .D (new_AGEMA_signal_5309), .Q (new_AGEMA_signal_5310) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_5318) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C (clk), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_5326) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C (clk), .D (new_AGEMA_signal_5333), .Q (new_AGEMA_signal_5334) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C (clk), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_5342) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C (clk), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_5350) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C (clk), .D (new_AGEMA_signal_5357), .Q (new_AGEMA_signal_5358) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C (clk), .D (new_AGEMA_signal_5365), .Q (new_AGEMA_signal_5366) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C (clk), .D (new_AGEMA_signal_5373), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C (clk), .D (new_AGEMA_signal_5381), .Q (new_AGEMA_signal_5382) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C (clk), .D (new_AGEMA_signal_5389), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C (clk), .D (new_AGEMA_signal_5397), .Q (new_AGEMA_signal_5398) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C (clk), .D (new_AGEMA_signal_5405), .Q (new_AGEMA_signal_5406) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C (clk), .D (new_AGEMA_signal_5413), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C (clk), .D (new_AGEMA_signal_5421), .Q (new_AGEMA_signal_5422) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C (clk), .D (new_AGEMA_signal_5429), .Q (new_AGEMA_signal_5430) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C (clk), .D (new_AGEMA_signal_5437), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C (clk), .D (new_AGEMA_signal_5445), .Q (new_AGEMA_signal_5446) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C (clk), .D (new_AGEMA_signal_5453), .Q (new_AGEMA_signal_5454) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C (clk), .D (new_AGEMA_signal_5461), .Q (new_AGEMA_signal_5462) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C (clk), .D (new_AGEMA_signal_5469), .Q (new_AGEMA_signal_5470) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C (clk), .D (new_AGEMA_signal_5477), .Q (new_AGEMA_signal_5478) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C (clk), .D (new_AGEMA_signal_5485), .Q (new_AGEMA_signal_5486) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C (clk), .D (new_AGEMA_signal_5493), .Q (new_AGEMA_signal_5494) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C (clk), .D (new_AGEMA_signal_5501), .Q (new_AGEMA_signal_5502) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C (clk), .D (new_AGEMA_signal_5509), .Q (new_AGEMA_signal_5510) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C (clk), .D (new_AGEMA_signal_5517), .Q (new_AGEMA_signal_5518) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C (clk), .D (new_AGEMA_signal_5525), .Q (new_AGEMA_signal_5526) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C (clk), .D (new_AGEMA_signal_5533), .Q (new_AGEMA_signal_5534) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C (clk), .D (new_AGEMA_signal_5541), .Q (new_AGEMA_signal_5542) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C (clk), .D (new_AGEMA_signal_5549), .Q (new_AGEMA_signal_5550) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C (clk), .D (new_AGEMA_signal_5557), .Q (new_AGEMA_signal_5558) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C (clk), .D (new_AGEMA_signal_5565), .Q (new_AGEMA_signal_5566) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C (clk), .D (new_AGEMA_signal_5573), .Q (new_AGEMA_signal_5574) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C (clk), .D (new_AGEMA_signal_5581), .Q (new_AGEMA_signal_5582) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C (clk), .D (new_AGEMA_signal_5589), .Q (new_AGEMA_signal_5590) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C (clk), .D (new_AGEMA_signal_5597), .Q (new_AGEMA_signal_5598) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C (clk), .D (new_AGEMA_signal_5605), .Q (new_AGEMA_signal_5606) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C (clk), .D (new_AGEMA_signal_5613), .Q (new_AGEMA_signal_5614) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C (clk), .D (new_AGEMA_signal_5621), .Q (new_AGEMA_signal_5622) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C (clk), .D (new_AGEMA_signal_5629), .Q (new_AGEMA_signal_5630) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C (clk), .D (new_AGEMA_signal_5637), .Q (new_AGEMA_signal_5638) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C (clk), .D (new_AGEMA_signal_5645), .Q (new_AGEMA_signal_5646) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C (clk), .D (new_AGEMA_signal_5653), .Q (new_AGEMA_signal_5654) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C (clk), .D (new_AGEMA_signal_5661), .Q (new_AGEMA_signal_5662) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C (clk), .D (new_AGEMA_signal_5669), .Q (new_AGEMA_signal_5670) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C (clk), .D (new_AGEMA_signal_5677), .Q (new_AGEMA_signal_5678) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C (clk), .D (new_AGEMA_signal_5685), .Q (new_AGEMA_signal_5686) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C (clk), .D (new_AGEMA_signal_5693), .Q (new_AGEMA_signal_5694) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C (clk), .D (new_AGEMA_signal_5701), .Q (new_AGEMA_signal_5702) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C (clk), .D (new_AGEMA_signal_5709), .Q (new_AGEMA_signal_5710) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C (clk), .D (new_AGEMA_signal_5717), .Q (new_AGEMA_signal_5718) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C (clk), .D (new_AGEMA_signal_5725), .Q (new_AGEMA_signal_5726) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_5736) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_5744) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_5752) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_5760) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_5784) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_5792) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_5832) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_5840) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_5880) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_5888) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_5904) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_5912) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_5952) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_5960) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_6000) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_6008) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_6048) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_6055), .Q (new_AGEMA_signal_6056) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_6072) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_6079), .Q (new_AGEMA_signal_6080) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_6120) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_6128) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_6168) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_6176) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_6216) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_6224) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_6239), .Q (new_AGEMA_signal_6240) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_0_n13), .Q (new_AGEMA_signal_6250) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_1922), .Q (new_AGEMA_signal_6254) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_1_n13), .Q (new_AGEMA_signal_6262) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_6266) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_2_n13), .Q (new_AGEMA_signal_6274) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_1934), .Q (new_AGEMA_signal_6278) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_3_n13), .Q (new_AGEMA_signal_6286) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C (clk), .D (new_AGEMA_signal_1940), .Q (new_AGEMA_signal_6290) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_4_n13), .Q (new_AGEMA_signal_6298) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_6302) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_5_n13), .Q (new_AGEMA_signal_6310) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C (clk), .D (new_AGEMA_signal_1952), .Q (new_AGEMA_signal_6314) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_6_n13), .Q (new_AGEMA_signal_6322) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_1958), .Q (new_AGEMA_signal_6326) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_7_n13), .Q (new_AGEMA_signal_6334) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C (clk), .D (new_AGEMA_signal_1964), .Q (new_AGEMA_signal_6338) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_8_n13), .Q (new_AGEMA_signal_6346) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_1970), .Q (new_AGEMA_signal_6350) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_9_n13), .Q (new_AGEMA_signal_6358) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C (clk), .D (new_AGEMA_signal_1976), .Q (new_AGEMA_signal_6362) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_10_n13), .Q (new_AGEMA_signal_6370) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_1982), .Q (new_AGEMA_signal_6374) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_11_n13), .Q (new_AGEMA_signal_6382) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C (clk), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_6386) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_12_n13), .Q (new_AGEMA_signal_6394) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C (clk), .D (new_AGEMA_signal_1994), .Q (new_AGEMA_signal_6398) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_13_n13), .Q (new_AGEMA_signal_6406) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C (clk), .D (new_AGEMA_signal_2000), .Q (new_AGEMA_signal_6410) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_14_n13), .Q (new_AGEMA_signal_6418) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C (clk), .D (new_AGEMA_signal_2006), .Q (new_AGEMA_signal_6422) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C (clk), .D (Midori_rounds_sub_sBox_PRINCE_15_n13), .Q (new_AGEMA_signal_6430) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C (clk), .D (new_AGEMA_signal_2012), .Q (new_AGEMA_signal_6434) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C (clk), .D (new_AGEMA_signal_6441), .Q (new_AGEMA_signal_6442) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C (clk), .D (new_AGEMA_signal_6449), .Q (new_AGEMA_signal_6450) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C (clk), .D (new_AGEMA_signal_6457), .Q (new_AGEMA_signal_6458) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C (clk), .D (new_AGEMA_signal_6465), .Q (new_AGEMA_signal_6466) ) ;

    /* cells in depth 4 */
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .a ({new_AGEMA_signal_1922, Midori_rounds_sub_sBox_PRINCE_0_n13}), .b ({new_AGEMA_signal_3099, new_AGEMA_signal_3097}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_2065, Midori_rounds_sub_sBox_PRINCE_0_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .a ({new_AGEMA_signal_1663, Midori_rounds_sub_sBox_PRINCE_0_n10}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3101}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_1917, Midori_rounds_sub_sBox_PRINCE_0_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3105}), .b ({new_AGEMA_signal_1919, Midori_rounds_sub_sBox_PRINCE_0_n4}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_2067, Midori_rounds_sub_sBox_PRINCE_0_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3109}), .b ({new_AGEMA_signal_1665, Midori_rounds_sub_sBox_PRINCE_0_n1}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_1921, Midori_rounds_sub_sBox_PRINCE_0_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .a ({new_AGEMA_signal_1928, Midori_rounds_sub_sBox_PRINCE_1_n13}), .b ({new_AGEMA_signal_3115, new_AGEMA_signal_3113}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_1_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .a ({new_AGEMA_signal_1671, Midori_rounds_sub_sBox_PRINCE_1_n10}), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3117}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_1923, Midori_rounds_sub_sBox_PRINCE_1_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3121}), .b ({new_AGEMA_signal_1925, Midori_rounds_sub_sBox_PRINCE_1_n4}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_1_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .a ({new_AGEMA_signal_3127, new_AGEMA_signal_3125}), .b ({new_AGEMA_signal_1673, Midori_rounds_sub_sBox_PRINCE_1_n1}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_1927, Midori_rounds_sub_sBox_PRINCE_1_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .a ({new_AGEMA_signal_1934, Midori_rounds_sub_sBox_PRINCE_2_n13}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3129}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_2075, Midori_rounds_sub_sBox_PRINCE_2_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .a ({new_AGEMA_signal_1679, Midori_rounds_sub_sBox_PRINCE_2_n10}), .b ({new_AGEMA_signal_3135, new_AGEMA_signal_3133}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_1929, Midori_rounds_sub_sBox_PRINCE_2_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3137}), .b ({new_AGEMA_signal_1931, Midori_rounds_sub_sBox_PRINCE_2_n4}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_2077, Midori_rounds_sub_sBox_PRINCE_2_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .a ({new_AGEMA_signal_3143, new_AGEMA_signal_3141}), .b ({new_AGEMA_signal_1681, Midori_rounds_sub_sBox_PRINCE_2_n1}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_1933, Midori_rounds_sub_sBox_PRINCE_2_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .a ({new_AGEMA_signal_1940, Midori_rounds_sub_sBox_PRINCE_3_n13}), .b ({new_AGEMA_signal_3147, new_AGEMA_signal_3145}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_2080, Midori_rounds_sub_sBox_PRINCE_3_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .a ({new_AGEMA_signal_1687, Midori_rounds_sub_sBox_PRINCE_3_n10}), .b ({new_AGEMA_signal_3151, new_AGEMA_signal_3149}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_1935, Midori_rounds_sub_sBox_PRINCE_3_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3153}), .b ({new_AGEMA_signal_1937, Midori_rounds_sub_sBox_PRINCE_3_n4}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_3_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3157}), .b ({new_AGEMA_signal_1689, Midori_rounds_sub_sBox_PRINCE_3_n1}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_1939, Midori_rounds_sub_sBox_PRINCE_3_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .a ({new_AGEMA_signal_1946, Midori_rounds_sub_sBox_PRINCE_4_n13}), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3161}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_2085, Midori_rounds_sub_sBox_PRINCE_4_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .a ({new_AGEMA_signal_1695, Midori_rounds_sub_sBox_PRINCE_4_n10}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3165}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_1941, Midori_rounds_sub_sBox_PRINCE_4_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3169}), .b ({new_AGEMA_signal_1943, Midori_rounds_sub_sBox_PRINCE_4_n4}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_2087, Midori_rounds_sub_sBox_PRINCE_4_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3173}), .b ({new_AGEMA_signal_1697, Midori_rounds_sub_sBox_PRINCE_4_n1}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_1945, Midori_rounds_sub_sBox_PRINCE_4_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .a ({new_AGEMA_signal_1952, Midori_rounds_sub_sBox_PRINCE_5_n13}), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3177}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_2090, Midori_rounds_sub_sBox_PRINCE_5_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .a ({new_AGEMA_signal_1703, Midori_rounds_sub_sBox_PRINCE_5_n10}), .b ({new_AGEMA_signal_3183, new_AGEMA_signal_3181}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_1947, Midori_rounds_sub_sBox_PRINCE_5_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3185}), .b ({new_AGEMA_signal_1949, Midori_rounds_sub_sBox_PRINCE_5_n4}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_2092, Midori_rounds_sub_sBox_PRINCE_5_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3189}), .b ({new_AGEMA_signal_1705, Midori_rounds_sub_sBox_PRINCE_5_n1}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_1951, Midori_rounds_sub_sBox_PRINCE_5_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .a ({new_AGEMA_signal_1958, Midori_rounds_sub_sBox_PRINCE_6_n13}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3193}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_2095, Midori_rounds_sub_sBox_PRINCE_6_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .a ({new_AGEMA_signal_1711, Midori_rounds_sub_sBox_PRINCE_6_n10}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3197}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_1953, Midori_rounds_sub_sBox_PRINCE_6_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3201}), .b ({new_AGEMA_signal_1955, Midori_rounds_sub_sBox_PRINCE_6_n4}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_2097, Midori_rounds_sub_sBox_PRINCE_6_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .a ({new_AGEMA_signal_3207, new_AGEMA_signal_3205}), .b ({new_AGEMA_signal_1713, Midori_rounds_sub_sBox_PRINCE_6_n1}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_1957, Midori_rounds_sub_sBox_PRINCE_6_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .a ({new_AGEMA_signal_1964, Midori_rounds_sub_sBox_PRINCE_7_n13}), .b ({new_AGEMA_signal_3211, new_AGEMA_signal_3209}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_7_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .a ({new_AGEMA_signal_1719, Midori_rounds_sub_sBox_PRINCE_7_n10}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3213}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_1959, Midori_rounds_sub_sBox_PRINCE_7_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3217}), .b ({new_AGEMA_signal_1961, Midori_rounds_sub_sBox_PRINCE_7_n4}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_7_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .a ({new_AGEMA_signal_3223, new_AGEMA_signal_3221}), .b ({new_AGEMA_signal_1721, Midori_rounds_sub_sBox_PRINCE_7_n1}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_1963, Midori_rounds_sub_sBox_PRINCE_7_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .a ({new_AGEMA_signal_1970, Midori_rounds_sub_sBox_PRINCE_8_n13}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3225}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_2105, Midori_rounds_sub_sBox_PRINCE_8_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .a ({new_AGEMA_signal_1727, Midori_rounds_sub_sBox_PRINCE_8_n10}), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3229}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_1965, Midori_rounds_sub_sBox_PRINCE_8_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3233}), .b ({new_AGEMA_signal_1967, Midori_rounds_sub_sBox_PRINCE_8_n4}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_2107, Midori_rounds_sub_sBox_PRINCE_8_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3237}), .b ({new_AGEMA_signal_1729, Midori_rounds_sub_sBox_PRINCE_8_n1}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_1969, Midori_rounds_sub_sBox_PRINCE_8_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .a ({new_AGEMA_signal_1976, Midori_rounds_sub_sBox_PRINCE_9_n13}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3241}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_9_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .a ({new_AGEMA_signal_1735, Midori_rounds_sub_sBox_PRINCE_9_n10}), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3245}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_1971, Midori_rounds_sub_sBox_PRINCE_9_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3249}), .b ({new_AGEMA_signal_1973, Midori_rounds_sub_sBox_PRINCE_9_n4}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_2112, Midori_rounds_sub_sBox_PRINCE_9_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .a ({new_AGEMA_signal_3255, new_AGEMA_signal_3253}), .b ({new_AGEMA_signal_1737, Midori_rounds_sub_sBox_PRINCE_9_n1}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_1975, Midori_rounds_sub_sBox_PRINCE_9_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .a ({new_AGEMA_signal_1982, Midori_rounds_sub_sBox_PRINCE_10_n13}), .b ({new_AGEMA_signal_3259, new_AGEMA_signal_3257}), .clk (clk), .r (Fresh[136]), .c ({new_AGEMA_signal_2115, Midori_rounds_sub_sBox_PRINCE_10_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .a ({new_AGEMA_signal_1743, Midori_rounds_sub_sBox_PRINCE_10_n10}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3261}), .clk (clk), .r (Fresh[137]), .c ({new_AGEMA_signal_1977, Midori_rounds_sub_sBox_PRINCE_10_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3265}), .b ({new_AGEMA_signal_1979, Midori_rounds_sub_sBox_PRINCE_10_n4}), .clk (clk), .r (Fresh[138]), .c ({new_AGEMA_signal_2117, Midori_rounds_sub_sBox_PRINCE_10_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3269}), .b ({new_AGEMA_signal_1745, Midori_rounds_sub_sBox_PRINCE_10_n1}), .clk (clk), .r (Fresh[139]), .c ({new_AGEMA_signal_1981, Midori_rounds_sub_sBox_PRINCE_10_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .a ({new_AGEMA_signal_1988, Midori_rounds_sub_sBox_PRINCE_11_n13}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3273}), .clk (clk), .r (Fresh[140]), .c ({new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_11_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .a ({new_AGEMA_signal_1751, Midori_rounds_sub_sBox_PRINCE_11_n10}), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3277}), .clk (clk), .r (Fresh[141]), .c ({new_AGEMA_signal_1983, Midori_rounds_sub_sBox_PRINCE_11_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .a ({new_AGEMA_signal_3283, new_AGEMA_signal_3281}), .b ({new_AGEMA_signal_1985, Midori_rounds_sub_sBox_PRINCE_11_n4}), .clk (clk), .r (Fresh[142]), .c ({new_AGEMA_signal_2122, Midori_rounds_sub_sBox_PRINCE_11_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .a ({new_AGEMA_signal_3287, new_AGEMA_signal_3285}), .b ({new_AGEMA_signal_1753, Midori_rounds_sub_sBox_PRINCE_11_n1}), .clk (clk), .r (Fresh[143]), .c ({new_AGEMA_signal_1987, Midori_rounds_sub_sBox_PRINCE_11_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .a ({new_AGEMA_signal_1994, Midori_rounds_sub_sBox_PRINCE_12_n13}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3289}), .clk (clk), .r (Fresh[144]), .c ({new_AGEMA_signal_2125, Midori_rounds_sub_sBox_PRINCE_12_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .a ({new_AGEMA_signal_1759, Midori_rounds_sub_sBox_PRINCE_12_n10}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3293}), .clk (clk), .r (Fresh[145]), .c ({new_AGEMA_signal_1989, Midori_rounds_sub_sBox_PRINCE_12_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .a ({new_AGEMA_signal_3299, new_AGEMA_signal_3297}), .b ({new_AGEMA_signal_1991, Midori_rounds_sub_sBox_PRINCE_12_n4}), .clk (clk), .r (Fresh[146]), .c ({new_AGEMA_signal_2127, Midori_rounds_sub_sBox_PRINCE_12_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .a ({new_AGEMA_signal_3303, new_AGEMA_signal_3301}), .b ({new_AGEMA_signal_1761, Midori_rounds_sub_sBox_PRINCE_12_n1}), .clk (clk), .r (Fresh[147]), .c ({new_AGEMA_signal_1993, Midori_rounds_sub_sBox_PRINCE_12_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .a ({new_AGEMA_signal_2000, Midori_rounds_sub_sBox_PRINCE_13_n13}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3305}), .clk (clk), .r (Fresh[148]), .c ({new_AGEMA_signal_2130, Midori_rounds_sub_sBox_PRINCE_13_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .a ({new_AGEMA_signal_1767, Midori_rounds_sub_sBox_PRINCE_13_n10}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3309}), .clk (clk), .r (Fresh[149]), .c ({new_AGEMA_signal_1995, Midori_rounds_sub_sBox_PRINCE_13_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .a ({new_AGEMA_signal_3315, new_AGEMA_signal_3313}), .b ({new_AGEMA_signal_1997, Midori_rounds_sub_sBox_PRINCE_13_n4}), .clk (clk), .r (Fresh[150]), .c ({new_AGEMA_signal_2132, Midori_rounds_sub_sBox_PRINCE_13_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .a ({new_AGEMA_signal_3319, new_AGEMA_signal_3317}), .b ({new_AGEMA_signal_1769, Midori_rounds_sub_sBox_PRINCE_13_n1}), .clk (clk), .r (Fresh[151]), .c ({new_AGEMA_signal_1999, Midori_rounds_sub_sBox_PRINCE_13_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .a ({new_AGEMA_signal_2006, Midori_rounds_sub_sBox_PRINCE_14_n13}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3321}), .clk (clk), .r (Fresh[152]), .c ({new_AGEMA_signal_2135, Midori_rounds_sub_sBox_PRINCE_14_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .a ({new_AGEMA_signal_1775, Midori_rounds_sub_sBox_PRINCE_14_n10}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3325}), .clk (clk), .r (Fresh[153]), .c ({new_AGEMA_signal_2001, Midori_rounds_sub_sBox_PRINCE_14_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3329}), .b ({new_AGEMA_signal_2003, Midori_rounds_sub_sBox_PRINCE_14_n4}), .clk (clk), .r (Fresh[154]), .c ({new_AGEMA_signal_2137, Midori_rounds_sub_sBox_PRINCE_14_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3333}), .b ({new_AGEMA_signal_1777, Midori_rounds_sub_sBox_PRINCE_14_n1}), .clk (clk), .r (Fresh[155]), .c ({new_AGEMA_signal_2005, Midori_rounds_sub_sBox_PRINCE_14_n2}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .a ({new_AGEMA_signal_2012, Midori_rounds_sub_sBox_PRINCE_15_n13}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3337}), .clk (clk), .r (Fresh[156]), .c ({new_AGEMA_signal_2140, Midori_rounds_sub_sBox_PRINCE_15_n14}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .a ({new_AGEMA_signal_1783, Midori_rounds_sub_sBox_PRINCE_15_n10}), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3341}), .clk (clk), .r (Fresh[157]), .c ({new_AGEMA_signal_2007, Midori_rounds_sub_sBox_PRINCE_15_n11}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3345}), .b ({new_AGEMA_signal_2009, Midori_rounds_sub_sBox_PRINCE_15_n4}), .clk (clk), .r (Fresh[158]), .c ({new_AGEMA_signal_2142, Midori_rounds_sub_sBox_PRINCE_15_n5}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3349}), .b ({new_AGEMA_signal_1785, Midori_rounds_sub_sBox_PRINCE_15_n1}), .clk (clk), .r (Fresh[159]), .c ({new_AGEMA_signal_2011, Midori_rounds_sub_sBox_PRINCE_15_n2}) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (new_AGEMA_signal_3027), .Q (new_AGEMA_signal_3028) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (clk), .D (new_AGEMA_signal_3354), .Q (new_AGEMA_signal_3355) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (clk), .D (new_AGEMA_signal_3360), .Q (new_AGEMA_signal_3361) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (clk), .D (new_AGEMA_signal_3366), .Q (new_AGEMA_signal_3367) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (clk), .D (new_AGEMA_signal_3372), .Q (new_AGEMA_signal_3373) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (clk), .D (new_AGEMA_signal_3378), .Q (new_AGEMA_signal_3379) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (clk), .D (new_AGEMA_signal_3384), .Q (new_AGEMA_signal_3385) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (clk), .D (new_AGEMA_signal_3390), .Q (new_AGEMA_signal_3391) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (clk), .D (new_AGEMA_signal_3396), .Q (new_AGEMA_signal_3397) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (clk), .D (new_AGEMA_signal_3402), .Q (new_AGEMA_signal_3403) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (clk), .D (new_AGEMA_signal_3408), .Q (new_AGEMA_signal_3409) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (clk), .D (new_AGEMA_signal_3414), .Q (new_AGEMA_signal_3415) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (clk), .D (new_AGEMA_signal_3420), .Q (new_AGEMA_signal_3421) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (clk), .D (new_AGEMA_signal_3426), .Q (new_AGEMA_signal_3427) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (clk), .D (new_AGEMA_signal_3432), .Q (new_AGEMA_signal_3433) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (clk), .D (new_AGEMA_signal_3438), .Q (new_AGEMA_signal_3439) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (clk), .D (new_AGEMA_signal_3444), .Q (new_AGEMA_signal_3445) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (clk), .D (new_AGEMA_signal_3450), .Q (new_AGEMA_signal_3451) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (clk), .D (new_AGEMA_signal_3456), .Q (new_AGEMA_signal_3457) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (clk), .D (new_AGEMA_signal_3462), .Q (new_AGEMA_signal_3463) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (clk), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_3469) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (clk), .D (new_AGEMA_signal_3474), .Q (new_AGEMA_signal_3475) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (clk), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_3481) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (clk), .D (new_AGEMA_signal_3486), .Q (new_AGEMA_signal_3487) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (clk), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_3493) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (clk), .D (new_AGEMA_signal_3498), .Q (new_AGEMA_signal_3499) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (clk), .D (new_AGEMA_signal_3504), .Q (new_AGEMA_signal_3505) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (clk), .D (new_AGEMA_signal_3510), .Q (new_AGEMA_signal_3511) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (clk), .D (new_AGEMA_signal_3516), .Q (new_AGEMA_signal_3517) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (clk), .D (new_AGEMA_signal_3522), .Q (new_AGEMA_signal_3523) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (clk), .D (new_AGEMA_signal_3528), .Q (new_AGEMA_signal_3529) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (clk), .D (new_AGEMA_signal_3534), .Q (new_AGEMA_signal_3535) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (clk), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_3541) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (clk), .D (new_AGEMA_signal_3546), .Q (new_AGEMA_signal_3547) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (clk), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_3553) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (clk), .D (new_AGEMA_signal_3558), .Q (new_AGEMA_signal_3559) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (clk), .D (new_AGEMA_signal_3564), .Q (new_AGEMA_signal_3565) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (clk), .D (new_AGEMA_signal_3570), .Q (new_AGEMA_signal_3571) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (clk), .D (new_AGEMA_signal_3576), .Q (new_AGEMA_signal_3577) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (clk), .D (new_AGEMA_signal_3582), .Q (new_AGEMA_signal_3583) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (clk), .D (new_AGEMA_signal_3588), .Q (new_AGEMA_signal_3589) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (clk), .D (new_AGEMA_signal_3594), .Q (new_AGEMA_signal_3595) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (clk), .D (new_AGEMA_signal_3600), .Q (new_AGEMA_signal_3601) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (clk), .D (new_AGEMA_signal_3606), .Q (new_AGEMA_signal_3607) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (clk), .D (new_AGEMA_signal_3612), .Q (new_AGEMA_signal_3613) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (clk), .D (new_AGEMA_signal_3618), .Q (new_AGEMA_signal_3619) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (clk), .D (new_AGEMA_signal_3624), .Q (new_AGEMA_signal_3625) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (clk), .D (new_AGEMA_signal_3630), .Q (new_AGEMA_signal_3631) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (clk), .D (new_AGEMA_signal_3636), .Q (new_AGEMA_signal_3637) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (clk), .D (new_AGEMA_signal_3642), .Q (new_AGEMA_signal_3643) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (clk), .D (new_AGEMA_signal_3648), .Q (new_AGEMA_signal_3649) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (clk), .D (new_AGEMA_signal_3654), .Q (new_AGEMA_signal_3655) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (clk), .D (new_AGEMA_signal_3660), .Q (new_AGEMA_signal_3661) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (clk), .D (new_AGEMA_signal_3666), .Q (new_AGEMA_signal_3667) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (clk), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (clk), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (clk), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (clk), .D (new_AGEMA_signal_3690), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (clk), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (clk), .D (new_AGEMA_signal_3702), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (clk), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (clk), .D (new_AGEMA_signal_3714), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (clk), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (clk), .D (new_AGEMA_signal_3726), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (clk), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (clk), .D (new_AGEMA_signal_3738), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (clk), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (clk), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (clk), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_3757) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (clk), .D (new_AGEMA_signal_3762), .Q (new_AGEMA_signal_3763) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_3769) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_3774), .Q (new_AGEMA_signal_3775) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_3780), .Q (new_AGEMA_signal_3781) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_3786), .Q (new_AGEMA_signal_3787) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_3792), .Q (new_AGEMA_signal_3793) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_3798), .Q (new_AGEMA_signal_3799) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_3804), .Q (new_AGEMA_signal_3805) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_3810), .Q (new_AGEMA_signal_3811) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_3817) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_3822), .Q (new_AGEMA_signal_3823) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_3828), .Q (new_AGEMA_signal_3829) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_3834), .Q (new_AGEMA_signal_3835) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_3841) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_3846), .Q (new_AGEMA_signal_3847) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_3853) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_3858), .Q (new_AGEMA_signal_3859) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_3865) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_3870), .Q (new_AGEMA_signal_3871) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_3876), .Q (new_AGEMA_signal_3877) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_3882), .Q (new_AGEMA_signal_3883) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_3889) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_3894), .Q (new_AGEMA_signal_3895) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_3906), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_3930), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_3954), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_3966), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_3978), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_3990), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_4002), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_4008), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_4014), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_4020), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_4026), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_4032), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_4038), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_4044), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_4050), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_4056), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_4062), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_4068), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_4074), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_4080), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_4086), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_4092), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_4098), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_4104), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_4110), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_4116), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_4122), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_4128), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_4134), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_4140), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_4146), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_4152), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_4158), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_4164), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_4170), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_4176), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_4182), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_4188), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_4194), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_4200), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_4206), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_4212), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_4218), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_4224), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_4230), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_4236), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_4242), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_4248), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_4254), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_4260), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_4266), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_4272), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_4278), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_4284), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_4290), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_4296), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_4302), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_4308), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_4314), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_4320), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_4326), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_4332), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_4338), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_4344), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_4350), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_4356), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_4362), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_4368), .Q (new_AGEMA_signal_4369) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_4374), .Q (new_AGEMA_signal_4375) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_4380), .Q (new_AGEMA_signal_4381) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_4386), .Q (new_AGEMA_signal_4387) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_4392), .Q (new_AGEMA_signal_4393) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_4398), .Q (new_AGEMA_signal_4399) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_4404), .Q (new_AGEMA_signal_4405) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_4410), .Q (new_AGEMA_signal_4411) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_4416), .Q (new_AGEMA_signal_4417) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_4422), .Q (new_AGEMA_signal_4423) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_4428), .Q (new_AGEMA_signal_4429) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_4434), .Q (new_AGEMA_signal_4435) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_4440), .Q (new_AGEMA_signal_4441) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_4446), .Q (new_AGEMA_signal_4447) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_4452), .Q (new_AGEMA_signal_4453) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_4458), .Q (new_AGEMA_signal_4459) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_4464), .Q (new_AGEMA_signal_4465) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_4470), .Q (new_AGEMA_signal_4471) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_4476), .Q (new_AGEMA_signal_4477) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_4482), .Q (new_AGEMA_signal_4483) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_4488), .Q (new_AGEMA_signal_4489) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_4494), .Q (new_AGEMA_signal_4495) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_4500), .Q (new_AGEMA_signal_4501) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_4506), .Q (new_AGEMA_signal_4507) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_4510), .Q (new_AGEMA_signal_4511) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_4512), .Q (new_AGEMA_signal_4513) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_4514), .Q (new_AGEMA_signal_4515) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_4516), .Q (new_AGEMA_signal_4517) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_4518), .Q (new_AGEMA_signal_4519) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_4520), .Q (new_AGEMA_signal_4521) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_4522), .Q (new_AGEMA_signal_4523) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_4524), .Q (new_AGEMA_signal_4525) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_4526), .Q (new_AGEMA_signal_4527) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_4528), .Q (new_AGEMA_signal_4529) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_4530), .Q (new_AGEMA_signal_4531) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_4532), .Q (new_AGEMA_signal_4533) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_4534), .Q (new_AGEMA_signal_4535) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_4536), .Q (new_AGEMA_signal_4537) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_4538), .Q (new_AGEMA_signal_4539) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_4540), .Q (new_AGEMA_signal_4541) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_4542), .Q (new_AGEMA_signal_4543) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_4544), .Q (new_AGEMA_signal_4545) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_4546), .Q (new_AGEMA_signal_4547) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_4548), .Q (new_AGEMA_signal_4549) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_4550), .Q (new_AGEMA_signal_4551) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_4552), .Q (new_AGEMA_signal_4553) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_4554), .Q (new_AGEMA_signal_4555) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_4556), .Q (new_AGEMA_signal_4557) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_4558), .Q (new_AGEMA_signal_4559) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_4560), .Q (new_AGEMA_signal_4561) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_4562), .Q (new_AGEMA_signal_4563) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_4564), .Q (new_AGEMA_signal_4565) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_4566), .Q (new_AGEMA_signal_4567) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_4568), .Q (new_AGEMA_signal_4569) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_4570), .Q (new_AGEMA_signal_4571) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_4572), .Q (new_AGEMA_signal_4573) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_4574), .Q (new_AGEMA_signal_4575) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_4576), .Q (new_AGEMA_signal_4577) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_4578), .Q (new_AGEMA_signal_4579) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_4580), .Q (new_AGEMA_signal_4581) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_4582), .Q (new_AGEMA_signal_4583) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_4584), .Q (new_AGEMA_signal_4585) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_4586), .Q (new_AGEMA_signal_4587) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_4588), .Q (new_AGEMA_signal_4589) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_4590), .Q (new_AGEMA_signal_4591) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_4592), .Q (new_AGEMA_signal_4593) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_4594), .Q (new_AGEMA_signal_4595) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_4596), .Q (new_AGEMA_signal_4597) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_4598), .Q (new_AGEMA_signal_4599) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_4600), .Q (new_AGEMA_signal_4601) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_4602), .Q (new_AGEMA_signal_4603) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_4604), .Q (new_AGEMA_signal_4605) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_4606), .Q (new_AGEMA_signal_4607) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_4608), .Q (new_AGEMA_signal_4609) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_4610), .Q (new_AGEMA_signal_4611) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_4612), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_4614), .Q (new_AGEMA_signal_4615) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4617) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_4618), .Q (new_AGEMA_signal_4619) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_4620), .Q (new_AGEMA_signal_4621) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_4623) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_4625) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_4626), .Q (new_AGEMA_signal_4627) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_4628), .Q (new_AGEMA_signal_4629) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_4631) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_4632), .Q (new_AGEMA_signal_4633) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_4634), .Q (new_AGEMA_signal_4635) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_4636), .Q (new_AGEMA_signal_4637) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_4638), .Q (new_AGEMA_signal_4639) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_4641) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_4642), .Q (new_AGEMA_signal_4643) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_4644), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_4646), .Q (new_AGEMA_signal_4647) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_4648), .Q (new_AGEMA_signal_4649) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_4650), .Q (new_AGEMA_signal_4651) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_4652), .Q (new_AGEMA_signal_4653) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_4654), .Q (new_AGEMA_signal_4655) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_4656), .Q (new_AGEMA_signal_4657) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_4658), .Q (new_AGEMA_signal_4659) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_4660), .Q (new_AGEMA_signal_4661) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_4662), .Q (new_AGEMA_signal_4663) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_4664), .Q (new_AGEMA_signal_4665) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_4666), .Q (new_AGEMA_signal_4667) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_4668), .Q (new_AGEMA_signal_4669) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_4670), .Q (new_AGEMA_signal_4671) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_4672), .Q (new_AGEMA_signal_4673) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_4674), .Q (new_AGEMA_signal_4675) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_4676), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_4679) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_4681) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_4683) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_4685) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_4686), .Q (new_AGEMA_signal_4687) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_4689) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_4691) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_4692), .Q (new_AGEMA_signal_4693) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_4695) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_4697) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_4698), .Q (new_AGEMA_signal_4699) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_4701) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_4704), .Q (new_AGEMA_signal_4705) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_4710), .Q (new_AGEMA_signal_4711) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_4719) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_4735) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_4830), .Q (new_AGEMA_signal_4831) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_4855) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_4879) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_4887) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_4895) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_4902), .Q (new_AGEMA_signal_4903) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_4911) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_4919) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_4926), .Q (new_AGEMA_signal_4927) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_4935) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_4943) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_4950), .Q (new_AGEMA_signal_4951) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_4958), .Q (new_AGEMA_signal_4959) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_4967) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_4974), .Q (new_AGEMA_signal_4975) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_4982), .Q (new_AGEMA_signal_4983) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_4991) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_4998), .Q (new_AGEMA_signal_4999) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_5006), .Q (new_AGEMA_signal_5007) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_5015) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_5023) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_5030), .Q (new_AGEMA_signal_5031) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_5039) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_5047) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_5054), .Q (new_AGEMA_signal_5055) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_5063) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_5070), .Q (new_AGEMA_signal_5071) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_5078), .Q (new_AGEMA_signal_5079) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_5087) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_5095) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_5102), .Q (new_AGEMA_signal_5103) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_5111) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_5118), .Q (new_AGEMA_signal_5119) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_5126), .Q (new_AGEMA_signal_5127) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_5135) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_5143) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_5150), .Q (new_AGEMA_signal_5151) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_5159) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_5167) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_5174), .Q (new_AGEMA_signal_5175) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_5183) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_5191) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_5198), .Q (new_AGEMA_signal_5199) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_5207) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_5215) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_5222), .Q (new_AGEMA_signal_5223) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_5231) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_5239) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_5246), .Q (new_AGEMA_signal_5247) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_5255) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_5262), .Q (new_AGEMA_signal_5263) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_5270), .Q (new_AGEMA_signal_5271) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_5279) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_5287) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_5294), .Q (new_AGEMA_signal_5295) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_5303) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_5311) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_5318), .Q (new_AGEMA_signal_5319) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_5326), .Q (new_AGEMA_signal_5327) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_5334), .Q (new_AGEMA_signal_5335) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_5342), .Q (new_AGEMA_signal_5343) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_5350), .Q (new_AGEMA_signal_5351) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_5359) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_5366), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_5383) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_5399) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_5406), .Q (new_AGEMA_signal_5407) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_5414), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_5422), .Q (new_AGEMA_signal_5423) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_5430), .Q (new_AGEMA_signal_5431) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_5446), .Q (new_AGEMA_signal_5447) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_5455) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_5463) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_5471) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_5479) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_5486), .Q (new_AGEMA_signal_5487) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_5495) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_5503) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_5510), .Q (new_AGEMA_signal_5511) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_5519) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_5527) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_5535) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_5543) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_5550), .Q (new_AGEMA_signal_5551) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_5559) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_5566), .Q (new_AGEMA_signal_5567) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_5574), .Q (new_AGEMA_signal_5575) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_5583) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_5591) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_5599) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_5607) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_5615) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_5623) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_5630), .Q (new_AGEMA_signal_5631) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_5639) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_5646), .Q (new_AGEMA_signal_5647) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_5654), .Q (new_AGEMA_signal_5655) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_5663) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_5671) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_5679) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_5687) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_5694), .Q (new_AGEMA_signal_5695) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_5703) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_5711) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_5719) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_5727) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_5849) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_5897) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_5945) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_5993) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_6041) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_6089) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_6136), .Q (new_AGEMA_signal_6137) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_6185) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_6233) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_6251) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_6262), .Q (new_AGEMA_signal_6263) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_6266), .Q (new_AGEMA_signal_6267) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_6275) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_6286), .Q (new_AGEMA_signal_6287) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_6290), .Q (new_AGEMA_signal_6291) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_6298), .Q (new_AGEMA_signal_6299) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_6303) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_6311) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_6314), .Q (new_AGEMA_signal_6315) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_6322), .Q (new_AGEMA_signal_6323) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_6327) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_6335) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_6338), .Q (new_AGEMA_signal_6339) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_6346), .Q (new_AGEMA_signal_6347) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_6351) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_6359) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_6363) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_6370), .Q (new_AGEMA_signal_6371) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_6375) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_6383) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_6387) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_6394), .Q (new_AGEMA_signal_6395) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_6399) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_6407) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_6411) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_6418), .Q (new_AGEMA_signal_6419) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_6423) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_6431) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_6435) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_6442), .Q (new_AGEMA_signal_6443) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_6450), .Q (new_AGEMA_signal_6451) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_6459) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_6466), .Q (new_AGEMA_signal_6467) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_3028), .Q (new_AGEMA_signal_3029) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (clk), .D (new_AGEMA_signal_3355), .Q (new_AGEMA_signal_3356) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (clk), .D (new_AGEMA_signal_3361), .Q (new_AGEMA_signal_3362) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (clk), .D (new_AGEMA_signal_3367), .Q (new_AGEMA_signal_3368) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (clk), .D (new_AGEMA_signal_3373), .Q (new_AGEMA_signal_3374) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (clk), .D (new_AGEMA_signal_3379), .Q (new_AGEMA_signal_3380) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (clk), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_3386) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (clk), .D (new_AGEMA_signal_3391), .Q (new_AGEMA_signal_3392) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (clk), .D (new_AGEMA_signal_3397), .Q (new_AGEMA_signal_3398) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (clk), .D (new_AGEMA_signal_3403), .Q (new_AGEMA_signal_3404) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (clk), .D (new_AGEMA_signal_3409), .Q (new_AGEMA_signal_3410) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (clk), .D (new_AGEMA_signal_3415), .Q (new_AGEMA_signal_3416) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (clk), .D (new_AGEMA_signal_3421), .Q (new_AGEMA_signal_3422) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (clk), .D (new_AGEMA_signal_3427), .Q (new_AGEMA_signal_3428) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (clk), .D (new_AGEMA_signal_3433), .Q (new_AGEMA_signal_3434) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (clk), .D (new_AGEMA_signal_3439), .Q (new_AGEMA_signal_3440) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (clk), .D (new_AGEMA_signal_3445), .Q (new_AGEMA_signal_3446) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (clk), .D (new_AGEMA_signal_3451), .Q (new_AGEMA_signal_3452) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (clk), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_3458) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (clk), .D (new_AGEMA_signal_3463), .Q (new_AGEMA_signal_3464) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (clk), .D (new_AGEMA_signal_3469), .Q (new_AGEMA_signal_3470) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (clk), .D (new_AGEMA_signal_3475), .Q (new_AGEMA_signal_3476) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (clk), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_3482) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (clk), .D (new_AGEMA_signal_3487), .Q (new_AGEMA_signal_3488) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (clk), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_3494) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (clk), .D (new_AGEMA_signal_3499), .Q (new_AGEMA_signal_3500) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (clk), .D (new_AGEMA_signal_3505), .Q (new_AGEMA_signal_3506) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (clk), .D (new_AGEMA_signal_3511), .Q (new_AGEMA_signal_3512) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (clk), .D (new_AGEMA_signal_3517), .Q (new_AGEMA_signal_3518) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (clk), .D (new_AGEMA_signal_3523), .Q (new_AGEMA_signal_3524) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (clk), .D (new_AGEMA_signal_3529), .Q (new_AGEMA_signal_3530) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (clk), .D (new_AGEMA_signal_3535), .Q (new_AGEMA_signal_3536) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (clk), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_3542) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (clk), .D (new_AGEMA_signal_3547), .Q (new_AGEMA_signal_3548) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (clk), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_3554) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (clk), .D (new_AGEMA_signal_3559), .Q (new_AGEMA_signal_3560) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (clk), .D (new_AGEMA_signal_3565), .Q (new_AGEMA_signal_3566) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (clk), .D (new_AGEMA_signal_3571), .Q (new_AGEMA_signal_3572) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (clk), .D (new_AGEMA_signal_3577), .Q (new_AGEMA_signal_3578) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (clk), .D (new_AGEMA_signal_3583), .Q (new_AGEMA_signal_3584) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (clk), .D (new_AGEMA_signal_3589), .Q (new_AGEMA_signal_3590) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (clk), .D (new_AGEMA_signal_3595), .Q (new_AGEMA_signal_3596) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (clk), .D (new_AGEMA_signal_3601), .Q (new_AGEMA_signal_3602) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (clk), .D (new_AGEMA_signal_3607), .Q (new_AGEMA_signal_3608) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (clk), .D (new_AGEMA_signal_3613), .Q (new_AGEMA_signal_3614) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (clk), .D (new_AGEMA_signal_3619), .Q (new_AGEMA_signal_3620) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (clk), .D (new_AGEMA_signal_3625), .Q (new_AGEMA_signal_3626) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (clk), .D (new_AGEMA_signal_3631), .Q (new_AGEMA_signal_3632) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (clk), .D (new_AGEMA_signal_3637), .Q (new_AGEMA_signal_3638) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (clk), .D (new_AGEMA_signal_3643), .Q (new_AGEMA_signal_3644) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (clk), .D (new_AGEMA_signal_3649), .Q (new_AGEMA_signal_3650) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (clk), .D (new_AGEMA_signal_3655), .Q (new_AGEMA_signal_3656) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (clk), .D (new_AGEMA_signal_3661), .Q (new_AGEMA_signal_3662) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (clk), .D (new_AGEMA_signal_3667), .Q (new_AGEMA_signal_3668) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (clk), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (clk), .D (new_AGEMA_signal_3679), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (clk), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (clk), .D (new_AGEMA_signal_3691), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (clk), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (clk), .D (new_AGEMA_signal_3703), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (clk), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (clk), .D (new_AGEMA_signal_3715), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (clk), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (clk), .D (new_AGEMA_signal_3727), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (clk), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (clk), .D (new_AGEMA_signal_3739), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (clk), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (clk), .D (new_AGEMA_signal_3751), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (clk), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_3758) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (clk), .D (new_AGEMA_signal_3763), .Q (new_AGEMA_signal_3764) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (clk), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_3770) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (clk), .D (new_AGEMA_signal_3775), .Q (new_AGEMA_signal_3776) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (clk), .D (new_AGEMA_signal_3781), .Q (new_AGEMA_signal_3782) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (clk), .D (new_AGEMA_signal_3787), .Q (new_AGEMA_signal_3788) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (clk), .D (new_AGEMA_signal_3793), .Q (new_AGEMA_signal_3794) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (clk), .D (new_AGEMA_signal_3799), .Q (new_AGEMA_signal_3800) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (clk), .D (new_AGEMA_signal_3805), .Q (new_AGEMA_signal_3806) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (clk), .D (new_AGEMA_signal_3811), .Q (new_AGEMA_signal_3812) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (clk), .D (new_AGEMA_signal_3817), .Q (new_AGEMA_signal_3818) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (clk), .D (new_AGEMA_signal_3823), .Q (new_AGEMA_signal_3824) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_3829), .Q (new_AGEMA_signal_3830) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (clk), .D (new_AGEMA_signal_3835), .Q (new_AGEMA_signal_3836) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_3841), .Q (new_AGEMA_signal_3842) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (clk), .D (new_AGEMA_signal_3847), .Q (new_AGEMA_signal_3848) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_3853), .Q (new_AGEMA_signal_3854) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (clk), .D (new_AGEMA_signal_3859), .Q (new_AGEMA_signal_3860) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (clk), .D (new_AGEMA_signal_3865), .Q (new_AGEMA_signal_3866) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_3871), .Q (new_AGEMA_signal_3872) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (clk), .D (new_AGEMA_signal_3877), .Q (new_AGEMA_signal_3878) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_3883), .Q (new_AGEMA_signal_3884) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (clk), .D (new_AGEMA_signal_3889), .Q (new_AGEMA_signal_3890) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_3895), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (clk), .D (new_AGEMA_signal_3901), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_3907), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (clk), .D (new_AGEMA_signal_3913), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_3919), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (clk), .D (new_AGEMA_signal_3925), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_3931), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (clk), .D (new_AGEMA_signal_3937), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_3943), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (clk), .D (new_AGEMA_signal_3949), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_3955), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (clk), .D (new_AGEMA_signal_3961), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_3967), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (clk), .D (new_AGEMA_signal_3973), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_3979), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (clk), .D (new_AGEMA_signal_3985), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_3991), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (clk), .D (new_AGEMA_signal_3997), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_4003), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (clk), .D (new_AGEMA_signal_4009), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_4015), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (clk), .D (new_AGEMA_signal_4021), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_4027), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (clk), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_4039), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (clk), .D (new_AGEMA_signal_4045), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_4051), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (clk), .D (new_AGEMA_signal_4057), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_4063), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (clk), .D (new_AGEMA_signal_4069), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_4075), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (clk), .D (new_AGEMA_signal_4081), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_4087), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (clk), .D (new_AGEMA_signal_4093), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_4099), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (clk), .D (new_AGEMA_signal_4105), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_4111), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (clk), .D (new_AGEMA_signal_4117), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_4123), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_4129), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_4135), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_4147), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_4153), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_4159), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_4165), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_4171), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_4183), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_4189), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_4195), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_4207), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_4213), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_4219), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_4225), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_4231), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_4237), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_4243), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_4249), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_4255), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_4261), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_4267), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_4273), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_4279), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_4285), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_4291), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_4297), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_4303), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_4309), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_4315), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_4321), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_4327), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_4333), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_4339), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_4345), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_4351), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_4357), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_4363), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_4369), .Q (new_AGEMA_signal_4370) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_4375), .Q (new_AGEMA_signal_4376) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_4381), .Q (new_AGEMA_signal_4382) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_4387), .Q (new_AGEMA_signal_4388) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_4393), .Q (new_AGEMA_signal_4394) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_4399), .Q (new_AGEMA_signal_4400) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_4405), .Q (new_AGEMA_signal_4406) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_4411), .Q (new_AGEMA_signal_4412) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_4417), .Q (new_AGEMA_signal_4418) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_4423), .Q (new_AGEMA_signal_4424) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_4429), .Q (new_AGEMA_signal_4430) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_4435), .Q (new_AGEMA_signal_4436) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_4441), .Q (new_AGEMA_signal_4442) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_4447), .Q (new_AGEMA_signal_4448) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_4453), .Q (new_AGEMA_signal_4454) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_4459), .Q (new_AGEMA_signal_4460) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_4465), .Q (new_AGEMA_signal_4466) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_4471), .Q (new_AGEMA_signal_4472) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_4477), .Q (new_AGEMA_signal_4478) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_4483), .Q (new_AGEMA_signal_4484) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_4489), .Q (new_AGEMA_signal_4490) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_4495), .Q (new_AGEMA_signal_4496) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_4501), .Q (new_AGEMA_signal_4502) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_4507), .Q (new_AGEMA_signal_4508) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C (clk), .D (new_AGEMA_signal_4705), .Q (new_AGEMA_signal_4706) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_4712) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_4720) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_4728) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (new_AGEMA_signal_4736) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_4744) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_4752) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_4760) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_4768) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_4776) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_4784) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_4792) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_4800) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (new_AGEMA_signal_4808) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_4816) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_4824) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (new_AGEMA_signal_4832) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (new_AGEMA_signal_4840) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (new_AGEMA_signal_4848) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_4855), .Q (new_AGEMA_signal_4856) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (new_AGEMA_signal_4864) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (new_AGEMA_signal_4872) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (new_AGEMA_signal_4880) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_4888) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_4896) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_4904) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (new_AGEMA_signal_4912) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (new_AGEMA_signal_4920) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_4927), .Q (new_AGEMA_signal_4928) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_4936) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_4943), .Q (new_AGEMA_signal_4944) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_4951), .Q (new_AGEMA_signal_4952) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_4960) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_4967), .Q (new_AGEMA_signal_4968) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_4976) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_4984) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_4991), .Q (new_AGEMA_signal_4992) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_4999), .Q (new_AGEMA_signal_5000) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_5007), .Q (new_AGEMA_signal_5008) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_5015), .Q (new_AGEMA_signal_5016) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_5023), .Q (new_AGEMA_signal_5024) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_5032) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_5039), .Q (new_AGEMA_signal_5040) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_5047), .Q (new_AGEMA_signal_5048) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_5056) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_5063), .Q (new_AGEMA_signal_5064) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_5071), .Q (new_AGEMA_signal_5072) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_5079), .Q (new_AGEMA_signal_5080) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_5087), .Q (new_AGEMA_signal_5088) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_5095), .Q (new_AGEMA_signal_5096) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_5104) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_5111), .Q (new_AGEMA_signal_5112) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_5119), .Q (new_AGEMA_signal_5120) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_5127), .Q (new_AGEMA_signal_5128) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_5135), .Q (new_AGEMA_signal_5136) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_5144) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_5152) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_5159), .Q (new_AGEMA_signal_5160) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_5167), .Q (new_AGEMA_signal_5168) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_5176) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_5183), .Q (new_AGEMA_signal_5184) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_5192) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_5200) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_5207), .Q (new_AGEMA_signal_5208) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_5215), .Q (new_AGEMA_signal_5216) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_5224) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_5231), .Q (new_AGEMA_signal_5232) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_5239), .Q (new_AGEMA_signal_5240) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_5248) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_5255), .Q (new_AGEMA_signal_5256) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_5264) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_5272) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_5279), .Q (new_AGEMA_signal_5280) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_5287), .Q (new_AGEMA_signal_5288) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_5296) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_5303), .Q (new_AGEMA_signal_5304) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_5312) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_5320) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_5327), .Q (new_AGEMA_signal_5328) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_5336) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_5344) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_5351), .Q (new_AGEMA_signal_5352) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_5360) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_5367), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_5375), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_5384) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_5400) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_5408) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_5424) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_5431), .Q (new_AGEMA_signal_5432) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_5447), .Q (new_AGEMA_signal_5448) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_5456) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_5464) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_5471), .Q (new_AGEMA_signal_5472) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_5480) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_5487), .Q (new_AGEMA_signal_5488) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_5495), .Q (new_AGEMA_signal_5496) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_5504) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (new_AGEMA_signal_5512) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_5520) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_5528) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_5536) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_5544) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_5552) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_5560) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_5567), .Q (new_AGEMA_signal_5568) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (new_AGEMA_signal_5576) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_5584) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_5591), .Q (new_AGEMA_signal_5592) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_5600) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_5608) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_5615), .Q (new_AGEMA_signal_5616) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_5624) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_5631), .Q (new_AGEMA_signal_5632) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_5639), .Q (new_AGEMA_signal_5640) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_5647), .Q (new_AGEMA_signal_5648) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_5655), .Q (new_AGEMA_signal_5656) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_5663), .Q (new_AGEMA_signal_5664) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_5672) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_5680) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_5687), .Q (new_AGEMA_signal_5688) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_5696) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_5704) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_5711), .Q (new_AGEMA_signal_5712) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_5720) ) ;
    buf_clk new_AGEMA_reg_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_5728) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C (clk), .D (new_AGEMA_signal_5737), .Q (new_AGEMA_signal_5738) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C (clk), .D (new_AGEMA_signal_5745), .Q (new_AGEMA_signal_5746) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C (clk), .D (new_AGEMA_signal_5753), .Q (new_AGEMA_signal_5754) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C (clk), .D (new_AGEMA_signal_5761), .Q (new_AGEMA_signal_5762) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C (clk), .D (new_AGEMA_signal_5769), .Q (new_AGEMA_signal_5770) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C (clk), .D (new_AGEMA_signal_5777), .Q (new_AGEMA_signal_5778) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C (clk), .D (new_AGEMA_signal_5785), .Q (new_AGEMA_signal_5786) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C (clk), .D (new_AGEMA_signal_5793), .Q (new_AGEMA_signal_5794) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C (clk), .D (new_AGEMA_signal_5801), .Q (new_AGEMA_signal_5802) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C (clk), .D (new_AGEMA_signal_5809), .Q (new_AGEMA_signal_5810) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C (clk), .D (new_AGEMA_signal_5817), .Q (new_AGEMA_signal_5818) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C (clk), .D (new_AGEMA_signal_5825), .Q (new_AGEMA_signal_5826) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C (clk), .D (new_AGEMA_signal_5833), .Q (new_AGEMA_signal_5834) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C (clk), .D (new_AGEMA_signal_5841), .Q (new_AGEMA_signal_5842) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C (clk), .D (new_AGEMA_signal_5849), .Q (new_AGEMA_signal_5850) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C (clk), .D (new_AGEMA_signal_5857), .Q (new_AGEMA_signal_5858) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C (clk), .D (new_AGEMA_signal_5865), .Q (new_AGEMA_signal_5866) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C (clk), .D (new_AGEMA_signal_5873), .Q (new_AGEMA_signal_5874) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C (clk), .D (new_AGEMA_signal_5881), .Q (new_AGEMA_signal_5882) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C (clk), .D (new_AGEMA_signal_5889), .Q (new_AGEMA_signal_5890) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C (clk), .D (new_AGEMA_signal_5897), .Q (new_AGEMA_signal_5898) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C (clk), .D (new_AGEMA_signal_5905), .Q (new_AGEMA_signal_5906) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C (clk), .D (new_AGEMA_signal_5913), .Q (new_AGEMA_signal_5914) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C (clk), .D (new_AGEMA_signal_5921), .Q (new_AGEMA_signal_5922) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C (clk), .D (new_AGEMA_signal_5929), .Q (new_AGEMA_signal_5930) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C (clk), .D (new_AGEMA_signal_5937), .Q (new_AGEMA_signal_5938) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C (clk), .D (new_AGEMA_signal_5945), .Q (new_AGEMA_signal_5946) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C (clk), .D (new_AGEMA_signal_5953), .Q (new_AGEMA_signal_5954) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C (clk), .D (new_AGEMA_signal_5961), .Q (new_AGEMA_signal_5962) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C (clk), .D (new_AGEMA_signal_5969), .Q (new_AGEMA_signal_5970) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C (clk), .D (new_AGEMA_signal_5977), .Q (new_AGEMA_signal_5978) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C (clk), .D (new_AGEMA_signal_5985), .Q (new_AGEMA_signal_5986) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C (clk), .D (new_AGEMA_signal_5993), .Q (new_AGEMA_signal_5994) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C (clk), .D (new_AGEMA_signal_6001), .Q (new_AGEMA_signal_6002) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C (clk), .D (new_AGEMA_signal_6009), .Q (new_AGEMA_signal_6010) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C (clk), .D (new_AGEMA_signal_6017), .Q (new_AGEMA_signal_6018) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C (clk), .D (new_AGEMA_signal_6025), .Q (new_AGEMA_signal_6026) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C (clk), .D (new_AGEMA_signal_6033), .Q (new_AGEMA_signal_6034) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C (clk), .D (new_AGEMA_signal_6041), .Q (new_AGEMA_signal_6042) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C (clk), .D (new_AGEMA_signal_6049), .Q (new_AGEMA_signal_6050) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C (clk), .D (new_AGEMA_signal_6057), .Q (new_AGEMA_signal_6058) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C (clk), .D (new_AGEMA_signal_6065), .Q (new_AGEMA_signal_6066) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C (clk), .D (new_AGEMA_signal_6073), .Q (new_AGEMA_signal_6074) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C (clk), .D (new_AGEMA_signal_6081), .Q (new_AGEMA_signal_6082) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C (clk), .D (new_AGEMA_signal_6089), .Q (new_AGEMA_signal_6090) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C (clk), .D (new_AGEMA_signal_6097), .Q (new_AGEMA_signal_6098) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C (clk), .D (new_AGEMA_signal_6105), .Q (new_AGEMA_signal_6106) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C (clk), .D (new_AGEMA_signal_6113), .Q (new_AGEMA_signal_6114) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C (clk), .D (new_AGEMA_signal_6121), .Q (new_AGEMA_signal_6122) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C (clk), .D (new_AGEMA_signal_6129), .Q (new_AGEMA_signal_6130) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C (clk), .D (new_AGEMA_signal_6137), .Q (new_AGEMA_signal_6138) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C (clk), .D (new_AGEMA_signal_6145), .Q (new_AGEMA_signal_6146) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C (clk), .D (new_AGEMA_signal_6153), .Q (new_AGEMA_signal_6154) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C (clk), .D (new_AGEMA_signal_6161), .Q (new_AGEMA_signal_6162) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C (clk), .D (new_AGEMA_signal_6169), .Q (new_AGEMA_signal_6170) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C (clk), .D (new_AGEMA_signal_6177), .Q (new_AGEMA_signal_6178) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C (clk), .D (new_AGEMA_signal_6185), .Q (new_AGEMA_signal_6186) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C (clk), .D (new_AGEMA_signal_6193), .Q (new_AGEMA_signal_6194) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C (clk), .D (new_AGEMA_signal_6201), .Q (new_AGEMA_signal_6202) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C (clk), .D (new_AGEMA_signal_6209), .Q (new_AGEMA_signal_6210) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C (clk), .D (new_AGEMA_signal_6217), .Q (new_AGEMA_signal_6218) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C (clk), .D (new_AGEMA_signal_6225), .Q (new_AGEMA_signal_6226) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C (clk), .D (new_AGEMA_signal_6233), .Q (new_AGEMA_signal_6234) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C (clk), .D (new_AGEMA_signal_6241), .Q (new_AGEMA_signal_6242) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C (clk), .D (new_AGEMA_signal_4511), .Q (new_AGEMA_signal_6246) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_4513), .Q (new_AGEMA_signal_6248) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_6252) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C (clk), .D (new_AGEMA_signal_4523), .Q (new_AGEMA_signal_6258) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_4525), .Q (new_AGEMA_signal_6260) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C (clk), .D (new_AGEMA_signal_4535), .Q (new_AGEMA_signal_6270) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_4537), .Q (new_AGEMA_signal_6272) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C (clk), .D (new_AGEMA_signal_4547), .Q (new_AGEMA_signal_6282) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_4549), .Q (new_AGEMA_signal_6284) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_6287), .Q (new_AGEMA_signal_6288) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C (clk), .D (new_AGEMA_signal_4559), .Q (new_AGEMA_signal_6294) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_4561), .Q (new_AGEMA_signal_6296) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_6299), .Q (new_AGEMA_signal_6300) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_6304) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C (clk), .D (new_AGEMA_signal_4571), .Q (new_AGEMA_signal_6306) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_4573), .Q (new_AGEMA_signal_6308) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_6312) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C (clk), .D (new_AGEMA_signal_4583), .Q (new_AGEMA_signal_6318) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_4585), .Q (new_AGEMA_signal_6320) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_6324) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C (clk), .D (new_AGEMA_signal_4595), .Q (new_AGEMA_signal_6330) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_4597), .Q (new_AGEMA_signal_6332) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_6336) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_6340) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C (clk), .D (new_AGEMA_signal_4607), .Q (new_AGEMA_signal_6342) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_4609), .Q (new_AGEMA_signal_6344) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_6347), .Q (new_AGEMA_signal_6348) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_6352) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C (clk), .D (new_AGEMA_signal_4619), .Q (new_AGEMA_signal_6354) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_4621), .Q (new_AGEMA_signal_6356) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_6360) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_6366) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_6368) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_6371), .Q (new_AGEMA_signal_6372) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_6376) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C (clk), .D (new_AGEMA_signal_4643), .Q (new_AGEMA_signal_6378) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_4645), .Q (new_AGEMA_signal_6380) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_6384) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_6388) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_4655), .Q (new_AGEMA_signal_6390) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_4657), .Q (new_AGEMA_signal_6392) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_6396) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C (clk), .D (new_AGEMA_signal_4667), .Q (new_AGEMA_signal_6402) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_4669), .Q (new_AGEMA_signal_6404) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_6408) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_6412) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_6414) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_4681), .Q (new_AGEMA_signal_6416) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_6419), .Q (new_AGEMA_signal_6420) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_6424) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_6426) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_4693), .Q (new_AGEMA_signal_6428) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_6432) ) ;
    buf_clk new_AGEMA_reg_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_6436) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_6443), .Q (new_AGEMA_signal_6444) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_6451), .Q (new_AGEMA_signal_6452) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_6460) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_6467), .Q (new_AGEMA_signal_6468) ) ;

    /* cells in depth 6 */
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U128 ( .a ({new_AGEMA_signal_3363, new_AGEMA_signal_3357}), .b ({new_AGEMA_signal_2154, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_3032, new_AGEMA_signal_3014}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U126 ( .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3369}), .b ({new_AGEMA_signal_2148, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_3034, new_AGEMA_signal_3016}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U124 ( .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3381}), .b ({new_AGEMA_signal_2204, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_3036, new_AGEMA_signal_2960}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U122 ( .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3393}), .b ({new_AGEMA_signal_2206, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_3038, new_AGEMA_signal_2962}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U120 ( .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3405}), .b ({new_AGEMA_signal_2150, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_3040, new_AGEMA_signal_3018}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U119 ( .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3417}), .b ({new_AGEMA_signal_2200, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_3042, new_AGEMA_signal_2964}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U117 ( .a ({new_AGEMA_signal_3435, new_AGEMA_signal_3429}), .b ({new_AGEMA_signal_2202, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_3044, new_AGEMA_signal_2966}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U115 ( .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3441}), .b ({new_AGEMA_signal_2196, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_3046, new_AGEMA_signal_2968}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U113 ( .a ({new_AGEMA_signal_3459, new_AGEMA_signal_3453}), .b ({new_AGEMA_signal_2198, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_3048, new_AGEMA_signal_2970}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U111 ( .a ({new_AGEMA_signal_3471, new_AGEMA_signal_3465}), .b ({new_AGEMA_signal_2192, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_3050, new_AGEMA_signal_2972}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U108 ( .a ({new_AGEMA_signal_3483, new_AGEMA_signal_3477}), .b ({new_AGEMA_signal_2194, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_3052, new_AGEMA_signal_2974}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U106 ( .a ({new_AGEMA_signal_3495, new_AGEMA_signal_3489}), .b ({new_AGEMA_signal_2188, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_3054, new_AGEMA_signal_2976}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U104 ( .a ({new_AGEMA_signal_3507, new_AGEMA_signal_3501}), .b ({new_AGEMA_signal_2190, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_3056, new_AGEMA_signal_2978}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U102 ( .a ({new_AGEMA_signal_3519, new_AGEMA_signal_3513}), .b ({new_AGEMA_signal_2184, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_3058, new_AGEMA_signal_2980}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U100 ( .a ({new_AGEMA_signal_3531, new_AGEMA_signal_3525}), .b ({new_AGEMA_signal_2186, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_3060, new_AGEMA_signal_2982}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U98 ( .a ({new_AGEMA_signal_3543, new_AGEMA_signal_3537}), .b ({new_AGEMA_signal_2144, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_3062, new_AGEMA_signal_3020}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U97 ( .a ({new_AGEMA_signal_3555, new_AGEMA_signal_3549}), .b ({new_AGEMA_signal_2180, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_3064, new_AGEMA_signal_2984}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U95 ( .a ({new_AGEMA_signal_3567, new_AGEMA_signal_3561}), .b ({new_AGEMA_signal_2182, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_3066, new_AGEMA_signal_2986}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U93 ( .a ({new_AGEMA_signal_3579, new_AGEMA_signal_3573}), .b ({new_AGEMA_signal_2176, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_3068, new_AGEMA_signal_2988}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U91 ( .a ({new_AGEMA_signal_3591, new_AGEMA_signal_3585}), .b ({new_AGEMA_signal_2178, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_3070, new_AGEMA_signal_2990}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U89 ( .a ({new_AGEMA_signal_3603, new_AGEMA_signal_3597}), .b ({new_AGEMA_signal_2172, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_3072, new_AGEMA_signal_2992}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U86 ( .a ({new_AGEMA_signal_3615, new_AGEMA_signal_3609}), .b ({new_AGEMA_signal_2174, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_3074, new_AGEMA_signal_2994}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U84 ( .a ({new_AGEMA_signal_3627, new_AGEMA_signal_3621}), .b ({new_AGEMA_signal_2168, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_3076, new_AGEMA_signal_2996}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U82 ( .a ({new_AGEMA_signal_3639, new_AGEMA_signal_3633}), .b ({new_AGEMA_signal_2170, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_3078, new_AGEMA_signal_2998}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U80 ( .a ({new_AGEMA_signal_3651, new_AGEMA_signal_3645}), .b ({new_AGEMA_signal_2164, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_3080, new_AGEMA_signal_3000}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U78 ( .a ({new_AGEMA_signal_3663, new_AGEMA_signal_3657}), .b ({new_AGEMA_signal_2166, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_3082, new_AGEMA_signal_3002}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U76 ( .a ({new_AGEMA_signal_3675, new_AGEMA_signal_3669}), .b ({new_AGEMA_signal_2146, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_3084, new_AGEMA_signal_3022}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U75 ( .a ({new_AGEMA_signal_3687, new_AGEMA_signal_3681}), .b ({new_AGEMA_signal_2160, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_3086, new_AGEMA_signal_3004}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U73 ( .a ({new_AGEMA_signal_3699, new_AGEMA_signal_3693}), .b ({new_AGEMA_signal_2162, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_3088, new_AGEMA_signal_3006}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U71 ( .a ({new_AGEMA_signal_3711, new_AGEMA_signal_3705}), .b ({new_AGEMA_signal_2156, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_3090, new_AGEMA_signal_3008}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U69 ( .a ({new_AGEMA_signal_3723, new_AGEMA_signal_3717}), .b ({new_AGEMA_signal_2158, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_3092, new_AGEMA_signal_3010}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U67 ( .a ({new_AGEMA_signal_3735, new_AGEMA_signal_3729}), .b ({new_AGEMA_signal_2152, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_3094, new_AGEMA_signal_3012}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U144 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3741}), .b ({new_AGEMA_signal_2154, Midori_rounds_SR_Result[9]}), .c ({new_AGEMA_signal_2272, Midori_rounds_sub_ResultXORkey[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U142 ( .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3753}), .b ({new_AGEMA_signal_2148, Midori_rounds_SR_Result[47]}), .c ({new_AGEMA_signal_2273, Midori_rounds_sub_ResultXORkey[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U140 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3765}), .b ({new_AGEMA_signal_2204, Midori_rounds_SR_Result[63]}), .c ({new_AGEMA_signal_2275, Midori_rounds_sub_ResultXORkey[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U138 ( .a ({new_AGEMA_signal_3783, new_AGEMA_signal_3777}), .b ({new_AGEMA_signal_2206, Midori_rounds_SR_Result[61]}), .c ({new_AGEMA_signal_2277, Midori_rounds_sub_ResultXORkey[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U136 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3789}), .b ({new_AGEMA_signal_2150, Midori_rounds_SR_Result[45]}), .c ({new_AGEMA_signal_2278, Midori_rounds_sub_ResultXORkey[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U135 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3801}), .b ({new_AGEMA_signal_2200, Midori_rounds_SR_Result[35]}), .c ({new_AGEMA_signal_2279, Midori_rounds_sub_ResultXORkey[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U133 ( .a ({new_AGEMA_signal_3819, new_AGEMA_signal_3813}), .b ({new_AGEMA_signal_2202, Midori_rounds_SR_Result[33]}), .c ({new_AGEMA_signal_2281, Midori_rounds_sub_ResultXORkey[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U131 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3825}), .b ({new_AGEMA_signal_2196, Midori_rounds_SR_Result[7]}), .c ({new_AGEMA_signal_2282, Midori_rounds_sub_ResultXORkey[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U129 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3837}), .b ({new_AGEMA_signal_2198, Midori_rounds_SR_Result[5]}), .c ({new_AGEMA_signal_2284, Midori_rounds_sub_ResultXORkey[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U127 ( .a ({new_AGEMA_signal_3855, new_AGEMA_signal_3849}), .b ({new_AGEMA_signal_2192, Midori_rounds_SR_Result[27]}), .c ({new_AGEMA_signal_2285, Midori_rounds_sub_ResultXORkey[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U124 ( .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3861}), .b ({new_AGEMA_signal_2194, Midori_rounds_SR_Result[25]}), .c ({new_AGEMA_signal_2287, Midori_rounds_sub_ResultXORkey[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U122 ( .a ({new_AGEMA_signal_3879, new_AGEMA_signal_3873}), .b ({new_AGEMA_signal_2188, Midori_rounds_SR_Result[43]}), .c ({new_AGEMA_signal_2288, Midori_rounds_sub_ResultXORkey[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U120 ( .a ({new_AGEMA_signal_3891, new_AGEMA_signal_3885}), .b ({new_AGEMA_signal_2190, Midori_rounds_SR_Result[41]}), .c ({new_AGEMA_signal_2290, Midori_rounds_sub_ResultXORkey[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U118 ( .a ({new_AGEMA_signal_3903, new_AGEMA_signal_3897}), .b ({new_AGEMA_signal_2184, Midori_rounds_SR_Result[55]}), .c ({new_AGEMA_signal_2291, Midori_rounds_sub_ResultXORkey[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U116 ( .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3909}), .b ({new_AGEMA_signal_2186, Midori_rounds_SR_Result[53]}), .c ({new_AGEMA_signal_2293, Midori_rounds_sub_ResultXORkey[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U114 ( .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3921}), .b ({new_AGEMA_signal_2144, Midori_rounds_SR_Result[51]}), .c ({new_AGEMA_signal_2294, Midori_rounds_sub_ResultXORkey[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U113 ( .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3933}), .b ({new_AGEMA_signal_2180, Midori_rounds_SR_Result[19]}), .c ({new_AGEMA_signal_2295, Midori_rounds_sub_ResultXORkey[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U111 ( .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3945}), .b ({new_AGEMA_signal_2182, Midori_rounds_SR_Result[17]}), .c ({new_AGEMA_signal_2297, Midori_rounds_sub_ResultXORkey[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U109 ( .a ({new_AGEMA_signal_3963, new_AGEMA_signal_3957}), .b ({new_AGEMA_signal_2176, Midori_rounds_SR_Result[15]}), .c ({new_AGEMA_signal_2298, Midori_rounds_sub_ResultXORkey[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U107 ( .a ({new_AGEMA_signal_3975, new_AGEMA_signal_3969}), .b ({new_AGEMA_signal_2178, Midori_rounds_SR_Result[13]}), .c ({new_AGEMA_signal_2300, Midori_rounds_sub_ResultXORkey[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U105 ( .a ({new_AGEMA_signal_3987, new_AGEMA_signal_3981}), .b ({new_AGEMA_signal_2172, Midori_rounds_SR_Result[3]}), .c ({new_AGEMA_signal_2301, Midori_rounds_sub_ResultXORkey[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U102 ( .a ({new_AGEMA_signal_3999, new_AGEMA_signal_3993}), .b ({new_AGEMA_signal_2174, Midori_rounds_SR_Result[1]}), .c ({new_AGEMA_signal_2304, Midori_rounds_sub_ResultXORkey[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U100 ( .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4005}), .b ({new_AGEMA_signal_2168, Midori_rounds_SR_Result[31]}), .c ({new_AGEMA_signal_2305, Midori_rounds_sub_ResultXORkey[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U98 ( .a ({new_AGEMA_signal_4023, new_AGEMA_signal_4017}), .b ({new_AGEMA_signal_2170, Midori_rounds_SR_Result[29]}), .c ({new_AGEMA_signal_2307, Midori_rounds_sub_ResultXORkey[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U96 ( .a ({new_AGEMA_signal_4035, new_AGEMA_signal_4029}), .b ({new_AGEMA_signal_2164, Midori_rounds_SR_Result[59]}), .c ({new_AGEMA_signal_2308, Midori_rounds_sub_ResultXORkey[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U94 ( .a ({new_AGEMA_signal_4047, new_AGEMA_signal_4041}), .b ({new_AGEMA_signal_2166, Midori_rounds_SR_Result[57]}), .c ({new_AGEMA_signal_2310, Midori_rounds_sub_ResultXORkey[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U92 ( .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4053}), .b ({new_AGEMA_signal_2146, Midori_rounds_SR_Result[49]}), .c ({new_AGEMA_signal_2311, Midori_rounds_sub_ResultXORkey[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U91 ( .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4065}), .b ({new_AGEMA_signal_2160, Midori_rounds_SR_Result[39]}), .c ({new_AGEMA_signal_2312, Midori_rounds_sub_ResultXORkey[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U89 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4077}), .b ({new_AGEMA_signal_2162, Midori_rounds_SR_Result[37]}), .c ({new_AGEMA_signal_2314, Midori_rounds_sub_ResultXORkey[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U87 ( .a ({new_AGEMA_signal_4095, new_AGEMA_signal_4089}), .b ({new_AGEMA_signal_2156, Midori_rounds_SR_Result[23]}), .c ({new_AGEMA_signal_2315, Midori_rounds_sub_ResultXORkey[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U85 ( .a ({new_AGEMA_signal_4107, new_AGEMA_signal_4101}), .b ({new_AGEMA_signal_2158, Midori_rounds_SR_Result[21]}), .c ({new_AGEMA_signal_2317, Midori_rounds_sub_ResultXORkey[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U83 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4113}), .b ({new_AGEMA_signal_2152, Midori_rounds_SR_Result[11]}), .c ({new_AGEMA_signal_2318, Midori_rounds_sub_ResultXORkey[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U80 ( .a ({new_AGEMA_signal_3747, new_AGEMA_signal_3741}), .b ({new_AGEMA_signal_2428, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_2440, Midori_rounds_mul_ResultXORkey[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U77 ( .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3753}), .b ({new_AGEMA_signal_2429, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_2442, Midori_rounds_mul_ResultXORkey[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U75 ( .a ({new_AGEMA_signal_3771, new_AGEMA_signal_3765}), .b ({new_AGEMA_signal_2399, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_2444, Midori_rounds_mul_ResultXORkey[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U73 ( .a ({new_AGEMA_signal_3783, new_AGEMA_signal_3777}), .b ({new_AGEMA_signal_2401, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_2446, Midori_rounds_mul_ResultXORkey[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U70 ( .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3789}), .b ({new_AGEMA_signal_2431, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_2447, Midori_rounds_mul_ResultXORkey[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U69 ( .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3801}), .b ({new_AGEMA_signal_2402, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_2448, Midori_rounds_mul_ResultXORkey[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U67 ( .a ({new_AGEMA_signal_3819, new_AGEMA_signal_3813}), .b ({new_AGEMA_signal_2392, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_2450, Midori_rounds_mul_ResultXORkey[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U64 ( .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3825}), .b ({new_AGEMA_signal_2393, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_2451, Midori_rounds_mul_ResultXORkey[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U62 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3837}), .b ({new_AGEMA_signal_2395, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_2453, Midori_rounds_mul_ResultXORkey[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U59 ( .a ({new_AGEMA_signal_3855, new_AGEMA_signal_3849}), .b ({new_AGEMA_signal_2396, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_2454, Midori_rounds_mul_ResultXORkey[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U55 ( .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3861}), .b ({new_AGEMA_signal_2398, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_2456, Midori_rounds_mul_ResultXORkey[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U52 ( .a ({new_AGEMA_signal_3879, new_AGEMA_signal_3873}), .b ({new_AGEMA_signal_2411, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_2457, Midori_rounds_mul_ResultXORkey[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U50 ( .a ({new_AGEMA_signal_3891, new_AGEMA_signal_3885}), .b ({new_AGEMA_signal_2413, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_2459, Midori_rounds_mul_ResultXORkey[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U47 ( .a ({new_AGEMA_signal_3903, new_AGEMA_signal_3897}), .b ({new_AGEMA_signal_2414, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_2461, Midori_rounds_mul_ResultXORkey[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U45 ( .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3909}), .b ({new_AGEMA_signal_2404, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_2463, Midori_rounds_mul_ResultXORkey[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U42 ( .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3921}), .b ({new_AGEMA_signal_2432, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_2464, Midori_rounds_mul_ResultXORkey[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U41 ( .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3933}), .b ({new_AGEMA_signal_2405, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_2465, Midori_rounds_mul_ResultXORkey[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U39 ( .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3945}), .b ({new_AGEMA_signal_2407, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_2467, Midori_rounds_mul_ResultXORkey[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U36 ( .a ({new_AGEMA_signal_3963, new_AGEMA_signal_3957}), .b ({new_AGEMA_signal_2408, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_2469, Midori_rounds_mul_ResultXORkey[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U34 ( .a ({new_AGEMA_signal_3975, new_AGEMA_signal_3969}), .b ({new_AGEMA_signal_2410, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_2471, Midori_rounds_mul_ResultXORkey[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U31 ( .a ({new_AGEMA_signal_3987, new_AGEMA_signal_3981}), .b ({new_AGEMA_signal_2423, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_2472, Midori_rounds_mul_ResultXORkey[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U28 ( .a ({new_AGEMA_signal_3999, new_AGEMA_signal_3993}), .b ({new_AGEMA_signal_2425, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_2475, Midori_rounds_mul_ResultXORkey[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U25 ( .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4005}), .b ({new_AGEMA_signal_2426, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_2476, Midori_rounds_mul_ResultXORkey[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U23 ( .a ({new_AGEMA_signal_4023, new_AGEMA_signal_4017}), .b ({new_AGEMA_signal_2416, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_2478, Midori_rounds_mul_ResultXORkey[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U20 ( .a ({new_AGEMA_signal_4035, new_AGEMA_signal_4029}), .b ({new_AGEMA_signal_2417, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_2479, Midori_rounds_mul_ResultXORkey[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U18 ( .a ({new_AGEMA_signal_4047, new_AGEMA_signal_4041}), .b ({new_AGEMA_signal_2419, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_2481, Midori_rounds_mul_ResultXORkey[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U15 ( .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4053}), .b ({new_AGEMA_signal_2434, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_2483, Midori_rounds_mul_ResultXORkey[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U14 ( .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4065}), .b ({new_AGEMA_signal_2420, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_2484, Midori_rounds_mul_ResultXORkey[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U12 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4077}), .b ({new_AGEMA_signal_2422, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_2486, Midori_rounds_mul_ResultXORkey[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U9 ( .a ({new_AGEMA_signal_4095, new_AGEMA_signal_4089}), .b ({new_AGEMA_signal_2435, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_2487, Midori_rounds_mul_ResultXORkey[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U7 ( .a ({new_AGEMA_signal_4107, new_AGEMA_signal_4101}), .b ({new_AGEMA_signal_2437, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_2489, Midori_rounds_mul_ResultXORkey[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U4 ( .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4113}), .b ({new_AGEMA_signal_2438, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_2490, Midori_rounds_mul_ResultXORkey[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2506, Midori_rounds_round_Result[1]}), .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4131}), .c ({new_AGEMA_signal_2565, Midori_rounds_roundResult_Reg_SFF_1_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2508, Midori_rounds_round_Result[3]}), .a ({new_AGEMA_signal_4149, new_AGEMA_signal_4143}), .c ({new_AGEMA_signal_2567, Midori_rounds_roundResult_Reg_SFF_3_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2509, Midori_rounds_round_Result[5]}), .a ({new_AGEMA_signal_4161, new_AGEMA_signal_4155}), .c ({new_AGEMA_signal_2568, Midori_rounds_roundResult_Reg_SFF_5_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2511, Midori_rounds_round_Result[7]}), .a ({new_AGEMA_signal_4173, new_AGEMA_signal_4167}), .c ({new_AGEMA_signal_2570, Midori_rounds_roundResult_Reg_SFF_7_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2512, Midori_rounds_round_Result[9]}), .a ({new_AGEMA_signal_4185, new_AGEMA_signal_4179}), .c ({new_AGEMA_signal_2571, Midori_rounds_roundResult_Reg_SFF_9_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2514, Midori_rounds_round_Result[11]}), .a ({new_AGEMA_signal_4197, new_AGEMA_signal_4191}), .c ({new_AGEMA_signal_2573, Midori_rounds_roundResult_Reg_SFF_11_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2515, Midori_rounds_round_Result[13]}), .a ({new_AGEMA_signal_4209, new_AGEMA_signal_4203}), .c ({new_AGEMA_signal_2574, Midori_rounds_roundResult_Reg_SFF_13_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2517, Midori_rounds_round_Result[15]}), .a ({new_AGEMA_signal_4221, new_AGEMA_signal_4215}), .c ({new_AGEMA_signal_2576, Midori_rounds_roundResult_Reg_SFF_15_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2518, Midori_rounds_round_Result[17]}), .a ({new_AGEMA_signal_4233, new_AGEMA_signal_4227}), .c ({new_AGEMA_signal_2577, Midori_rounds_roundResult_Reg_SFF_17_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2520, Midori_rounds_round_Result[19]}), .a ({new_AGEMA_signal_4245, new_AGEMA_signal_4239}), .c ({new_AGEMA_signal_2579, Midori_rounds_roundResult_Reg_SFF_19_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2521, Midori_rounds_round_Result[21]}), .a ({new_AGEMA_signal_4257, new_AGEMA_signal_4251}), .c ({new_AGEMA_signal_2580, Midori_rounds_roundResult_Reg_SFF_21_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2523, Midori_rounds_round_Result[23]}), .a ({new_AGEMA_signal_4269, new_AGEMA_signal_4263}), .c ({new_AGEMA_signal_2582, Midori_rounds_roundResult_Reg_SFF_23_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2524, Midori_rounds_round_Result[25]}), .a ({new_AGEMA_signal_4281, new_AGEMA_signal_4275}), .c ({new_AGEMA_signal_2583, Midori_rounds_roundResult_Reg_SFF_25_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2526, Midori_rounds_round_Result[27]}), .a ({new_AGEMA_signal_4293, new_AGEMA_signal_4287}), .c ({new_AGEMA_signal_2585, Midori_rounds_roundResult_Reg_SFF_27_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2527, Midori_rounds_round_Result[29]}), .a ({new_AGEMA_signal_4305, new_AGEMA_signal_4299}), .c ({new_AGEMA_signal_2586, Midori_rounds_roundResult_Reg_SFF_29_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2529, Midori_rounds_round_Result[31]}), .a ({new_AGEMA_signal_4317, new_AGEMA_signal_4311}), .c ({new_AGEMA_signal_2588, Midori_rounds_roundResult_Reg_SFF_31_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2530, Midori_rounds_round_Result[33]}), .a ({new_AGEMA_signal_4329, new_AGEMA_signal_4323}), .c ({new_AGEMA_signal_2589, Midori_rounds_roundResult_Reg_SFF_33_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2532, Midori_rounds_round_Result[35]}), .a ({new_AGEMA_signal_4341, new_AGEMA_signal_4335}), .c ({new_AGEMA_signal_2591, Midori_rounds_roundResult_Reg_SFF_35_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2533, Midori_rounds_round_Result[37]}), .a ({new_AGEMA_signal_4353, new_AGEMA_signal_4347}), .c ({new_AGEMA_signal_2592, Midori_rounds_roundResult_Reg_SFF_37_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2535, Midori_rounds_round_Result[39]}), .a ({new_AGEMA_signal_4365, new_AGEMA_signal_4359}), .c ({new_AGEMA_signal_2594, Midori_rounds_roundResult_Reg_SFF_39_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2536, Midori_rounds_round_Result[41]}), .a ({new_AGEMA_signal_4377, new_AGEMA_signal_4371}), .c ({new_AGEMA_signal_2595, Midori_rounds_roundResult_Reg_SFF_41_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2538, Midori_rounds_round_Result[43]}), .a ({new_AGEMA_signal_4389, new_AGEMA_signal_4383}), .c ({new_AGEMA_signal_2597, Midori_rounds_roundResult_Reg_SFF_43_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2539, Midori_rounds_round_Result[45]}), .a ({new_AGEMA_signal_4401, new_AGEMA_signal_4395}), .c ({new_AGEMA_signal_2598, Midori_rounds_roundResult_Reg_SFF_45_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2541, Midori_rounds_round_Result[47]}), .a ({new_AGEMA_signal_4413, new_AGEMA_signal_4407}), .c ({new_AGEMA_signal_2600, Midori_rounds_roundResult_Reg_SFF_47_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2542, Midori_rounds_round_Result[49]}), .a ({new_AGEMA_signal_4425, new_AGEMA_signal_4419}), .c ({new_AGEMA_signal_2601, Midori_rounds_roundResult_Reg_SFF_49_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2544, Midori_rounds_round_Result[51]}), .a ({new_AGEMA_signal_4437, new_AGEMA_signal_4431}), .c ({new_AGEMA_signal_2603, Midori_rounds_roundResult_Reg_SFF_51_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2545, Midori_rounds_round_Result[53]}), .a ({new_AGEMA_signal_4449, new_AGEMA_signal_4443}), .c ({new_AGEMA_signal_2604, Midori_rounds_roundResult_Reg_SFF_53_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2547, Midori_rounds_round_Result[55]}), .a ({new_AGEMA_signal_4461, new_AGEMA_signal_4455}), .c ({new_AGEMA_signal_2606, Midori_rounds_roundResult_Reg_SFF_55_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2548, Midori_rounds_round_Result[57]}), .a ({new_AGEMA_signal_4473, new_AGEMA_signal_4467}), .c ({new_AGEMA_signal_2607, Midori_rounds_roundResult_Reg_SFF_57_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2550, Midori_rounds_round_Result[59]}), .a ({new_AGEMA_signal_4485, new_AGEMA_signal_4479}), .c ({new_AGEMA_signal_2609, Midori_rounds_roundResult_Reg_SFF_59_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2551, Midori_rounds_round_Result[61]}), .a ({new_AGEMA_signal_4497, new_AGEMA_signal_4491}), .c ({new_AGEMA_signal_2610, Midori_rounds_roundResult_Reg_SFF_61_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1 ( .s (new_AGEMA_signal_4125), .b ({new_AGEMA_signal_2553, Midori_rounds_round_Result[63]}), .a ({new_AGEMA_signal_4509, new_AGEMA_signal_4503}), .c ({new_AGEMA_signal_2612, Midori_rounds_roundResult_Reg_SFF_63_DQ}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .a ({new_AGEMA_signal_4513, new_AGEMA_signal_4511}), .b ({new_AGEMA_signal_2065, Midori_rounds_sub_sBox_PRINCE_0_n14}), .clk (clk), .r (Fresh[160]), .c ({new_AGEMA_signal_2144, Midori_rounds_SR_Result[51]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .a ({new_AGEMA_signal_1917, Midori_rounds_sub_sBox_PRINCE_0_n11}), .b ({new_AGEMA_signal_4517, new_AGEMA_signal_4515}), .clk (clk), .r (Fresh[161]), .c ({new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_0_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .a ({new_AGEMA_signal_4521, new_AGEMA_signal_4519}), .b ({new_AGEMA_signal_2067, Midori_rounds_sub_sBox_PRINCE_0_n5}), .clk (clk), .r (Fresh[162]), .c ({new_AGEMA_signal_2146, Midori_rounds_SR_Result[49]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .a ({new_AGEMA_signal_4517, new_AGEMA_signal_4515}), .b ({new_AGEMA_signal_1921, Midori_rounds_sub_sBox_PRINCE_0_n2}), .clk (clk), .r (Fresh[163]), .c ({new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_0_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .a ({new_AGEMA_signal_4525, new_AGEMA_signal_4523}), .b ({new_AGEMA_signal_2070, Midori_rounds_sub_sBox_PRINCE_1_n14}), .clk (clk), .r (Fresh[164]), .c ({new_AGEMA_signal_2148, Midori_rounds_SR_Result[47]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .a ({new_AGEMA_signal_1923, Midori_rounds_sub_sBox_PRINCE_1_n11}), .b ({new_AGEMA_signal_4529, new_AGEMA_signal_4527}), .clk (clk), .r (Fresh[165]), .c ({new_AGEMA_signal_2071, Midori_rounds_sub_sBox_PRINCE_1_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .a ({new_AGEMA_signal_4533, new_AGEMA_signal_4531}), .b ({new_AGEMA_signal_2072, Midori_rounds_sub_sBox_PRINCE_1_n5}), .clk (clk), .r (Fresh[166]), .c ({new_AGEMA_signal_2150, Midori_rounds_SR_Result[45]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .a ({new_AGEMA_signal_4529, new_AGEMA_signal_4527}), .b ({new_AGEMA_signal_1927, Midori_rounds_sub_sBox_PRINCE_1_n2}), .clk (clk), .r (Fresh[167]), .c ({new_AGEMA_signal_2073, Midori_rounds_sub_sBox_PRINCE_1_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .a ({new_AGEMA_signal_4537, new_AGEMA_signal_4535}), .b ({new_AGEMA_signal_2075, Midori_rounds_sub_sBox_PRINCE_2_n14}), .clk (clk), .r (Fresh[168]), .c ({new_AGEMA_signal_2152, Midori_rounds_SR_Result[11]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .a ({new_AGEMA_signal_1929, Midori_rounds_sub_sBox_PRINCE_2_n11}), .b ({new_AGEMA_signal_4541, new_AGEMA_signal_4539}), .clk (clk), .r (Fresh[169]), .c ({new_AGEMA_signal_2076, Midori_rounds_sub_sBox_PRINCE_2_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .a ({new_AGEMA_signal_4545, new_AGEMA_signal_4543}), .b ({new_AGEMA_signal_2077, Midori_rounds_sub_sBox_PRINCE_2_n5}), .clk (clk), .r (Fresh[170]), .c ({new_AGEMA_signal_2154, Midori_rounds_SR_Result[9]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .a ({new_AGEMA_signal_4541, new_AGEMA_signal_4539}), .b ({new_AGEMA_signal_1933, Midori_rounds_sub_sBox_PRINCE_2_n2}), .clk (clk), .r (Fresh[171]), .c ({new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_2_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .a ({new_AGEMA_signal_4549, new_AGEMA_signal_4547}), .b ({new_AGEMA_signal_2080, Midori_rounds_sub_sBox_PRINCE_3_n14}), .clk (clk), .r (Fresh[172]), .c ({new_AGEMA_signal_2156, Midori_rounds_SR_Result[23]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .a ({new_AGEMA_signal_1935, Midori_rounds_sub_sBox_PRINCE_3_n11}), .b ({new_AGEMA_signal_4553, new_AGEMA_signal_4551}), .clk (clk), .r (Fresh[173]), .c ({new_AGEMA_signal_2081, Midori_rounds_sub_sBox_PRINCE_3_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .a ({new_AGEMA_signal_4557, new_AGEMA_signal_4555}), .b ({new_AGEMA_signal_2082, Midori_rounds_sub_sBox_PRINCE_3_n5}), .clk (clk), .r (Fresh[174]), .c ({new_AGEMA_signal_2158, Midori_rounds_SR_Result[21]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .a ({new_AGEMA_signal_4553, new_AGEMA_signal_4551}), .b ({new_AGEMA_signal_1939, Midori_rounds_sub_sBox_PRINCE_3_n2}), .clk (clk), .r (Fresh[175]), .c ({new_AGEMA_signal_2083, Midori_rounds_sub_sBox_PRINCE_3_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .a ({new_AGEMA_signal_4561, new_AGEMA_signal_4559}), .b ({new_AGEMA_signal_2085, Midori_rounds_sub_sBox_PRINCE_4_n14}), .clk (clk), .r (Fresh[176]), .c ({new_AGEMA_signal_2160, Midori_rounds_SR_Result[39]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .a ({new_AGEMA_signal_1941, Midori_rounds_sub_sBox_PRINCE_4_n11}), .b ({new_AGEMA_signal_4565, new_AGEMA_signal_4563}), .clk (clk), .r (Fresh[177]), .c ({new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_4_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .a ({new_AGEMA_signal_4569, new_AGEMA_signal_4567}), .b ({new_AGEMA_signal_2087, Midori_rounds_sub_sBox_PRINCE_4_n5}), .clk (clk), .r (Fresh[178]), .c ({new_AGEMA_signal_2162, Midori_rounds_SR_Result[37]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .a ({new_AGEMA_signal_4565, new_AGEMA_signal_4563}), .b ({new_AGEMA_signal_1945, Midori_rounds_sub_sBox_PRINCE_4_n2}), .clk (clk), .r (Fresh[179]), .c ({new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_4_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .a ({new_AGEMA_signal_4573, new_AGEMA_signal_4571}), .b ({new_AGEMA_signal_2090, Midori_rounds_sub_sBox_PRINCE_5_n14}), .clk (clk), .r (Fresh[180]), .c ({new_AGEMA_signal_2164, Midori_rounds_SR_Result[59]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .a ({new_AGEMA_signal_1947, Midori_rounds_sub_sBox_PRINCE_5_n11}), .b ({new_AGEMA_signal_4577, new_AGEMA_signal_4575}), .clk (clk), .r (Fresh[181]), .c ({new_AGEMA_signal_2091, Midori_rounds_sub_sBox_PRINCE_5_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .a ({new_AGEMA_signal_4581, new_AGEMA_signal_4579}), .b ({new_AGEMA_signal_2092, Midori_rounds_sub_sBox_PRINCE_5_n5}), .clk (clk), .r (Fresh[182]), .c ({new_AGEMA_signal_2166, Midori_rounds_SR_Result[57]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .a ({new_AGEMA_signal_4577, new_AGEMA_signal_4575}), .b ({new_AGEMA_signal_1951, Midori_rounds_sub_sBox_PRINCE_5_n2}), .clk (clk), .r (Fresh[183]), .c ({new_AGEMA_signal_2093, Midori_rounds_sub_sBox_PRINCE_5_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .a ({new_AGEMA_signal_4585, new_AGEMA_signal_4583}), .b ({new_AGEMA_signal_2095, Midori_rounds_sub_sBox_PRINCE_6_n14}), .clk (clk), .r (Fresh[184]), .c ({new_AGEMA_signal_2168, Midori_rounds_SR_Result[31]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .a ({new_AGEMA_signal_1953, Midori_rounds_sub_sBox_PRINCE_6_n11}), .b ({new_AGEMA_signal_4589, new_AGEMA_signal_4587}), .clk (clk), .r (Fresh[185]), .c ({new_AGEMA_signal_2096, Midori_rounds_sub_sBox_PRINCE_6_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4591}), .b ({new_AGEMA_signal_2097, Midori_rounds_sub_sBox_PRINCE_6_n5}), .clk (clk), .r (Fresh[186]), .c ({new_AGEMA_signal_2170, Midori_rounds_SR_Result[29]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .a ({new_AGEMA_signal_4589, new_AGEMA_signal_4587}), .b ({new_AGEMA_signal_1957, Midori_rounds_sub_sBox_PRINCE_6_n2}), .clk (clk), .r (Fresh[187]), .c ({new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_6_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .a ({new_AGEMA_signal_4597, new_AGEMA_signal_4595}), .b ({new_AGEMA_signal_2100, Midori_rounds_sub_sBox_PRINCE_7_n14}), .clk (clk), .r (Fresh[188]), .c ({new_AGEMA_signal_2172, Midori_rounds_SR_Result[3]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .a ({new_AGEMA_signal_1959, Midori_rounds_sub_sBox_PRINCE_7_n11}), .b ({new_AGEMA_signal_4601, new_AGEMA_signal_4599}), .clk (clk), .r (Fresh[189]), .c ({new_AGEMA_signal_2101, Midori_rounds_sub_sBox_PRINCE_7_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .a ({new_AGEMA_signal_4605, new_AGEMA_signal_4603}), .b ({new_AGEMA_signal_2102, Midori_rounds_sub_sBox_PRINCE_7_n5}), .clk (clk), .r (Fresh[190]), .c ({new_AGEMA_signal_2174, Midori_rounds_SR_Result[1]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .a ({new_AGEMA_signal_4601, new_AGEMA_signal_4599}), .b ({new_AGEMA_signal_1963, Midori_rounds_sub_sBox_PRINCE_7_n2}), .clk (clk), .r (Fresh[191]), .c ({new_AGEMA_signal_2103, Midori_rounds_sub_sBox_PRINCE_7_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .a ({new_AGEMA_signal_4609, new_AGEMA_signal_4607}), .b ({new_AGEMA_signal_2105, Midori_rounds_sub_sBox_PRINCE_8_n14}), .clk (clk), .r (Fresh[192]), .c ({new_AGEMA_signal_2176, Midori_rounds_SR_Result[15]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .a ({new_AGEMA_signal_1965, Midori_rounds_sub_sBox_PRINCE_8_n11}), .b ({new_AGEMA_signal_4613, new_AGEMA_signal_4611}), .clk (clk), .r (Fresh[193]), .c ({new_AGEMA_signal_2106, Midori_rounds_sub_sBox_PRINCE_8_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .a ({new_AGEMA_signal_4617, new_AGEMA_signal_4615}), .b ({new_AGEMA_signal_2107, Midori_rounds_sub_sBox_PRINCE_8_n5}), .clk (clk), .r (Fresh[194]), .c ({new_AGEMA_signal_2178, Midori_rounds_SR_Result[13]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .a ({new_AGEMA_signal_4613, new_AGEMA_signal_4611}), .b ({new_AGEMA_signal_1969, Midori_rounds_sub_sBox_PRINCE_8_n2}), .clk (clk), .r (Fresh[195]), .c ({new_AGEMA_signal_2108, Midori_rounds_sub_sBox_PRINCE_8_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .a ({new_AGEMA_signal_4621, new_AGEMA_signal_4619}), .b ({new_AGEMA_signal_2110, Midori_rounds_sub_sBox_PRINCE_9_n14}), .clk (clk), .r (Fresh[196]), .c ({new_AGEMA_signal_2180, Midori_rounds_SR_Result[19]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .a ({new_AGEMA_signal_1971, Midori_rounds_sub_sBox_PRINCE_9_n11}), .b ({new_AGEMA_signal_4625, new_AGEMA_signal_4623}), .clk (clk), .r (Fresh[197]), .c ({new_AGEMA_signal_2111, Midori_rounds_sub_sBox_PRINCE_9_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .a ({new_AGEMA_signal_4629, new_AGEMA_signal_4627}), .b ({new_AGEMA_signal_2112, Midori_rounds_sub_sBox_PRINCE_9_n5}), .clk (clk), .r (Fresh[198]), .c ({new_AGEMA_signal_2182, Midori_rounds_SR_Result[17]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .a ({new_AGEMA_signal_4625, new_AGEMA_signal_4623}), .b ({new_AGEMA_signal_1975, Midori_rounds_sub_sBox_PRINCE_9_n2}), .clk (clk), .r (Fresh[199]), .c ({new_AGEMA_signal_2113, Midori_rounds_sub_sBox_PRINCE_9_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .a ({new_AGEMA_signal_4633, new_AGEMA_signal_4631}), .b ({new_AGEMA_signal_2115, Midori_rounds_sub_sBox_PRINCE_10_n14}), .clk (clk), .r (Fresh[200]), .c ({new_AGEMA_signal_2184, Midori_rounds_SR_Result[55]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .a ({new_AGEMA_signal_1977, Midori_rounds_sub_sBox_PRINCE_10_n11}), .b ({new_AGEMA_signal_4637, new_AGEMA_signal_4635}), .clk (clk), .r (Fresh[201]), .c ({new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_10_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .a ({new_AGEMA_signal_4641, new_AGEMA_signal_4639}), .b ({new_AGEMA_signal_2117, Midori_rounds_sub_sBox_PRINCE_10_n5}), .clk (clk), .r (Fresh[202]), .c ({new_AGEMA_signal_2186, Midori_rounds_SR_Result[53]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .a ({new_AGEMA_signal_4637, new_AGEMA_signal_4635}), .b ({new_AGEMA_signal_1981, Midori_rounds_sub_sBox_PRINCE_10_n2}), .clk (clk), .r (Fresh[203]), .c ({new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_10_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .a ({new_AGEMA_signal_4645, new_AGEMA_signal_4643}), .b ({new_AGEMA_signal_2120, Midori_rounds_sub_sBox_PRINCE_11_n14}), .clk (clk), .r (Fresh[204]), .c ({new_AGEMA_signal_2188, Midori_rounds_SR_Result[43]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .a ({new_AGEMA_signal_1983, Midori_rounds_sub_sBox_PRINCE_11_n11}), .b ({new_AGEMA_signal_4649, new_AGEMA_signal_4647}), .clk (clk), .r (Fresh[205]), .c ({new_AGEMA_signal_2121, Midori_rounds_sub_sBox_PRINCE_11_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .a ({new_AGEMA_signal_4653, new_AGEMA_signal_4651}), .b ({new_AGEMA_signal_2122, Midori_rounds_sub_sBox_PRINCE_11_n5}), .clk (clk), .r (Fresh[206]), .c ({new_AGEMA_signal_2190, Midori_rounds_SR_Result[41]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .a ({new_AGEMA_signal_4649, new_AGEMA_signal_4647}), .b ({new_AGEMA_signal_1987, Midori_rounds_sub_sBox_PRINCE_11_n2}), .clk (clk), .r (Fresh[207]), .c ({new_AGEMA_signal_2123, Midori_rounds_sub_sBox_PRINCE_11_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .a ({new_AGEMA_signal_4657, new_AGEMA_signal_4655}), .b ({new_AGEMA_signal_2125, Midori_rounds_sub_sBox_PRINCE_12_n14}), .clk (clk), .r (Fresh[208]), .c ({new_AGEMA_signal_2192, Midori_rounds_SR_Result[27]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .a ({new_AGEMA_signal_1989, Midori_rounds_sub_sBox_PRINCE_12_n11}), .b ({new_AGEMA_signal_4661, new_AGEMA_signal_4659}), .clk (clk), .r (Fresh[209]), .c ({new_AGEMA_signal_2126, Midori_rounds_sub_sBox_PRINCE_12_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .a ({new_AGEMA_signal_4665, new_AGEMA_signal_4663}), .b ({new_AGEMA_signal_2127, Midori_rounds_sub_sBox_PRINCE_12_n5}), .clk (clk), .r (Fresh[210]), .c ({new_AGEMA_signal_2194, Midori_rounds_SR_Result[25]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .a ({new_AGEMA_signal_4661, new_AGEMA_signal_4659}), .b ({new_AGEMA_signal_1993, Midori_rounds_sub_sBox_PRINCE_12_n2}), .clk (clk), .r (Fresh[211]), .c ({new_AGEMA_signal_2128, Midori_rounds_sub_sBox_PRINCE_12_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .a ({new_AGEMA_signal_4669, new_AGEMA_signal_4667}), .b ({new_AGEMA_signal_2130, Midori_rounds_sub_sBox_PRINCE_13_n14}), .clk (clk), .r (Fresh[212]), .c ({new_AGEMA_signal_2196, Midori_rounds_SR_Result[7]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .a ({new_AGEMA_signal_1995, Midori_rounds_sub_sBox_PRINCE_13_n11}), .b ({new_AGEMA_signal_4673, new_AGEMA_signal_4671}), .clk (clk), .r (Fresh[213]), .c ({new_AGEMA_signal_2131, Midori_rounds_sub_sBox_PRINCE_13_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .a ({new_AGEMA_signal_4677, new_AGEMA_signal_4675}), .b ({new_AGEMA_signal_2132, Midori_rounds_sub_sBox_PRINCE_13_n5}), .clk (clk), .r (Fresh[214]), .c ({new_AGEMA_signal_2198, Midori_rounds_SR_Result[5]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .a ({new_AGEMA_signal_4673, new_AGEMA_signal_4671}), .b ({new_AGEMA_signal_1999, Midori_rounds_sub_sBox_PRINCE_13_n2}), .clk (clk), .r (Fresh[215]), .c ({new_AGEMA_signal_2133, Midori_rounds_sub_sBox_PRINCE_13_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .a ({new_AGEMA_signal_4681, new_AGEMA_signal_4679}), .b ({new_AGEMA_signal_2135, Midori_rounds_sub_sBox_PRINCE_14_n14}), .clk (clk), .r (Fresh[216]), .c ({new_AGEMA_signal_2200, Midori_rounds_SR_Result[35]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .a ({new_AGEMA_signal_2001, Midori_rounds_sub_sBox_PRINCE_14_n11}), .b ({new_AGEMA_signal_4685, new_AGEMA_signal_4683}), .clk (clk), .r (Fresh[217]), .c ({new_AGEMA_signal_2136, Midori_rounds_sub_sBox_PRINCE_14_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .a ({new_AGEMA_signal_4689, new_AGEMA_signal_4687}), .b ({new_AGEMA_signal_2137, Midori_rounds_sub_sBox_PRINCE_14_n5}), .clk (clk), .r (Fresh[218]), .c ({new_AGEMA_signal_2202, Midori_rounds_SR_Result[33]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .a ({new_AGEMA_signal_4685, new_AGEMA_signal_4683}), .b ({new_AGEMA_signal_2005, Midori_rounds_sub_sBox_PRINCE_14_n2}), .clk (clk), .r (Fresh[219]), .c ({new_AGEMA_signal_2138, Midori_rounds_sub_sBox_PRINCE_14_n3}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .a ({new_AGEMA_signal_4693, new_AGEMA_signal_4691}), .b ({new_AGEMA_signal_2140, Midori_rounds_sub_sBox_PRINCE_15_n14}), .clk (clk), .r (Fresh[220]), .c ({new_AGEMA_signal_2204, Midori_rounds_SR_Result[63]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .a ({new_AGEMA_signal_2007, Midori_rounds_sub_sBox_PRINCE_15_n11}), .b ({new_AGEMA_signal_4697, new_AGEMA_signal_4695}), .clk (clk), .r (Fresh[221]), .c ({new_AGEMA_signal_2141, Midori_rounds_sub_sBox_PRINCE_15_n12}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .a ({new_AGEMA_signal_4701, new_AGEMA_signal_4699}), .b ({new_AGEMA_signal_2142, Midori_rounds_sub_sBox_PRINCE_15_n5}), .clk (clk), .r (Fresh[222]), .c ({new_AGEMA_signal_2206, Midori_rounds_SR_Result[61]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .a ({new_AGEMA_signal_4697, new_AGEMA_signal_4695}), .b ({new_AGEMA_signal_2011, Midori_rounds_sub_sBox_PRINCE_15_n2}), .clk (clk), .r (Fresh[223]), .c ({new_AGEMA_signal_2143, Midori_rounds_sub_sBox_PRINCE_15_n3}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_1_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2174, Midori_rounds_SR_Result[1]}), .a ({new_AGEMA_signal_2311, Midori_rounds_sub_ResultXORkey[1]}), .c ({new_AGEMA_signal_2320, Midori_rounds_mul_input[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_3_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2172, Midori_rounds_SR_Result[3]}), .a ({new_AGEMA_signal_2294, Midori_rounds_sub_ResultXORkey[3]}), .c ({new_AGEMA_signal_2322, Midori_rounds_mul_input[3]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_5_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2198, Midori_rounds_SR_Result[5]}), .a ({new_AGEMA_signal_2278, Midori_rounds_sub_ResultXORkey[5]}), .c ({new_AGEMA_signal_2323, Midori_rounds_mul_input[5]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_7_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2196, Midori_rounds_SR_Result[7]}), .a ({new_AGEMA_signal_2273, Midori_rounds_sub_ResultXORkey[7]}), .c ({new_AGEMA_signal_2325, Midori_rounds_mul_input[7]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_9_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2154, Midori_rounds_SR_Result[9]}), .a ({new_AGEMA_signal_2272, Midori_rounds_sub_ResultXORkey[9]}), .c ({new_AGEMA_signal_2326, Midori_rounds_mul_input[9]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_11_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2152, Midori_rounds_SR_Result[11]}), .a ({new_AGEMA_signal_2318, Midori_rounds_sub_ResultXORkey[11]}), .c ({new_AGEMA_signal_2328, Midori_rounds_mul_input[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_13_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2178, Midori_rounds_SR_Result[13]}), .a ({new_AGEMA_signal_2317, Midori_rounds_sub_ResultXORkey[13]}), .c ({new_AGEMA_signal_2329, Midori_rounds_mul_input[13]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_15_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2176, Midori_rounds_SR_Result[15]}), .a ({new_AGEMA_signal_2315, Midori_rounds_sub_ResultXORkey[15]}), .c ({new_AGEMA_signal_2331, Midori_rounds_mul_input[15]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_17_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2182, Midori_rounds_SR_Result[17]}), .a ({new_AGEMA_signal_2314, Midori_rounds_sub_ResultXORkey[17]}), .c ({new_AGEMA_signal_2332, Midori_rounds_mul_input[17]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_19_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2180, Midori_rounds_SR_Result[19]}), .a ({new_AGEMA_signal_2312, Midori_rounds_sub_ResultXORkey[19]}), .c ({new_AGEMA_signal_2334, Midori_rounds_mul_input[19]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_21_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2158, Midori_rounds_SR_Result[21]}), .a ({new_AGEMA_signal_2310, Midori_rounds_sub_ResultXORkey[21]}), .c ({new_AGEMA_signal_2335, Midori_rounds_mul_input[21]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_23_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2156, Midori_rounds_SR_Result[23]}), .a ({new_AGEMA_signal_2308, Midori_rounds_sub_ResultXORkey[23]}), .c ({new_AGEMA_signal_2337, Midori_rounds_mul_input[23]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_25_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2194, Midori_rounds_SR_Result[25]}), .a ({new_AGEMA_signal_2307, Midori_rounds_sub_ResultXORkey[25]}), .c ({new_AGEMA_signal_2338, Midori_rounds_mul_input[25]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_27_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2192, Midori_rounds_SR_Result[27]}), .a ({new_AGEMA_signal_2305, Midori_rounds_sub_ResultXORkey[27]}), .c ({new_AGEMA_signal_2340, Midori_rounds_mul_input[27]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_29_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2170, Midori_rounds_SR_Result[29]}), .a ({new_AGEMA_signal_2304, Midori_rounds_sub_ResultXORkey[29]}), .c ({new_AGEMA_signal_2341, Midori_rounds_mul_input[29]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_31_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2168, Midori_rounds_SR_Result[31]}), .a ({new_AGEMA_signal_2301, Midori_rounds_sub_ResultXORkey[31]}), .c ({new_AGEMA_signal_2343, Midori_rounds_mul_input[31]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_33_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2202, Midori_rounds_SR_Result[33]}), .a ({new_AGEMA_signal_2300, Midori_rounds_sub_ResultXORkey[33]}), .c ({new_AGEMA_signal_2344, Midori_rounds_mul_input[33]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_35_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2200, Midori_rounds_SR_Result[35]}), .a ({new_AGEMA_signal_2298, Midori_rounds_sub_ResultXORkey[35]}), .c ({new_AGEMA_signal_2346, Midori_rounds_mul_input[35]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_37_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2162, Midori_rounds_SR_Result[37]}), .a ({new_AGEMA_signal_2297, Midori_rounds_sub_ResultXORkey[37]}), .c ({new_AGEMA_signal_2347, Midori_rounds_mul_input[37]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_39_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2160, Midori_rounds_SR_Result[39]}), .a ({new_AGEMA_signal_2295, Midori_rounds_sub_ResultXORkey[39]}), .c ({new_AGEMA_signal_2349, Midori_rounds_mul_input[39]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_41_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2190, Midori_rounds_SR_Result[41]}), .a ({new_AGEMA_signal_2293, Midori_rounds_sub_ResultXORkey[41]}), .c ({new_AGEMA_signal_2350, Midori_rounds_mul_input[41]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_43_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2188, Midori_rounds_SR_Result[43]}), .a ({new_AGEMA_signal_2291, Midori_rounds_sub_ResultXORkey[43]}), .c ({new_AGEMA_signal_2352, Midori_rounds_mul_input[43]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_45_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2150, Midori_rounds_SR_Result[45]}), .a ({new_AGEMA_signal_2290, Midori_rounds_sub_ResultXORkey[45]}), .c ({new_AGEMA_signal_2353, Midori_rounds_mul_input[45]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_47_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2148, Midori_rounds_SR_Result[47]}), .a ({new_AGEMA_signal_2288, Midori_rounds_sub_ResultXORkey[47]}), .c ({new_AGEMA_signal_2355, Midori_rounds_mul_input[47]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_49_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2146, Midori_rounds_SR_Result[49]}), .a ({new_AGEMA_signal_2287, Midori_rounds_sub_ResultXORkey[49]}), .c ({new_AGEMA_signal_2356, Midori_rounds_mul_input[49]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_51_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2144, Midori_rounds_SR_Result[51]}), .a ({new_AGEMA_signal_2285, Midori_rounds_sub_ResultXORkey[51]}), .c ({new_AGEMA_signal_2358, Midori_rounds_mul_input[51]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_53_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2186, Midori_rounds_SR_Result[53]}), .a ({new_AGEMA_signal_2284, Midori_rounds_sub_ResultXORkey[53]}), .c ({new_AGEMA_signal_2359, Midori_rounds_mul_input[53]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_55_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2184, Midori_rounds_SR_Result[55]}), .a ({new_AGEMA_signal_2282, Midori_rounds_sub_ResultXORkey[55]}), .c ({new_AGEMA_signal_2361, Midori_rounds_mul_input[55]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_57_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2166, Midori_rounds_SR_Result[57]}), .a ({new_AGEMA_signal_2281, Midori_rounds_sub_ResultXORkey[57]}), .c ({new_AGEMA_signal_2362, Midori_rounds_mul_input[57]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_59_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2164, Midori_rounds_SR_Result[59]}), .a ({new_AGEMA_signal_2279, Midori_rounds_sub_ResultXORkey[59]}), .c ({new_AGEMA_signal_2364, Midori_rounds_mul_input[59]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_61_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2206, Midori_rounds_SR_Result[61]}), .a ({new_AGEMA_signal_2277, Midori_rounds_sub_ResultXORkey[61]}), .c ({new_AGEMA_signal_2365, Midori_rounds_mul_input[61]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_63_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2204, Midori_rounds_SR_Result[63]}), .a ({new_AGEMA_signal_2275, Midori_rounds_sub_ResultXORkey[63]}), .c ({new_AGEMA_signal_2367, Midori_rounds_mul_input[63]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U24 ( .a ({new_AGEMA_signal_2365, Midori_rounds_mul_input[61]}), .b ({new_AGEMA_signal_2371, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_2392, Midori_rounds_SR_Inv_Result[21]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U22 ( .a ({new_AGEMA_signal_2358, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_2368, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_2393, Midori_rounds_SR_Inv_Result[43]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U20 ( .a ({new_AGEMA_signal_2356, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_2370, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_2395, Midori_rounds_SR_Inv_Result[41]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U18 ( .a ({new_AGEMA_signal_2361, Midori_rounds_mul_input[55]}), .b ({new_AGEMA_signal_2368, Midori_rounds_mul_MC1_n6}), .c ({new_AGEMA_signal_2396, Midori_rounds_SR_Inv_Result[3]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U17 ( .a ({new_AGEMA_signal_2367, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_2364, Midori_rounds_mul_input[59]}), .c ({new_AGEMA_signal_2368, Midori_rounds_mul_MC1_n6}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U14 ( .a ({new_AGEMA_signal_2359, Midori_rounds_mul_input[53]}), .b ({new_AGEMA_signal_2370, Midori_rounds_mul_MC1_n4}), .c ({new_AGEMA_signal_2398, Midori_rounds_SR_Inv_Result[1]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U13 ( .a ({new_AGEMA_signal_2362, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_2365, Midori_rounds_mul_input[61]}), .c ({new_AGEMA_signal_2370, Midori_rounds_mul_MC1_n4}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U12 ( .a ({new_AGEMA_signal_2364, Midori_rounds_mul_input[59]}), .b ({new_AGEMA_signal_2372, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_2399, Midori_rounds_SR_Inv_Result[63]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U10 ( .a ({new_AGEMA_signal_2362, Midori_rounds_mul_input[57]}), .b ({new_AGEMA_signal_2371, Midori_rounds_mul_MC1_n8}), .c ({new_AGEMA_signal_2401, Midori_rounds_SR_Inv_Result[61]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U9 ( .a ({new_AGEMA_signal_2356, Midori_rounds_mul_input[49]}), .b ({new_AGEMA_signal_2359, Midori_rounds_mul_input[53]}), .c ({new_AGEMA_signal_2371, Midori_rounds_mul_MC1_n8}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U6 ( .a ({new_AGEMA_signal_2367, Midori_rounds_mul_input[63]}), .b ({new_AGEMA_signal_2372, Midori_rounds_mul_MC1_n2}), .c ({new_AGEMA_signal_2402, Midori_rounds_SR_Inv_Result[23]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U5 ( .a ({new_AGEMA_signal_2358, Midori_rounds_mul_input[51]}), .b ({new_AGEMA_signal_2361, Midori_rounds_mul_input[55]}), .c ({new_AGEMA_signal_2372, Midori_rounds_mul_MC1_n2}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U24 ( .a ({new_AGEMA_signal_2353, Midori_rounds_mul_input[45]}), .b ({new_AGEMA_signal_2377, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_2404, Midori_rounds_SR_Inv_Result[45]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U22 ( .a ({new_AGEMA_signal_2346, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_2374, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_2405, Midori_rounds_SR_Inv_Result[19]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U20 ( .a ({new_AGEMA_signal_2344, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_2376, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_2407, Midori_rounds_SR_Inv_Result[17]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U18 ( .a ({new_AGEMA_signal_2349, Midori_rounds_mul_input[39]}), .b ({new_AGEMA_signal_2374, Midori_rounds_mul_MC2_n6}), .c ({new_AGEMA_signal_2408, Midori_rounds_SR_Inv_Result[59]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U17 ( .a ({new_AGEMA_signal_2355, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_2352, Midori_rounds_mul_input[43]}), .c ({new_AGEMA_signal_2374, Midori_rounds_mul_MC2_n6}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U14 ( .a ({new_AGEMA_signal_2347, Midori_rounds_mul_input[37]}), .b ({new_AGEMA_signal_2376, Midori_rounds_mul_MC2_n4}), .c ({new_AGEMA_signal_2410, Midori_rounds_SR_Inv_Result[57]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U13 ( .a ({new_AGEMA_signal_2350, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_2353, Midori_rounds_mul_input[45]}), .c ({new_AGEMA_signal_2376, Midori_rounds_mul_MC2_n4}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U12 ( .a ({new_AGEMA_signal_2352, Midori_rounds_mul_input[43]}), .b ({new_AGEMA_signal_2378, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_2411, Midori_rounds_SR_Inv_Result[7]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U10 ( .a ({new_AGEMA_signal_2350, Midori_rounds_mul_input[41]}), .b ({new_AGEMA_signal_2377, Midori_rounds_mul_MC2_n8}), .c ({new_AGEMA_signal_2413, Midori_rounds_SR_Inv_Result[5]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U9 ( .a ({new_AGEMA_signal_2344, Midori_rounds_mul_input[33]}), .b ({new_AGEMA_signal_2347, Midori_rounds_mul_input[37]}), .c ({new_AGEMA_signal_2377, Midori_rounds_mul_MC2_n8}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U6 ( .a ({new_AGEMA_signal_2355, Midori_rounds_mul_input[47]}), .b ({new_AGEMA_signal_2378, Midori_rounds_mul_MC2_n2}), .c ({new_AGEMA_signal_2414, Midori_rounds_SR_Inv_Result[47]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U5 ( .a ({new_AGEMA_signal_2346, Midori_rounds_mul_input[35]}), .b ({new_AGEMA_signal_2349, Midori_rounds_mul_input[39]}), .c ({new_AGEMA_signal_2378, Midori_rounds_mul_MC2_n2}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U24 ( .a ({new_AGEMA_signal_2341, Midori_rounds_mul_input[29]}), .b ({new_AGEMA_signal_2383, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_2416, Midori_rounds_SR_Inv_Result[49]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U22 ( .a ({new_AGEMA_signal_2334, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_2380, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_2417, Midori_rounds_SR_Inv_Result[15]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U20 ( .a ({new_AGEMA_signal_2332, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_2382, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_2419, Midori_rounds_SR_Inv_Result[13]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U18 ( .a ({new_AGEMA_signal_2337, Midori_rounds_mul_input[23]}), .b ({new_AGEMA_signal_2380, Midori_rounds_mul_MC3_n6}), .c ({new_AGEMA_signal_2420, Midori_rounds_SR_Inv_Result[39]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U17 ( .a ({new_AGEMA_signal_2343, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_2340, Midori_rounds_mul_input[27]}), .c ({new_AGEMA_signal_2380, Midori_rounds_mul_MC3_n6}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U14 ( .a ({new_AGEMA_signal_2335, Midori_rounds_mul_input[21]}), .b ({new_AGEMA_signal_2382, Midori_rounds_mul_MC3_n4}), .c ({new_AGEMA_signal_2422, Midori_rounds_SR_Inv_Result[37]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U13 ( .a ({new_AGEMA_signal_2338, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_2341, Midori_rounds_mul_input[29]}), .c ({new_AGEMA_signal_2382, Midori_rounds_mul_MC3_n4}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U12 ( .a ({new_AGEMA_signal_2340, Midori_rounds_mul_input[27]}), .b ({new_AGEMA_signal_2384, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_2423, Midori_rounds_SR_Inv_Result[27]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U10 ( .a ({new_AGEMA_signal_2338, Midori_rounds_mul_input[25]}), .b ({new_AGEMA_signal_2383, Midori_rounds_mul_MC3_n8}), .c ({new_AGEMA_signal_2425, Midori_rounds_SR_Inv_Result[25]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U9 ( .a ({new_AGEMA_signal_2332, Midori_rounds_mul_input[17]}), .b ({new_AGEMA_signal_2335, Midori_rounds_mul_input[21]}), .c ({new_AGEMA_signal_2383, Midori_rounds_mul_MC3_n8}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U6 ( .a ({new_AGEMA_signal_2343, Midori_rounds_mul_input[31]}), .b ({new_AGEMA_signal_2384, Midori_rounds_mul_MC3_n2}), .c ({new_AGEMA_signal_2426, Midori_rounds_SR_Inv_Result[51]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U5 ( .a ({new_AGEMA_signal_2334, Midori_rounds_mul_input[19]}), .b ({new_AGEMA_signal_2337, Midori_rounds_mul_input[23]}), .c ({new_AGEMA_signal_2384, Midori_rounds_mul_MC3_n2}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U24 ( .a ({new_AGEMA_signal_2329, Midori_rounds_mul_input[13]}), .b ({new_AGEMA_signal_2389, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_2428, Midori_rounds_SR_Inv_Result[9]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U22 ( .a ({new_AGEMA_signal_2322, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_2386, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_2429, Midori_rounds_SR_Inv_Result[55]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U20 ( .a ({new_AGEMA_signal_2320, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_2388, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_2431, Midori_rounds_SR_Inv_Result[53]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U18 ( .a ({new_AGEMA_signal_2325, Midori_rounds_mul_input[7]}), .b ({new_AGEMA_signal_2386, Midori_rounds_mul_MC4_n6}), .c ({new_AGEMA_signal_2432, Midori_rounds_SR_Inv_Result[31]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U17 ( .a ({new_AGEMA_signal_2331, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_2328, Midori_rounds_mul_input[11]}), .c ({new_AGEMA_signal_2386, Midori_rounds_mul_MC4_n6}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U14 ( .a ({new_AGEMA_signal_2323, Midori_rounds_mul_input[5]}), .b ({new_AGEMA_signal_2388, Midori_rounds_mul_MC4_n4}), .c ({new_AGEMA_signal_2434, Midori_rounds_SR_Inv_Result[29]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U13 ( .a ({new_AGEMA_signal_2326, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_2329, Midori_rounds_mul_input[13]}), .c ({new_AGEMA_signal_2388, Midori_rounds_mul_MC4_n4}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U12 ( .a ({new_AGEMA_signal_2328, Midori_rounds_mul_input[11]}), .b ({new_AGEMA_signal_2390, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_2435, Midori_rounds_SR_Inv_Result[35]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U10 ( .a ({new_AGEMA_signal_2326, Midori_rounds_mul_input[9]}), .b ({new_AGEMA_signal_2389, Midori_rounds_mul_MC4_n8}), .c ({new_AGEMA_signal_2437, Midori_rounds_SR_Inv_Result[33]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U9 ( .a ({new_AGEMA_signal_2320, Midori_rounds_mul_input[1]}), .b ({new_AGEMA_signal_2323, Midori_rounds_mul_input[5]}), .c ({new_AGEMA_signal_2389, Midori_rounds_mul_MC4_n8}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U6 ( .a ({new_AGEMA_signal_2331, Midori_rounds_mul_input[15]}), .b ({new_AGEMA_signal_2390, Midori_rounds_mul_MC4_n2}), .c ({new_AGEMA_signal_2438, Midori_rounds_SR_Inv_Result[11]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U5 ( .a ({new_AGEMA_signal_2322, Midori_rounds_mul_input[3]}), .b ({new_AGEMA_signal_2325, Midori_rounds_mul_input[7]}), .c ({new_AGEMA_signal_2390, Midori_rounds_mul_MC4_n2}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_1_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2483, Midori_rounds_mul_ResultXORkey[1]}), .a ({new_AGEMA_signal_2398, Midori_rounds_SR_Inv_Result[1]}), .c ({new_AGEMA_signal_2506, Midori_rounds_round_Result[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_3_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2464, Midori_rounds_mul_ResultXORkey[3]}), .a ({new_AGEMA_signal_2396, Midori_rounds_SR_Inv_Result[3]}), .c ({new_AGEMA_signal_2508, Midori_rounds_round_Result[3]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_5_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2447, Midori_rounds_mul_ResultXORkey[5]}), .a ({new_AGEMA_signal_2413, Midori_rounds_SR_Inv_Result[5]}), .c ({new_AGEMA_signal_2509, Midori_rounds_round_Result[5]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_7_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2442, Midori_rounds_mul_ResultXORkey[7]}), .a ({new_AGEMA_signal_2411, Midori_rounds_SR_Inv_Result[7]}), .c ({new_AGEMA_signal_2511, Midori_rounds_round_Result[7]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_9_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2440, Midori_rounds_mul_ResultXORkey[9]}), .a ({new_AGEMA_signal_2428, Midori_rounds_SR_Inv_Result[9]}), .c ({new_AGEMA_signal_2512, Midori_rounds_round_Result[9]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_11_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2490, Midori_rounds_mul_ResultXORkey[11]}), .a ({new_AGEMA_signal_2438, Midori_rounds_SR_Inv_Result[11]}), .c ({new_AGEMA_signal_2514, Midori_rounds_round_Result[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_13_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2489, Midori_rounds_mul_ResultXORkey[13]}), .a ({new_AGEMA_signal_2419, Midori_rounds_SR_Inv_Result[13]}), .c ({new_AGEMA_signal_2515, Midori_rounds_round_Result[13]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_15_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2487, Midori_rounds_mul_ResultXORkey[15]}), .a ({new_AGEMA_signal_2417, Midori_rounds_SR_Inv_Result[15]}), .c ({new_AGEMA_signal_2517, Midori_rounds_round_Result[15]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_17_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2486, Midori_rounds_mul_ResultXORkey[17]}), .a ({new_AGEMA_signal_2407, Midori_rounds_SR_Inv_Result[17]}), .c ({new_AGEMA_signal_2518, Midori_rounds_round_Result[17]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_19_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2484, Midori_rounds_mul_ResultXORkey[19]}), .a ({new_AGEMA_signal_2405, Midori_rounds_SR_Inv_Result[19]}), .c ({new_AGEMA_signal_2520, Midori_rounds_round_Result[19]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_21_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2481, Midori_rounds_mul_ResultXORkey[21]}), .a ({new_AGEMA_signal_2392, Midori_rounds_SR_Inv_Result[21]}), .c ({new_AGEMA_signal_2521, Midori_rounds_round_Result[21]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_23_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2479, Midori_rounds_mul_ResultXORkey[23]}), .a ({new_AGEMA_signal_2402, Midori_rounds_SR_Inv_Result[23]}), .c ({new_AGEMA_signal_2523, Midori_rounds_round_Result[23]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_25_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2478, Midori_rounds_mul_ResultXORkey[25]}), .a ({new_AGEMA_signal_2425, Midori_rounds_SR_Inv_Result[25]}), .c ({new_AGEMA_signal_2524, Midori_rounds_round_Result[25]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_27_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2476, Midori_rounds_mul_ResultXORkey[27]}), .a ({new_AGEMA_signal_2423, Midori_rounds_SR_Inv_Result[27]}), .c ({new_AGEMA_signal_2526, Midori_rounds_round_Result[27]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_29_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2475, Midori_rounds_mul_ResultXORkey[29]}), .a ({new_AGEMA_signal_2434, Midori_rounds_SR_Inv_Result[29]}), .c ({new_AGEMA_signal_2527, Midori_rounds_round_Result[29]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_31_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2472, Midori_rounds_mul_ResultXORkey[31]}), .a ({new_AGEMA_signal_2432, Midori_rounds_SR_Inv_Result[31]}), .c ({new_AGEMA_signal_2529, Midori_rounds_round_Result[31]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_33_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2471, Midori_rounds_mul_ResultXORkey[33]}), .a ({new_AGEMA_signal_2437, Midori_rounds_SR_Inv_Result[33]}), .c ({new_AGEMA_signal_2530, Midori_rounds_round_Result[33]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_35_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2469, Midori_rounds_mul_ResultXORkey[35]}), .a ({new_AGEMA_signal_2435, Midori_rounds_SR_Inv_Result[35]}), .c ({new_AGEMA_signal_2532, Midori_rounds_round_Result[35]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_37_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2467, Midori_rounds_mul_ResultXORkey[37]}), .a ({new_AGEMA_signal_2422, Midori_rounds_SR_Inv_Result[37]}), .c ({new_AGEMA_signal_2533, Midori_rounds_round_Result[37]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_39_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2465, Midori_rounds_mul_ResultXORkey[39]}), .a ({new_AGEMA_signal_2420, Midori_rounds_SR_Inv_Result[39]}), .c ({new_AGEMA_signal_2535, Midori_rounds_round_Result[39]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_41_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2463, Midori_rounds_mul_ResultXORkey[41]}), .a ({new_AGEMA_signal_2395, Midori_rounds_SR_Inv_Result[41]}), .c ({new_AGEMA_signal_2536, Midori_rounds_round_Result[41]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_43_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2461, Midori_rounds_mul_ResultXORkey[43]}), .a ({new_AGEMA_signal_2393, Midori_rounds_SR_Inv_Result[43]}), .c ({new_AGEMA_signal_2538, Midori_rounds_round_Result[43]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_45_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2459, Midori_rounds_mul_ResultXORkey[45]}), .a ({new_AGEMA_signal_2404, Midori_rounds_SR_Inv_Result[45]}), .c ({new_AGEMA_signal_2539, Midori_rounds_round_Result[45]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_47_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2457, Midori_rounds_mul_ResultXORkey[47]}), .a ({new_AGEMA_signal_2414, Midori_rounds_SR_Inv_Result[47]}), .c ({new_AGEMA_signal_2541, Midori_rounds_round_Result[47]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_49_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2456, Midori_rounds_mul_ResultXORkey[49]}), .a ({new_AGEMA_signal_2416, Midori_rounds_SR_Inv_Result[49]}), .c ({new_AGEMA_signal_2542, Midori_rounds_round_Result[49]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_51_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2454, Midori_rounds_mul_ResultXORkey[51]}), .a ({new_AGEMA_signal_2426, Midori_rounds_SR_Inv_Result[51]}), .c ({new_AGEMA_signal_2544, Midori_rounds_round_Result[51]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_53_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2453, Midori_rounds_mul_ResultXORkey[53]}), .a ({new_AGEMA_signal_2431, Midori_rounds_SR_Inv_Result[53]}), .c ({new_AGEMA_signal_2545, Midori_rounds_round_Result[53]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_55_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2451, Midori_rounds_mul_ResultXORkey[55]}), .a ({new_AGEMA_signal_2429, Midori_rounds_SR_Inv_Result[55]}), .c ({new_AGEMA_signal_2547, Midori_rounds_round_Result[55]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_57_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2450, Midori_rounds_mul_ResultXORkey[57]}), .a ({new_AGEMA_signal_2410, Midori_rounds_SR_Inv_Result[57]}), .c ({new_AGEMA_signal_2548, Midori_rounds_round_Result[57]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_59_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2448, Midori_rounds_mul_ResultXORkey[59]}), .a ({new_AGEMA_signal_2408, Midori_rounds_SR_Inv_Result[59]}), .c ({new_AGEMA_signal_2550, Midori_rounds_round_Result[59]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_61_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2446, Midori_rounds_mul_ResultXORkey[61]}), .a ({new_AGEMA_signal_2401, Midori_rounds_SR_Inv_Result[61]}), .c ({new_AGEMA_signal_2551, Midori_rounds_round_Result[61]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_63_U1 ( .s (new_AGEMA_signal_4707), .b ({new_AGEMA_signal_2444, Midori_rounds_mul_ResultXORkey[63]}), .a ({new_AGEMA_signal_2399, Midori_rounds_SR_Inv_Result[63]}), .c ({new_AGEMA_signal_2553, Midori_rounds_round_Result[63]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_3029), .Q (new_AGEMA_signal_3030) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (clk), .D (new_AGEMA_signal_3356), .Q (new_AGEMA_signal_3357) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (clk), .D (new_AGEMA_signal_3362), .Q (new_AGEMA_signal_3363) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (clk), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_3369) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (clk), .D (new_AGEMA_signal_3374), .Q (new_AGEMA_signal_3375) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (clk), .D (new_AGEMA_signal_3380), .Q (new_AGEMA_signal_3381) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (clk), .D (new_AGEMA_signal_3386), .Q (new_AGEMA_signal_3387) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (clk), .D (new_AGEMA_signal_3392), .Q (new_AGEMA_signal_3393) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (clk), .D (new_AGEMA_signal_3398), .Q (new_AGEMA_signal_3399) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (clk), .D (new_AGEMA_signal_3404), .Q (new_AGEMA_signal_3405) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (clk), .D (new_AGEMA_signal_3410), .Q (new_AGEMA_signal_3411) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (clk), .D (new_AGEMA_signal_3416), .Q (new_AGEMA_signal_3417) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (clk), .D (new_AGEMA_signal_3422), .Q (new_AGEMA_signal_3423) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (clk), .D (new_AGEMA_signal_3428), .Q (new_AGEMA_signal_3429) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (clk), .D (new_AGEMA_signal_3434), .Q (new_AGEMA_signal_3435) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (clk), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_3441) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (clk), .D (new_AGEMA_signal_3446), .Q (new_AGEMA_signal_3447) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (clk), .D (new_AGEMA_signal_3452), .Q (new_AGEMA_signal_3453) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (clk), .D (new_AGEMA_signal_3458), .Q (new_AGEMA_signal_3459) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (clk), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_3465) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (clk), .D (new_AGEMA_signal_3470), .Q (new_AGEMA_signal_3471) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (clk), .D (new_AGEMA_signal_3476), .Q (new_AGEMA_signal_3477) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (clk), .D (new_AGEMA_signal_3482), .Q (new_AGEMA_signal_3483) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (clk), .D (new_AGEMA_signal_3488), .Q (new_AGEMA_signal_3489) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (clk), .D (new_AGEMA_signal_3494), .Q (new_AGEMA_signal_3495) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (clk), .D (new_AGEMA_signal_3500), .Q (new_AGEMA_signal_3501) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (clk), .D (new_AGEMA_signal_3506), .Q (new_AGEMA_signal_3507) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (clk), .D (new_AGEMA_signal_3512), .Q (new_AGEMA_signal_3513) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (clk), .D (new_AGEMA_signal_3518), .Q (new_AGEMA_signal_3519) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (clk), .D (new_AGEMA_signal_3524), .Q (new_AGEMA_signal_3525) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (clk), .D (new_AGEMA_signal_3530), .Q (new_AGEMA_signal_3531) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (clk), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_3537) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (clk), .D (new_AGEMA_signal_3542), .Q (new_AGEMA_signal_3543) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (clk), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_3549) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (clk), .D (new_AGEMA_signal_3554), .Q (new_AGEMA_signal_3555) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (clk), .D (new_AGEMA_signal_3560), .Q (new_AGEMA_signal_3561) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (clk), .D (new_AGEMA_signal_3566), .Q (new_AGEMA_signal_3567) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (clk), .D (new_AGEMA_signal_3572), .Q (new_AGEMA_signal_3573) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (clk), .D (new_AGEMA_signal_3578), .Q (new_AGEMA_signal_3579) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (clk), .D (new_AGEMA_signal_3584), .Q (new_AGEMA_signal_3585) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (clk), .D (new_AGEMA_signal_3590), .Q (new_AGEMA_signal_3591) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (clk), .D (new_AGEMA_signal_3596), .Q (new_AGEMA_signal_3597) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (clk), .D (new_AGEMA_signal_3602), .Q (new_AGEMA_signal_3603) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (clk), .D (new_AGEMA_signal_3608), .Q (new_AGEMA_signal_3609) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (clk), .D (new_AGEMA_signal_3614), .Q (new_AGEMA_signal_3615) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (clk), .D (new_AGEMA_signal_3620), .Q (new_AGEMA_signal_3621) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (clk), .D (new_AGEMA_signal_3626), .Q (new_AGEMA_signal_3627) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (clk), .D (new_AGEMA_signal_3632), .Q (new_AGEMA_signal_3633) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (clk), .D (new_AGEMA_signal_3638), .Q (new_AGEMA_signal_3639) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (clk), .D (new_AGEMA_signal_3644), .Q (new_AGEMA_signal_3645) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (clk), .D (new_AGEMA_signal_3650), .Q (new_AGEMA_signal_3651) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (clk), .D (new_AGEMA_signal_3656), .Q (new_AGEMA_signal_3657) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (clk), .D (new_AGEMA_signal_3662), .Q (new_AGEMA_signal_3663) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (clk), .D (new_AGEMA_signal_3668), .Q (new_AGEMA_signal_3669) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (clk), .D (new_AGEMA_signal_3674), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (clk), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (clk), .D (new_AGEMA_signal_3686), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (clk), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (clk), .D (new_AGEMA_signal_3698), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (clk), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (clk), .D (new_AGEMA_signal_3710), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (clk), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (clk), .D (new_AGEMA_signal_3722), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (clk), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (clk), .D (new_AGEMA_signal_3734), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (clk), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (clk), .D (new_AGEMA_signal_3746), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (clk), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (clk), .D (new_AGEMA_signal_3758), .Q (new_AGEMA_signal_3759) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (clk), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_3765) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_3770), .Q (new_AGEMA_signal_3771) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_3776), .Q (new_AGEMA_signal_3777) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_3782), .Q (new_AGEMA_signal_3783) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_3788), .Q (new_AGEMA_signal_3789) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_3794), .Q (new_AGEMA_signal_3795) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_3800), .Q (new_AGEMA_signal_3801) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_3806), .Q (new_AGEMA_signal_3807) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_3813) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_3818), .Q (new_AGEMA_signal_3819) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_3824), .Q (new_AGEMA_signal_3825) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_3830), .Q (new_AGEMA_signal_3831) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_3837) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_3842), .Q (new_AGEMA_signal_3843) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_3848), .Q (new_AGEMA_signal_3849) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_3855) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_3861) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_3866), .Q (new_AGEMA_signal_3867) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_3872), .Q (new_AGEMA_signal_3873) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_3879) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_3885) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_3890), .Q (new_AGEMA_signal_3891) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_3914), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_3938), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_3962), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_4010), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_4034), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_4058), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_4082), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_4106), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_4130), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_4202), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_4226), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_4250), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_4274), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_4371) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_4376), .Q (new_AGEMA_signal_4377) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_4382), .Q (new_AGEMA_signal_4383) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_4388), .Q (new_AGEMA_signal_4389) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_4394), .Q (new_AGEMA_signal_4395) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_4400), .Q (new_AGEMA_signal_4401) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_4406), .Q (new_AGEMA_signal_4407) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_4412), .Q (new_AGEMA_signal_4413) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_4418), .Q (new_AGEMA_signal_4419) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_4424), .Q (new_AGEMA_signal_4425) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_4430), .Q (new_AGEMA_signal_4431) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_4436), .Q (new_AGEMA_signal_4437) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_4442), .Q (new_AGEMA_signal_4443) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_4448), .Q (new_AGEMA_signal_4449) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_4454), .Q (new_AGEMA_signal_4455) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_4460), .Q (new_AGEMA_signal_4461) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_4466), .Q (new_AGEMA_signal_4467) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_4472), .Q (new_AGEMA_signal_4473) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_4478), .Q (new_AGEMA_signal_4479) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_4484), .Q (new_AGEMA_signal_4485) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_4490), .Q (new_AGEMA_signal_4491) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_4496), .Q (new_AGEMA_signal_4497) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_4502), .Q (new_AGEMA_signal_4503) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_4508), .Q (new_AGEMA_signal_4509) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_4707) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_4713) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_4728), .Q (new_AGEMA_signal_4729) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_4848), .Q (new_AGEMA_signal_4849) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_4872), .Q (new_AGEMA_signal_4873) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_4889) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_4896), .Q (new_AGEMA_signal_4897) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_4905) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_4913) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_4920), .Q (new_AGEMA_signal_4921) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_4929) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_4944), .Q (new_AGEMA_signal_4945) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_4952), .Q (new_AGEMA_signal_4953) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_4961) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_4968), .Q (new_AGEMA_signal_4969) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_4976), .Q (new_AGEMA_signal_4977) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_4985) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_4992), .Q (new_AGEMA_signal_4993) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_5000), .Q (new_AGEMA_signal_5001) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_5009) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_5016), .Q (new_AGEMA_signal_5017) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_5024), .Q (new_AGEMA_signal_5025) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_5033) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_5041) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_5048), .Q (new_AGEMA_signal_5049) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_5057) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_5065) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_5072), .Q (new_AGEMA_signal_5073) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_5081) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_5088), .Q (new_AGEMA_signal_5089) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_5096), .Q (new_AGEMA_signal_5097) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_5105) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_5112), .Q (new_AGEMA_signal_5113) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_5120), .Q (new_AGEMA_signal_5121) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_5129) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_5136), .Q (new_AGEMA_signal_5137) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_5144), .Q (new_AGEMA_signal_5145) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_5153) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_5161) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_5168), .Q (new_AGEMA_signal_5169) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_5177) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_5185) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_5192), .Q (new_AGEMA_signal_5193) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_5201) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_5208), .Q (new_AGEMA_signal_5209) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_5216), .Q (new_AGEMA_signal_5217) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_5225) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_5233) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_5240), .Q (new_AGEMA_signal_5241) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_5249) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_5257) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_5264), .Q (new_AGEMA_signal_5265) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_5273) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_5280), .Q (new_AGEMA_signal_5281) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_5288), .Q (new_AGEMA_signal_5289) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_5297) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_5304), .Q (new_AGEMA_signal_5305) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_5312), .Q (new_AGEMA_signal_5313) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_5321) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_5328), .Q (new_AGEMA_signal_5329) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_5336), .Q (new_AGEMA_signal_5337) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_5345) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_5352), .Q (new_AGEMA_signal_5353) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_5360), .Q (new_AGEMA_signal_5361) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_5368), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_5385) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_5401) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_5409) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_5425) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_5739) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_5747) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_5754), .Q (new_AGEMA_signal_5755) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_5763) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_5771) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_5778), .Q (new_AGEMA_signal_5779) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_5787) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_5795) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_5803) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_5811) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_5818), .Q (new_AGEMA_signal_5819) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_5827) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_5835) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_5842), .Q (new_AGEMA_signal_5843) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_5851) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_5859) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_5866), .Q (new_AGEMA_signal_5867) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_5875) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_5883) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_5891) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_5899) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_5907) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_5915) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_5923) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_5931) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_5938), .Q (new_AGEMA_signal_5939) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_5947) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_5955) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_5962), .Q (new_AGEMA_signal_5963) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_5971) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_5979) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_5986), .Q (new_AGEMA_signal_5987) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_5995) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_6003) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_6011) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_6019) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_6027) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_6035) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_6043) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_6051) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_6058), .Q (new_AGEMA_signal_6059) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_6067) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_6075) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_6082), .Q (new_AGEMA_signal_6083) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_6091) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_6099) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_6106), .Q (new_AGEMA_signal_6107) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_6114), .Q (new_AGEMA_signal_6115) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_6123) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_6130), .Q (new_AGEMA_signal_6131) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_6138), .Q (new_AGEMA_signal_6139) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_6147) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_6155) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_6163) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_6171) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_6178), .Q (new_AGEMA_signal_6179) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_6187) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_6195) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_6202), .Q (new_AGEMA_signal_6203) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_6210), .Q (new_AGEMA_signal_6211) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_6219) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_6226), .Q (new_AGEMA_signal_6227) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_6234), .Q (new_AGEMA_signal_6235) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_6243) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_6259) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_6281) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_6283) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_6292), .Q (new_AGEMA_signal_6293) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_6301) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_6305) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_6307) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_6317) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_6319) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_6321) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_6325) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_6329) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_6331) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_6333) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_6337) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_6340), .Q (new_AGEMA_signal_6341) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_6343) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_6345) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_6349) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_6353) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_6355) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_6365) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_6367) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_6369) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_6373) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_6377) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_6379) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_6381) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_6385) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_6389) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_6391) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_6393) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_6397) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_6401) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_6403) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_6413) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_6415) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_6417) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_6421) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_6424), .Q (new_AGEMA_signal_6425) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_6426), .Q (new_AGEMA_signal_6427) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_6429) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_6433) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_6437) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_6445) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_6461) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_6469) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_2960), .Q (new_AGEMA_signal_2961) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_2962), .Q (new_AGEMA_signal_2963) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_2964), .Q (new_AGEMA_signal_2965) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_2966), .Q (new_AGEMA_signal_2967) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_2968), .Q (new_AGEMA_signal_2969) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_2970), .Q (new_AGEMA_signal_2971) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_2972), .Q (new_AGEMA_signal_2973) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_2974), .Q (new_AGEMA_signal_2975) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_2976), .Q (new_AGEMA_signal_2977) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_2978), .Q (new_AGEMA_signal_2979) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_2980), .Q (new_AGEMA_signal_2981) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_2982), .Q (new_AGEMA_signal_2983) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_2984), .Q (new_AGEMA_signal_2985) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_2986), .Q (new_AGEMA_signal_2987) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_2988), .Q (new_AGEMA_signal_2989) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_2990), .Q (new_AGEMA_signal_2991) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_2992), .Q (new_AGEMA_signal_2993) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_2994), .Q (new_AGEMA_signal_2995) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_2996), .Q (new_AGEMA_signal_2997) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_2998), .Q (new_AGEMA_signal_2999) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_3000), .Q (new_AGEMA_signal_3001) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_3002), .Q (new_AGEMA_signal_3003) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_3004), .Q (new_AGEMA_signal_3005) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_3006), .Q (new_AGEMA_signal_3007) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_3008), .Q (new_AGEMA_signal_3009) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_3010), .Q (new_AGEMA_signal_3011) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_3012), .Q (new_AGEMA_signal_3013) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_3014), .Q (new_AGEMA_signal_3015) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_3016), .Q (new_AGEMA_signal_3017) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_3018), .Q (new_AGEMA_signal_3019) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_3020), .Q (new_AGEMA_signal_3021) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_3022), .Q (new_AGEMA_signal_3023) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_3030), .Q (new_AGEMA_signal_3031) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_3032), .Q (new_AGEMA_signal_3033) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_3034), .Q (new_AGEMA_signal_3035) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_3036), .Q (new_AGEMA_signal_3037) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_3038), .Q (new_AGEMA_signal_3039) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_3040), .Q (new_AGEMA_signal_3041) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_3042), .Q (new_AGEMA_signal_3043) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_3044), .Q (new_AGEMA_signal_3045) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_3046), .Q (new_AGEMA_signal_3047) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_3048), .Q (new_AGEMA_signal_3049) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_3050), .Q (new_AGEMA_signal_3051) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_3052), .Q (new_AGEMA_signal_3053) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_3054), .Q (new_AGEMA_signal_3055) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_3056), .Q (new_AGEMA_signal_3057) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_3058), .Q (new_AGEMA_signal_3059) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_3060), .Q (new_AGEMA_signal_3061) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_3062), .Q (new_AGEMA_signal_3063) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_3064), .Q (new_AGEMA_signal_3065) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (clk), .D (new_AGEMA_signal_3066), .Q (new_AGEMA_signal_3067) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (clk), .D (new_AGEMA_signal_3068), .Q (new_AGEMA_signal_3069) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (clk), .D (new_AGEMA_signal_3070), .Q (new_AGEMA_signal_3071) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (clk), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_3073) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (clk), .D (new_AGEMA_signal_3074), .Q (new_AGEMA_signal_3075) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (clk), .D (new_AGEMA_signal_3076), .Q (new_AGEMA_signal_3077) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (clk), .D (new_AGEMA_signal_3078), .Q (new_AGEMA_signal_3079) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (clk), .D (new_AGEMA_signal_3080), .Q (new_AGEMA_signal_3081) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (clk), .D (new_AGEMA_signal_3082), .Q (new_AGEMA_signal_3083) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (clk), .D (new_AGEMA_signal_3084), .Q (new_AGEMA_signal_3085) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (clk), .D (new_AGEMA_signal_3086), .Q (new_AGEMA_signal_3087) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (clk), .D (new_AGEMA_signal_3088), .Q (new_AGEMA_signal_3089) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (clk), .D (new_AGEMA_signal_3090), .Q (new_AGEMA_signal_3091) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (clk), .D (new_AGEMA_signal_3092), .Q (new_AGEMA_signal_3093) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (clk), .D (new_AGEMA_signal_3094), .Q (new_AGEMA_signal_3095) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C (clk), .D (new_AGEMA_signal_4713), .Q (new_AGEMA_signal_4714) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C (clk), .D (new_AGEMA_signal_4721), .Q (new_AGEMA_signal_4722) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C (clk), .D (new_AGEMA_signal_4729), .Q (new_AGEMA_signal_4730) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C (clk), .D (new_AGEMA_signal_4737), .Q (new_AGEMA_signal_4738) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C (clk), .D (new_AGEMA_signal_4745), .Q (new_AGEMA_signal_4746) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C (clk), .D (new_AGEMA_signal_4753), .Q (new_AGEMA_signal_4754) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C (clk), .D (new_AGEMA_signal_4761), .Q (new_AGEMA_signal_4762) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C (clk), .D (new_AGEMA_signal_4769), .Q (new_AGEMA_signal_4770) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C (clk), .D (new_AGEMA_signal_4777), .Q (new_AGEMA_signal_4778) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C (clk), .D (new_AGEMA_signal_4785), .Q (new_AGEMA_signal_4786) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C (clk), .D (new_AGEMA_signal_4793), .Q (new_AGEMA_signal_4794) ) ;
    buf_clk new_AGEMA_reg_buffer_3097 ( .C (clk), .D (new_AGEMA_signal_4801), .Q (new_AGEMA_signal_4802) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C (clk), .D (new_AGEMA_signal_4809), .Q (new_AGEMA_signal_4810) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C (clk), .D (new_AGEMA_signal_4817), .Q (new_AGEMA_signal_4818) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C (clk), .D (new_AGEMA_signal_4825), .Q (new_AGEMA_signal_4826) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C (clk), .D (new_AGEMA_signal_4833), .Q (new_AGEMA_signal_4834) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C (clk), .D (new_AGEMA_signal_4841), .Q (new_AGEMA_signal_4842) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C (clk), .D (new_AGEMA_signal_4849), .Q (new_AGEMA_signal_4850) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C (clk), .D (new_AGEMA_signal_4857), .Q (new_AGEMA_signal_4858) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C (clk), .D (new_AGEMA_signal_4865), .Q (new_AGEMA_signal_4866) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C (clk), .D (new_AGEMA_signal_4873), .Q (new_AGEMA_signal_4874) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C (clk), .D (new_AGEMA_signal_4881), .Q (new_AGEMA_signal_4882) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C (clk), .D (new_AGEMA_signal_4889), .Q (new_AGEMA_signal_4890) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C (clk), .D (new_AGEMA_signal_4897), .Q (new_AGEMA_signal_4898) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C (clk), .D (new_AGEMA_signal_4905), .Q (new_AGEMA_signal_4906) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C (clk), .D (new_AGEMA_signal_4913), .Q (new_AGEMA_signal_4914) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C (clk), .D (new_AGEMA_signal_4921), .Q (new_AGEMA_signal_4922) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C (clk), .D (new_AGEMA_signal_4929), .Q (new_AGEMA_signal_4930) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C (clk), .D (new_AGEMA_signal_4937), .Q (new_AGEMA_signal_4938) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C (clk), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_4946) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C (clk), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_4954) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C (clk), .D (new_AGEMA_signal_4961), .Q (new_AGEMA_signal_4962) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C (clk), .D (new_AGEMA_signal_4969), .Q (new_AGEMA_signal_4970) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C (clk), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_4978) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C (clk), .D (new_AGEMA_signal_4985), .Q (new_AGEMA_signal_4986) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_4994) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C (clk), .D (new_AGEMA_signal_5001), .Q (new_AGEMA_signal_5002) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C (clk), .D (new_AGEMA_signal_5009), .Q (new_AGEMA_signal_5010) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C (clk), .D (new_AGEMA_signal_5017), .Q (new_AGEMA_signal_5018) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C (clk), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_5026) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C (clk), .D (new_AGEMA_signal_5033), .Q (new_AGEMA_signal_5034) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C (clk), .D (new_AGEMA_signal_5041), .Q (new_AGEMA_signal_5042) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C (clk), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_5050) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C (clk), .D (new_AGEMA_signal_5057), .Q (new_AGEMA_signal_5058) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_5066) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C (clk), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_5074) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C (clk), .D (new_AGEMA_signal_5081), .Q (new_AGEMA_signal_5082) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C (clk), .D (new_AGEMA_signal_5089), .Q (new_AGEMA_signal_5090) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C (clk), .D (new_AGEMA_signal_5097), .Q (new_AGEMA_signal_5098) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C (clk), .D (new_AGEMA_signal_5105), .Q (new_AGEMA_signal_5106) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_5114) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C (clk), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_5122) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C (clk), .D (new_AGEMA_signal_5129), .Q (new_AGEMA_signal_5130) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_5138) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_5146) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C (clk), .D (new_AGEMA_signal_5153), .Q (new_AGEMA_signal_5154) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C (clk), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_5162) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C (clk), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_5170) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C (clk), .D (new_AGEMA_signal_5177), .Q (new_AGEMA_signal_5178) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C (clk), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_5186) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_5194) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C (clk), .D (new_AGEMA_signal_5201), .Q (new_AGEMA_signal_5202) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_5210) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C (clk), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_5218) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C (clk), .D (new_AGEMA_signal_5225), .Q (new_AGEMA_signal_5226) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C (clk), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_5234) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C (clk), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_5242) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C (clk), .D (new_AGEMA_signal_5249), .Q (new_AGEMA_signal_5250) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C (clk), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_5258) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_5266) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C (clk), .D (new_AGEMA_signal_5273), .Q (new_AGEMA_signal_5274) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_5282) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C (clk), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_5290) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C (clk), .D (new_AGEMA_signal_5297), .Q (new_AGEMA_signal_5298) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C (clk), .D (new_AGEMA_signal_5305), .Q (new_AGEMA_signal_5306) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C (clk), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_5314) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C (clk), .D (new_AGEMA_signal_5321), .Q (new_AGEMA_signal_5322) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C (clk), .D (new_AGEMA_signal_5329), .Q (new_AGEMA_signal_5330) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_5338) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C (clk), .D (new_AGEMA_signal_5345), .Q (new_AGEMA_signal_5346) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C (clk), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_5354) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_5362) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C (clk), .D (new_AGEMA_signal_5369), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C (clk), .D (new_AGEMA_signal_5377), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C (clk), .D (new_AGEMA_signal_5385), .Q (new_AGEMA_signal_5386) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C (clk), .D (new_AGEMA_signal_5393), .Q (new_AGEMA_signal_5394) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C (clk), .D (new_AGEMA_signal_5401), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C (clk), .D (new_AGEMA_signal_5409), .Q (new_AGEMA_signal_5410) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C (clk), .D (new_AGEMA_signal_5417), .Q (new_AGEMA_signal_5418) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C (clk), .D (new_AGEMA_signal_5425), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C (clk), .D (new_AGEMA_signal_5433), .Q (new_AGEMA_signal_5434) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C (clk), .D (new_AGEMA_signal_5441), .Q (new_AGEMA_signal_5442) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C (clk), .D (new_AGEMA_signal_5449), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C (clk), .D (new_AGEMA_signal_5457), .Q (new_AGEMA_signal_5458) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C (clk), .D (new_AGEMA_signal_5465), .Q (new_AGEMA_signal_5466) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C (clk), .D (new_AGEMA_signal_5473), .Q (new_AGEMA_signal_5474) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C (clk), .D (new_AGEMA_signal_5481), .Q (new_AGEMA_signal_5482) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C (clk), .D (new_AGEMA_signal_5489), .Q (new_AGEMA_signal_5490) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C (clk), .D (new_AGEMA_signal_5497), .Q (new_AGEMA_signal_5498) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C (clk), .D (new_AGEMA_signal_5505), .Q (new_AGEMA_signal_5506) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C (clk), .D (new_AGEMA_signal_5513), .Q (new_AGEMA_signal_5514) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C (clk), .D (new_AGEMA_signal_5521), .Q (new_AGEMA_signal_5522) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C (clk), .D (new_AGEMA_signal_5529), .Q (new_AGEMA_signal_5530) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C (clk), .D (new_AGEMA_signal_5537), .Q (new_AGEMA_signal_5538) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C (clk), .D (new_AGEMA_signal_5545), .Q (new_AGEMA_signal_5546) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C (clk), .D (new_AGEMA_signal_5553), .Q (new_AGEMA_signal_5554) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C (clk), .D (new_AGEMA_signal_5561), .Q (new_AGEMA_signal_5562) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C (clk), .D (new_AGEMA_signal_5569), .Q (new_AGEMA_signal_5570) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C (clk), .D (new_AGEMA_signal_5577), .Q (new_AGEMA_signal_5578) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C (clk), .D (new_AGEMA_signal_5585), .Q (new_AGEMA_signal_5586) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C (clk), .D (new_AGEMA_signal_5593), .Q (new_AGEMA_signal_5594) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C (clk), .D (new_AGEMA_signal_5601), .Q (new_AGEMA_signal_5602) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C (clk), .D (new_AGEMA_signal_5609), .Q (new_AGEMA_signal_5610) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C (clk), .D (new_AGEMA_signal_5617), .Q (new_AGEMA_signal_5618) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C (clk), .D (new_AGEMA_signal_5625), .Q (new_AGEMA_signal_5626) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C (clk), .D (new_AGEMA_signal_5633), .Q (new_AGEMA_signal_5634) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C (clk), .D (new_AGEMA_signal_5641), .Q (new_AGEMA_signal_5642) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C (clk), .D (new_AGEMA_signal_5649), .Q (new_AGEMA_signal_5650) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C (clk), .D (new_AGEMA_signal_5657), .Q (new_AGEMA_signal_5658) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C (clk), .D (new_AGEMA_signal_5665), .Q (new_AGEMA_signal_5666) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C (clk), .D (new_AGEMA_signal_5673), .Q (new_AGEMA_signal_5674) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C (clk), .D (new_AGEMA_signal_5681), .Q (new_AGEMA_signal_5682) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C (clk), .D (new_AGEMA_signal_5689), .Q (new_AGEMA_signal_5690) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C (clk), .D (new_AGEMA_signal_5697), .Q (new_AGEMA_signal_5698) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C (clk), .D (new_AGEMA_signal_5705), .Q (new_AGEMA_signal_5706) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C (clk), .D (new_AGEMA_signal_5713), .Q (new_AGEMA_signal_5714) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C (clk), .D (new_AGEMA_signal_5721), .Q (new_AGEMA_signal_5722) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C (clk), .D (new_AGEMA_signal_5729), .Q (new_AGEMA_signal_5730) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_4125), .Q (new_AGEMA_signal_5732) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_5740) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_5747), .Q (new_AGEMA_signal_5748) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_5756) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_5772) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_5796) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_5804) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_5844) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_5852) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_5868) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_5876) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_5916) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_5924) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_5964) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_5972) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_6012) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_6020) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_6036) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_6044) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_6084) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_6092) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_6132) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_6139), .Q (new_AGEMA_signal_6140) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_6180) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_6188) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_6204) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_6212) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_6438) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C (clk), .D (new_AGEMA_signal_6445), .Q (new_AGEMA_signal_6446) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C (clk), .D (new_AGEMA_signal_6453), .Q (new_AGEMA_signal_6454) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C (clk), .D (new_AGEMA_signal_6461), .Q (new_AGEMA_signal_6462) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C (clk), .D (new_AGEMA_signal_6469), .Q (new_AGEMA_signal_6470) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_1_DQ), .Q (new_AGEMA_signal_6472) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C (clk), .D (new_AGEMA_signal_2565), .Q (new_AGEMA_signal_6474) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_3_DQ), .Q (new_AGEMA_signal_6476) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C (clk), .D (new_AGEMA_signal_2567), .Q (new_AGEMA_signal_6478) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_5_DQ), .Q (new_AGEMA_signal_6480) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C (clk), .D (new_AGEMA_signal_2568), .Q (new_AGEMA_signal_6482) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_7_DQ), .Q (new_AGEMA_signal_6484) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C (clk), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_6486) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_9_DQ), .Q (new_AGEMA_signal_6488) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C (clk), .D (new_AGEMA_signal_2571), .Q (new_AGEMA_signal_6490) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_11_DQ), .Q (new_AGEMA_signal_6492) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C (clk), .D (new_AGEMA_signal_2573), .Q (new_AGEMA_signal_6494) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_13_DQ), .Q (new_AGEMA_signal_6496) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C (clk), .D (new_AGEMA_signal_2574), .Q (new_AGEMA_signal_6498) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_15_DQ), .Q (new_AGEMA_signal_6500) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C (clk), .D (new_AGEMA_signal_2576), .Q (new_AGEMA_signal_6502) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_17_DQ), .Q (new_AGEMA_signal_6504) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C (clk), .D (new_AGEMA_signal_2577), .Q (new_AGEMA_signal_6506) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_19_DQ), .Q (new_AGEMA_signal_6508) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C (clk), .D (new_AGEMA_signal_2579), .Q (new_AGEMA_signal_6510) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_21_DQ), .Q (new_AGEMA_signal_6512) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C (clk), .D (new_AGEMA_signal_2580), .Q (new_AGEMA_signal_6514) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_23_DQ), .Q (new_AGEMA_signal_6516) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C (clk), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_6518) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_25_DQ), .Q (new_AGEMA_signal_6520) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C (clk), .D (new_AGEMA_signal_2583), .Q (new_AGEMA_signal_6522) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_27_DQ), .Q (new_AGEMA_signal_6524) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_6526) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_29_DQ), .Q (new_AGEMA_signal_6528) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C (clk), .D (new_AGEMA_signal_2586), .Q (new_AGEMA_signal_6530) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_31_DQ), .Q (new_AGEMA_signal_6532) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_6534) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_33_DQ), .Q (new_AGEMA_signal_6536) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C (clk), .D (new_AGEMA_signal_2589), .Q (new_AGEMA_signal_6538) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_35_DQ), .Q (new_AGEMA_signal_6540) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C (clk), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_6542) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_37_DQ), .Q (new_AGEMA_signal_6544) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C (clk), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_6546) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_39_DQ), .Q (new_AGEMA_signal_6548) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C (clk), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_6550) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_41_DQ), .Q (new_AGEMA_signal_6552) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C (clk), .D (new_AGEMA_signal_2595), .Q (new_AGEMA_signal_6554) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_43_DQ), .Q (new_AGEMA_signal_6556) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C (clk), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_6558) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_45_DQ), .Q (new_AGEMA_signal_6560) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C (clk), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_6562) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_47_DQ), .Q (new_AGEMA_signal_6564) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C (clk), .D (new_AGEMA_signal_2600), .Q (new_AGEMA_signal_6566) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_49_DQ), .Q (new_AGEMA_signal_6568) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C (clk), .D (new_AGEMA_signal_2601), .Q (new_AGEMA_signal_6570) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_51_DQ), .Q (new_AGEMA_signal_6572) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_6574) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_53_DQ), .Q (new_AGEMA_signal_6576) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C (clk), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_6578) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_55_DQ), .Q (new_AGEMA_signal_6580) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_6582) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_57_DQ), .Q (new_AGEMA_signal_6584) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C (clk), .D (new_AGEMA_signal_2607), .Q (new_AGEMA_signal_6586) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_59_DQ), .Q (new_AGEMA_signal_6588) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C (clk), .D (new_AGEMA_signal_2609), .Q (new_AGEMA_signal_6590) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_61_DQ), .Q (new_AGEMA_signal_6592) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C (clk), .D (new_AGEMA_signal_2610), .Q (new_AGEMA_signal_6594) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C (clk), .D (Midori_rounds_roundResult_Reg_SFF_63_DQ), .Q (new_AGEMA_signal_6596) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_6598) ) ;

    /* cells in depth 8 */
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U127 ( .a ({new_AGEMA_signal_4723, new_AGEMA_signal_4715}), .b ({new_AGEMA_signal_2155, Midori_rounds_SR_Result[8]}), .c ({DataOut_s1[8], DataOut_s0[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U125 ( .a ({new_AGEMA_signal_4739, new_AGEMA_signal_4731}), .b ({new_AGEMA_signal_2149, Midori_rounds_SR_Result[46]}), .c ({DataOut_s1[6], DataOut_s0[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U123 ( .a ({new_AGEMA_signal_4755, new_AGEMA_signal_4747}), .b ({new_AGEMA_signal_2205, Midori_rounds_SR_Result[62]}), .c ({DataOut_s1[62], DataOut_s0[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U121 ( .a ({new_AGEMA_signal_4771, new_AGEMA_signal_4763}), .b ({new_AGEMA_signal_2207, Midori_rounds_SR_Result[60]}), .c ({DataOut_s1[60], DataOut_s0[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U118 ( .a ({new_AGEMA_signal_4787, new_AGEMA_signal_4779}), .b ({new_AGEMA_signal_2201, Midori_rounds_SR_Result[34]}), .c ({DataOut_s1[58], DataOut_s0[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U116 ( .a ({new_AGEMA_signal_4803, new_AGEMA_signal_4795}), .b ({new_AGEMA_signal_2203, Midori_rounds_SR_Result[32]}), .c ({DataOut_s1[56], DataOut_s0[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U114 ( .a ({new_AGEMA_signal_4819, new_AGEMA_signal_4811}), .b ({new_AGEMA_signal_2197, Midori_rounds_SR_Result[6]}), .c ({DataOut_s1[54], DataOut_s0[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U112 ( .a ({new_AGEMA_signal_4835, new_AGEMA_signal_4827}), .b ({new_AGEMA_signal_2199, Midori_rounds_SR_Result[4]}), .c ({DataOut_s1[52], DataOut_s0[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U110 ( .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4843}), .b ({new_AGEMA_signal_2193, Midori_rounds_SR_Result[26]}), .c ({DataOut_s1[50], DataOut_s0[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U109 ( .a ({new_AGEMA_signal_4867, new_AGEMA_signal_4859}), .b ({new_AGEMA_signal_2151, Midori_rounds_SR_Result[44]}), .c ({DataOut_s1[4], DataOut_s0[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U107 ( .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4875}), .b ({new_AGEMA_signal_2195, Midori_rounds_SR_Result[24]}), .c ({DataOut_s1[48], DataOut_s0[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U105 ( .a ({new_AGEMA_signal_4899, new_AGEMA_signal_4891}), .b ({new_AGEMA_signal_2189, Midori_rounds_SR_Result[42]}), .c ({DataOut_s1[46], DataOut_s0[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U103 ( .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4907}), .b ({new_AGEMA_signal_2191, Midori_rounds_SR_Result[40]}), .c ({DataOut_s1[44], DataOut_s0[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U101 ( .a ({new_AGEMA_signal_4931, new_AGEMA_signal_4923}), .b ({new_AGEMA_signal_2185, Midori_rounds_SR_Result[54]}), .c ({DataOut_s1[42], DataOut_s0[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U99 ( .a ({new_AGEMA_signal_4947, new_AGEMA_signal_4939}), .b ({new_AGEMA_signal_2187, Midori_rounds_SR_Result[52]}), .c ({DataOut_s1[40], DataOut_s0[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U96 ( .a ({new_AGEMA_signal_4963, new_AGEMA_signal_4955}), .b ({new_AGEMA_signal_2181, Midori_rounds_SR_Result[18]}), .c ({DataOut_s1[38], DataOut_s0[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U94 ( .a ({new_AGEMA_signal_4979, new_AGEMA_signal_4971}), .b ({new_AGEMA_signal_2183, Midori_rounds_SR_Result[16]}), .c ({DataOut_s1[36], DataOut_s0[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U92 ( .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4987}), .b ({new_AGEMA_signal_2177, Midori_rounds_SR_Result[14]}), .c ({DataOut_s1[34], DataOut_s0[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U90 ( .a ({new_AGEMA_signal_5011, new_AGEMA_signal_5003}), .b ({new_AGEMA_signal_2179, Midori_rounds_SR_Result[12]}), .c ({DataOut_s1[32], DataOut_s0[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U88 ( .a ({new_AGEMA_signal_5027, new_AGEMA_signal_5019}), .b ({new_AGEMA_signal_2173, Midori_rounds_SR_Result[2]}), .c ({DataOut_s1[30], DataOut_s0[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U87 ( .a ({new_AGEMA_signal_5043, new_AGEMA_signal_5035}), .b ({new_AGEMA_signal_2145, Midori_rounds_SR_Result[50]}), .c ({DataOut_s1[2], DataOut_s0[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U85 ( .a ({new_AGEMA_signal_5059, new_AGEMA_signal_5051}), .b ({new_AGEMA_signal_2175, Midori_rounds_SR_Result[0]}), .c ({DataOut_s1[28], DataOut_s0[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U83 ( .a ({new_AGEMA_signal_5075, new_AGEMA_signal_5067}), .b ({new_AGEMA_signal_2169, Midori_rounds_SR_Result[30]}), .c ({DataOut_s1[26], DataOut_s0[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U81 ( .a ({new_AGEMA_signal_5091, new_AGEMA_signal_5083}), .b ({new_AGEMA_signal_2171, Midori_rounds_SR_Result[28]}), .c ({DataOut_s1[24], DataOut_s0[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U79 ( .a ({new_AGEMA_signal_5107, new_AGEMA_signal_5099}), .b ({new_AGEMA_signal_2165, Midori_rounds_SR_Result[58]}), .c ({DataOut_s1[22], DataOut_s0[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U77 ( .a ({new_AGEMA_signal_5123, new_AGEMA_signal_5115}), .b ({new_AGEMA_signal_2167, Midori_rounds_SR_Result[56]}), .c ({DataOut_s1[20], DataOut_s0[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U74 ( .a ({new_AGEMA_signal_5139, new_AGEMA_signal_5131}), .b ({new_AGEMA_signal_2161, Midori_rounds_SR_Result[38]}), .c ({DataOut_s1[18], DataOut_s0[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U72 ( .a ({new_AGEMA_signal_5155, new_AGEMA_signal_5147}), .b ({new_AGEMA_signal_2163, Midori_rounds_SR_Result[36]}), .c ({DataOut_s1[16], DataOut_s0[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U70 ( .a ({new_AGEMA_signal_5171, new_AGEMA_signal_5163}), .b ({new_AGEMA_signal_2157, Midori_rounds_SR_Result[22]}), .c ({DataOut_s1[14], DataOut_s0[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U68 ( .a ({new_AGEMA_signal_5187, new_AGEMA_signal_5179}), .b ({new_AGEMA_signal_2159, Midori_rounds_SR_Result[20]}), .c ({DataOut_s1[12], DataOut_s0[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U66 ( .a ({new_AGEMA_signal_5203, new_AGEMA_signal_5195}), .b ({new_AGEMA_signal_2153, Midori_rounds_SR_Result[10]}), .c ({DataOut_s1[10], DataOut_s0[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_U65 ( .a ({new_AGEMA_signal_5219, new_AGEMA_signal_5211}), .b ({new_AGEMA_signal_2147, Midori_rounds_SR_Result[48]}), .c ({DataOut_s1[0], DataOut_s0[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U143 ( .a ({new_AGEMA_signal_2155, Midori_rounds_SR_Result[8]}), .b ({new_AGEMA_signal_5235, new_AGEMA_signal_5227}), .c ({new_AGEMA_signal_2492, Midori_rounds_sub_ResultXORkey[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U141 ( .a ({new_AGEMA_signal_5251, new_AGEMA_signal_5243}), .b ({new_AGEMA_signal_2149, Midori_rounds_SR_Result[46]}), .c ({new_AGEMA_signal_2274, Midori_rounds_sub_ResultXORkey[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U139 ( .a ({new_AGEMA_signal_5267, new_AGEMA_signal_5259}), .b ({new_AGEMA_signal_2205, Midori_rounds_SR_Result[62]}), .c ({new_AGEMA_signal_2276, Midori_rounds_sub_ResultXORkey[62]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U137 ( .a ({new_AGEMA_signal_2207, Midori_rounds_SR_Result[60]}), .b ({new_AGEMA_signal_5283, new_AGEMA_signal_5275}), .c ({new_AGEMA_signal_2554, Midori_rounds_sub_ResultXORkey[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U134 ( .a ({new_AGEMA_signal_5299, new_AGEMA_signal_5291}), .b ({new_AGEMA_signal_2201, Midori_rounds_SR_Result[34]}), .c ({new_AGEMA_signal_2280, Midori_rounds_sub_ResultXORkey[58]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U132 ( .a ({new_AGEMA_signal_2203, Midori_rounds_SR_Result[32]}), .b ({new_AGEMA_signal_5315, new_AGEMA_signal_5307}), .c ({new_AGEMA_signal_2555, Midori_rounds_sub_ResultXORkey[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U130 ( .a ({new_AGEMA_signal_5331, new_AGEMA_signal_5323}), .b ({new_AGEMA_signal_2197, Midori_rounds_SR_Result[6]}), .c ({new_AGEMA_signal_2283, Midori_rounds_sub_ResultXORkey[54]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U128 ( .a ({new_AGEMA_signal_2199, Midori_rounds_SR_Result[4]}), .b ({new_AGEMA_signal_5347, new_AGEMA_signal_5339}), .c ({new_AGEMA_signal_2556, Midori_rounds_sub_ResultXORkey[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U126 ( .a ({new_AGEMA_signal_5363, new_AGEMA_signal_5355}), .b ({new_AGEMA_signal_2193, Midori_rounds_SR_Result[26]}), .c ({new_AGEMA_signal_2286, Midori_rounds_sub_ResultXORkey[50]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U125 ( .a ({new_AGEMA_signal_2151, Midori_rounds_SR_Result[44]}), .b ({new_AGEMA_signal_5379, new_AGEMA_signal_5371}), .c ({new_AGEMA_signal_2557, Midori_rounds_sub_ResultXORkey[4]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U123 ( .a ({new_AGEMA_signal_2195, Midori_rounds_SR_Result[24]}), .b ({new_AGEMA_signal_5395, new_AGEMA_signal_5387}), .c ({new_AGEMA_signal_2629, Midori_rounds_sub_ResultXORkey[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U121 ( .a ({new_AGEMA_signal_5411, new_AGEMA_signal_5403}), .b ({new_AGEMA_signal_2189, Midori_rounds_SR_Result[42]}), .c ({new_AGEMA_signal_2289, Midori_rounds_sub_ResultXORkey[46]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U119 ( .a ({new_AGEMA_signal_2191, Midori_rounds_SR_Result[40]}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5419}), .c ({new_AGEMA_signal_2493, Midori_rounds_sub_ResultXORkey[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U117 ( .a ({new_AGEMA_signal_5443, new_AGEMA_signal_5435}), .b ({new_AGEMA_signal_2185, Midori_rounds_SR_Result[54]}), .c ({new_AGEMA_signal_2292, Midori_rounds_sub_ResultXORkey[42]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U115 ( .a ({new_AGEMA_signal_2187, Midori_rounds_SR_Result[52]}), .b ({new_AGEMA_signal_5459, new_AGEMA_signal_5451}), .c ({new_AGEMA_signal_2558, Midori_rounds_sub_ResultXORkey[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U112 ( .a ({new_AGEMA_signal_5475, new_AGEMA_signal_5467}), .b ({new_AGEMA_signal_2181, Midori_rounds_SR_Result[18]}), .c ({new_AGEMA_signal_2296, Midori_rounds_sub_ResultXORkey[38]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U110 ( .a ({new_AGEMA_signal_2183, Midori_rounds_SR_Result[16]}), .b ({new_AGEMA_signal_5491, new_AGEMA_signal_5483}), .c ({new_AGEMA_signal_2494, Midori_rounds_sub_ResultXORkey[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U108 ( .a ({new_AGEMA_signal_5507, new_AGEMA_signal_5499}), .b ({new_AGEMA_signal_2177, Midori_rounds_SR_Result[14]}), .c ({new_AGEMA_signal_2299, Midori_rounds_sub_ResultXORkey[34]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U106 ( .a ({new_AGEMA_signal_2179, Midori_rounds_SR_Result[12]}), .b ({new_AGEMA_signal_5523, new_AGEMA_signal_5515}), .c ({new_AGEMA_signal_2559, Midori_rounds_sub_ResultXORkey[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U104 ( .a ({new_AGEMA_signal_5539, new_AGEMA_signal_5531}), .b ({new_AGEMA_signal_2173, Midori_rounds_SR_Result[2]}), .c ({new_AGEMA_signal_2302, Midori_rounds_sub_ResultXORkey[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U103 ( .a ({new_AGEMA_signal_5555, new_AGEMA_signal_5547}), .b ({new_AGEMA_signal_2145, Midori_rounds_SR_Result[50]}), .c ({new_AGEMA_signal_2303, Midori_rounds_sub_ResultXORkey[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U101 ( .a ({new_AGEMA_signal_2175, Midori_rounds_SR_Result[0]}), .b ({new_AGEMA_signal_5571, new_AGEMA_signal_5563}), .c ({new_AGEMA_signal_2617, Midori_rounds_sub_ResultXORkey[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U99 ( .a ({new_AGEMA_signal_5587, new_AGEMA_signal_5579}), .b ({new_AGEMA_signal_2169, Midori_rounds_SR_Result[30]}), .c ({new_AGEMA_signal_2306, Midori_rounds_sub_ResultXORkey[26]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U97 ( .a ({new_AGEMA_signal_2171, Midori_rounds_SR_Result[28]}), .b ({new_AGEMA_signal_5603, new_AGEMA_signal_5595}), .c ({new_AGEMA_signal_2560, Midori_rounds_sub_ResultXORkey[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U95 ( .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5611}), .b ({new_AGEMA_signal_2165, Midori_rounds_SR_Result[58]}), .c ({new_AGEMA_signal_2309, Midori_rounds_sub_ResultXORkey[22]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U93 ( .a ({new_AGEMA_signal_2167, Midori_rounds_SR_Result[56]}), .b ({new_AGEMA_signal_5635, new_AGEMA_signal_5627}), .c ({new_AGEMA_signal_2495, Midori_rounds_sub_ResultXORkey[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U90 ( .a ({new_AGEMA_signal_5651, new_AGEMA_signal_5643}), .b ({new_AGEMA_signal_2161, Midori_rounds_SR_Result[38]}), .c ({new_AGEMA_signal_2313, Midori_rounds_sub_ResultXORkey[18]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U88 ( .a ({new_AGEMA_signal_2163, Midori_rounds_SR_Result[36]}), .b ({new_AGEMA_signal_5667, new_AGEMA_signal_5659}), .c ({new_AGEMA_signal_2561, Midori_rounds_sub_ResultXORkey[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U86 ( .a ({new_AGEMA_signal_5683, new_AGEMA_signal_5675}), .b ({new_AGEMA_signal_2157, Midori_rounds_SR_Result[22]}), .c ({new_AGEMA_signal_2316, Midori_rounds_sub_ResultXORkey[14]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U84 ( .a ({new_AGEMA_signal_2159, Midori_rounds_SR_Result[20]}), .b ({new_AGEMA_signal_5699, new_AGEMA_signal_5691}), .c ({new_AGEMA_signal_2562, Midori_rounds_sub_ResultXORkey[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U82 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5707}), .b ({new_AGEMA_signal_2153, Midori_rounds_SR_Result[10]}), .c ({new_AGEMA_signal_2319, Midori_rounds_sub_ResultXORkey[10]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U81 ( .a ({new_AGEMA_signal_2147, Midori_rounds_SR_Result[48]}), .b ({new_AGEMA_signal_5731, new_AGEMA_signal_5723}), .c ({new_AGEMA_signal_2563, Midori_rounds_sub_ResultXORkey[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U79 ( .a ({new_AGEMA_signal_2646, Midori_rounds_SR_Inv_Result[8]}), .b ({new_AGEMA_signal_5235, new_AGEMA_signal_5227}), .c ({new_AGEMA_signal_2650, Midori_rounds_mul_ResultXORkey[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U76 ( .a ({new_AGEMA_signal_5251, new_AGEMA_signal_5243}), .b ({new_AGEMA_signal_2430, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_2443, Midori_rounds_mul_ResultXORkey[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U74 ( .a ({new_AGEMA_signal_5267, new_AGEMA_signal_5259}), .b ({new_AGEMA_signal_2400, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_2445, Midori_rounds_mul_ResultXORkey[62]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U72 ( .a ({new_AGEMA_signal_2669, Midori_rounds_SR_Inv_Result[60]}), .b ({new_AGEMA_signal_5283, new_AGEMA_signal_5275}), .c ({new_AGEMA_signal_2681, Midori_rounds_mul_ResultXORkey[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U68 ( .a ({new_AGEMA_signal_5299, new_AGEMA_signal_5291}), .b ({new_AGEMA_signal_2403, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_2449, Midori_rounds_mul_ResultXORkey[58]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U66 ( .a ({new_AGEMA_signal_2668, Midori_rounds_SR_Inv_Result[20]}), .b ({new_AGEMA_signal_5315, new_AGEMA_signal_5307}), .c ({new_AGEMA_signal_2682, Midori_rounds_mul_ResultXORkey[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U63 ( .a ({new_AGEMA_signal_5331, new_AGEMA_signal_5323}), .b ({new_AGEMA_signal_2394, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_2452, Midori_rounds_mul_ResultXORkey[54]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U61 ( .a ({new_AGEMA_signal_2661, Midori_rounds_SR_Inv_Result[40]}), .b ({new_AGEMA_signal_5347, new_AGEMA_signal_5339}), .c ({new_AGEMA_signal_2665, Midori_rounds_mul_ResultXORkey[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U58 ( .a ({new_AGEMA_signal_5363, new_AGEMA_signal_5355}), .b ({new_AGEMA_signal_2397, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_2455, Midori_rounds_mul_ResultXORkey[50]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U57 ( .a ({new_AGEMA_signal_2647, Midori_rounds_SR_Inv_Result[52]}), .b ({new_AGEMA_signal_5379, new_AGEMA_signal_5371}), .c ({new_AGEMA_signal_2651, Midori_rounds_mul_ResultXORkey[4]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U54 ( .a ({new_AGEMA_signal_2638, Midori_rounds_SR_Inv_Result[0]}), .b ({new_AGEMA_signal_5395, new_AGEMA_signal_5387}), .c ({new_AGEMA_signal_2652, Midori_rounds_mul_ResultXORkey[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U51 ( .a ({new_AGEMA_signal_5411, new_AGEMA_signal_5403}), .b ({new_AGEMA_signal_2412, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_2458, Midori_rounds_mul_ResultXORkey[46]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U49 ( .a ({new_AGEMA_signal_2641, Midori_rounds_SR_Inv_Result[4]}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5419}), .c ({new_AGEMA_signal_2653, Midori_rounds_mul_ResultXORkey[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U46 ( .a ({new_AGEMA_signal_5443, new_AGEMA_signal_5435}), .b ({new_AGEMA_signal_2415, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_2462, Midori_rounds_mul_ResultXORkey[42]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U44 ( .a ({new_AGEMA_signal_2639, Midori_rounds_SR_Inv_Result[44]}), .b ({new_AGEMA_signal_5459, new_AGEMA_signal_5451}), .c ({new_AGEMA_signal_2654, Midori_rounds_mul_ResultXORkey[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U40 ( .a ({new_AGEMA_signal_5475, new_AGEMA_signal_5467}), .b ({new_AGEMA_signal_2406, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_2466, Midori_rounds_mul_ResultXORkey[38]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U38 ( .a ({new_AGEMA_signal_2640, Midori_rounds_SR_Inv_Result[16]}), .b ({new_AGEMA_signal_5491, new_AGEMA_signal_5483}), .c ({new_AGEMA_signal_2655, Midori_rounds_mul_ResultXORkey[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U35 ( .a ({new_AGEMA_signal_5507, new_AGEMA_signal_5499}), .b ({new_AGEMA_signal_2409, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_2470, Midori_rounds_mul_ResultXORkey[34]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U33 ( .a ({new_AGEMA_signal_2642, Midori_rounds_SR_Inv_Result[56]}), .b ({new_AGEMA_signal_5523, new_AGEMA_signal_5515}), .c ({new_AGEMA_signal_2656, Midori_rounds_mul_ResultXORkey[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U30 ( .a ({new_AGEMA_signal_5539, new_AGEMA_signal_5531}), .b ({new_AGEMA_signal_2424, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_2473, Midori_rounds_mul_ResultXORkey[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U29 ( .a ({new_AGEMA_signal_5555, new_AGEMA_signal_5547}), .b ({new_AGEMA_signal_2433, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_2474, Midori_rounds_mul_ResultXORkey[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U27 ( .a ({new_AGEMA_signal_2644, Midori_rounds_SR_Inv_Result[24]}), .b ({new_AGEMA_signal_5571, new_AGEMA_signal_5563}), .c ({new_AGEMA_signal_2657, Midori_rounds_mul_ResultXORkey[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U24 ( .a ({new_AGEMA_signal_5587, new_AGEMA_signal_5579}), .b ({new_AGEMA_signal_2427, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_2477, Midori_rounds_mul_ResultXORkey[26]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U22 ( .a ({new_AGEMA_signal_2643, Midori_rounds_SR_Inv_Result[48]}), .b ({new_AGEMA_signal_5603, new_AGEMA_signal_5595}), .c ({new_AGEMA_signal_2658, Midori_rounds_mul_ResultXORkey[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U19 ( .a ({new_AGEMA_signal_5619, new_AGEMA_signal_5611}), .b ({new_AGEMA_signal_2418, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_2480, Midori_rounds_mul_ResultXORkey[22]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U17 ( .a ({new_AGEMA_signal_2663, Midori_rounds_SR_Inv_Result[12]}), .b ({new_AGEMA_signal_5635, new_AGEMA_signal_5627}), .c ({new_AGEMA_signal_2666, Midori_rounds_mul_ResultXORkey[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U13 ( .a ({new_AGEMA_signal_5651, new_AGEMA_signal_5643}), .b ({new_AGEMA_signal_2421, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_2485, Midori_rounds_mul_ResultXORkey[18]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U11 ( .a ({new_AGEMA_signal_2664, Midori_rounds_SR_Inv_Result[36]}), .b ({new_AGEMA_signal_5667, new_AGEMA_signal_5659}), .c ({new_AGEMA_signal_2667, Midori_rounds_mul_ResultXORkey[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U8 ( .a ({new_AGEMA_signal_5683, new_AGEMA_signal_5675}), .b ({new_AGEMA_signal_2436, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_2488, Midori_rounds_mul_ResultXORkey[14]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U6 ( .a ({new_AGEMA_signal_2648, Midori_rounds_SR_Inv_Result[32]}), .b ({new_AGEMA_signal_5699, new_AGEMA_signal_5691}), .c ({new_AGEMA_signal_2659, Midori_rounds_mul_ResultXORkey[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U3 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5707}), .b ({new_AGEMA_signal_2439, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_2491, Midori_rounds_mul_ResultXORkey[10]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_U2 ( .a ({new_AGEMA_signal_2649, Midori_rounds_SR_Inv_Result[28]}), .b ({new_AGEMA_signal_5731, new_AGEMA_signal_5723}), .c ({new_AGEMA_signal_2660, Midori_rounds_mul_ResultXORkey[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2670, Midori_rounds_round_Result[0]}), .a ({new_AGEMA_signal_5749, new_AGEMA_signal_5741}), .c ({new_AGEMA_signal_2683, Midori_rounds_roundResult_Reg_SFF_0_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2507, Midori_rounds_round_Result[2]}), .a ({new_AGEMA_signal_5765, new_AGEMA_signal_5757}), .c ({new_AGEMA_signal_2566, Midori_rounds_roundResult_Reg_SFF_2_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2671, Midori_rounds_round_Result[4]}), .a ({new_AGEMA_signal_5781, new_AGEMA_signal_5773}), .c ({new_AGEMA_signal_2684, Midori_rounds_roundResult_Reg_SFF_4_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2510, Midori_rounds_round_Result[6]}), .a ({new_AGEMA_signal_5797, new_AGEMA_signal_5789}), .c ({new_AGEMA_signal_2569, Midori_rounds_roundResult_Reg_SFF_6_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2672, Midori_rounds_round_Result[8]}), .a ({new_AGEMA_signal_5813, new_AGEMA_signal_5805}), .c ({new_AGEMA_signal_2685, Midori_rounds_roundResult_Reg_SFF_8_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2513, Midori_rounds_round_Result[10]}), .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5821}), .c ({new_AGEMA_signal_2572, Midori_rounds_roundResult_Reg_SFF_10_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2673, Midori_rounds_round_Result[12]}), .a ({new_AGEMA_signal_5845, new_AGEMA_signal_5837}), .c ({new_AGEMA_signal_2686, Midori_rounds_roundResult_Reg_SFF_12_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2516, Midori_rounds_round_Result[14]}), .a ({new_AGEMA_signal_5861, new_AGEMA_signal_5853}), .c ({new_AGEMA_signal_2575, Midori_rounds_roundResult_Reg_SFF_14_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2694, Midori_rounds_round_Result[16]}), .a ({new_AGEMA_signal_5877, new_AGEMA_signal_5869}), .c ({new_AGEMA_signal_2697, Midori_rounds_roundResult_Reg_SFF_16_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2519, Midori_rounds_round_Result[18]}), .a ({new_AGEMA_signal_5893, new_AGEMA_signal_5885}), .c ({new_AGEMA_signal_2578, Midori_rounds_roundResult_Reg_SFF_18_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2695, Midori_rounds_round_Result[20]}), .a ({new_AGEMA_signal_5909, new_AGEMA_signal_5901}), .c ({new_AGEMA_signal_2698, Midori_rounds_roundResult_Reg_SFF_20_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2522, Midori_rounds_round_Result[22]}), .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5917}), .c ({new_AGEMA_signal_2581, Midori_rounds_roundResult_Reg_SFF_22_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2674, Midori_rounds_round_Result[24]}), .a ({new_AGEMA_signal_5941, new_AGEMA_signal_5933}), .c ({new_AGEMA_signal_2687, Midori_rounds_roundResult_Reg_SFF_24_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2525, Midori_rounds_round_Result[26]}), .a ({new_AGEMA_signal_5957, new_AGEMA_signal_5949}), .c ({new_AGEMA_signal_2584, Midori_rounds_roundResult_Reg_SFF_26_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2675, Midori_rounds_round_Result[28]}), .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5965}), .c ({new_AGEMA_signal_2688, Midori_rounds_roundResult_Reg_SFF_28_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2528, Midori_rounds_round_Result[30]}), .a ({new_AGEMA_signal_5989, new_AGEMA_signal_5981}), .c ({new_AGEMA_signal_2587, Midori_rounds_roundResult_Reg_SFF_30_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2676, Midori_rounds_round_Result[32]}), .a ({new_AGEMA_signal_6005, new_AGEMA_signal_5997}), .c ({new_AGEMA_signal_2689, Midori_rounds_roundResult_Reg_SFF_32_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2531, Midori_rounds_round_Result[34]}), .a ({new_AGEMA_signal_6021, new_AGEMA_signal_6013}), .c ({new_AGEMA_signal_2590, Midori_rounds_roundResult_Reg_SFF_34_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2677, Midori_rounds_round_Result[36]}), .a ({new_AGEMA_signal_6037, new_AGEMA_signal_6029}), .c ({new_AGEMA_signal_2690, Midori_rounds_roundResult_Reg_SFF_36_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2534, Midori_rounds_round_Result[38]}), .a ({new_AGEMA_signal_6053, new_AGEMA_signal_6045}), .c ({new_AGEMA_signal_2593, Midori_rounds_roundResult_Reg_SFF_38_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2678, Midori_rounds_round_Result[40]}), .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6061}), .c ({new_AGEMA_signal_2691, Midori_rounds_roundResult_Reg_SFF_40_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2537, Midori_rounds_round_Result[42]}), .a ({new_AGEMA_signal_6085, new_AGEMA_signal_6077}), .c ({new_AGEMA_signal_2596, Midori_rounds_roundResult_Reg_SFF_42_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2679, Midori_rounds_round_Result[44]}), .a ({new_AGEMA_signal_6101, new_AGEMA_signal_6093}), .c ({new_AGEMA_signal_2692, Midori_rounds_roundResult_Reg_SFF_44_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2540, Midori_rounds_round_Result[46]}), .a ({new_AGEMA_signal_6117, new_AGEMA_signal_6109}), .c ({new_AGEMA_signal_2599, Midori_rounds_roundResult_Reg_SFF_46_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2680, Midori_rounds_round_Result[48]}), .a ({new_AGEMA_signal_6133, new_AGEMA_signal_6125}), .c ({new_AGEMA_signal_2693, Midori_rounds_roundResult_Reg_SFF_48_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2543, Midori_rounds_round_Result[50]}), .a ({new_AGEMA_signal_6149, new_AGEMA_signal_6141}), .c ({new_AGEMA_signal_2602, Midori_rounds_roundResult_Reg_SFF_50_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2696, Midori_rounds_round_Result[52]}), .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6157}), .c ({new_AGEMA_signal_2699, Midori_rounds_roundResult_Reg_SFF_52_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2546, Midori_rounds_round_Result[54]}), .a ({new_AGEMA_signal_6181, new_AGEMA_signal_6173}), .c ({new_AGEMA_signal_2605, Midori_rounds_roundResult_Reg_SFF_54_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2700, Midori_rounds_round_Result[56]}), .a ({new_AGEMA_signal_6197, new_AGEMA_signal_6189}), .c ({new_AGEMA_signal_2702, Midori_rounds_roundResult_Reg_SFF_56_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2549, Midori_rounds_round_Result[58]}), .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6205}), .c ({new_AGEMA_signal_2608, Midori_rounds_roundResult_Reg_SFF_58_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2701, Midori_rounds_round_Result[60]}), .a ({new_AGEMA_signal_6229, new_AGEMA_signal_6221}), .c ({new_AGEMA_signal_2703, Midori_rounds_roundResult_Reg_SFF_60_DQ}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1 ( .s (new_AGEMA_signal_5733), .b ({new_AGEMA_signal_2552, Midori_rounds_round_Result[62]}), .a ({new_AGEMA_signal_6245, new_AGEMA_signal_6237}), .c ({new_AGEMA_signal_2611, Midori_rounds_roundResult_Reg_SFF_62_DQ}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6247}), .b ({new_AGEMA_signal_2066, Midori_rounds_sub_sBox_PRINCE_0_n12}), .clk (clk), .r (Fresh[224]), .c ({new_AGEMA_signal_2145, Midori_rounds_SR_Result[50]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .a ({new_AGEMA_signal_6257, new_AGEMA_signal_6253}), .b ({new_AGEMA_signal_2068, Midori_rounds_sub_sBox_PRINCE_0_n3}), .clk (clk), .r (Fresh[225]), .c ({new_AGEMA_signal_2147, Midori_rounds_SR_Result[48]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .a ({new_AGEMA_signal_6261, new_AGEMA_signal_6259}), .b ({new_AGEMA_signal_2071, Midori_rounds_sub_sBox_PRINCE_1_n12}), .clk (clk), .r (Fresh[226]), .c ({new_AGEMA_signal_2149, Midori_rounds_SR_Result[46]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .a ({new_AGEMA_signal_6269, new_AGEMA_signal_6265}), .b ({new_AGEMA_signal_2073, Midori_rounds_sub_sBox_PRINCE_1_n3}), .clk (clk), .r (Fresh[227]), .c ({new_AGEMA_signal_2151, Midori_rounds_SR_Result[44]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6271}), .b ({new_AGEMA_signal_2076, Midori_rounds_sub_sBox_PRINCE_2_n12}), .clk (clk), .r (Fresh[228]), .c ({new_AGEMA_signal_2153, Midori_rounds_SR_Result[10]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .a ({new_AGEMA_signal_6281, new_AGEMA_signal_6277}), .b ({new_AGEMA_signal_2078, Midori_rounds_sub_sBox_PRINCE_2_n3}), .clk (clk), .r (Fresh[229]), .c ({new_AGEMA_signal_2155, Midori_rounds_SR_Result[8]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .a ({new_AGEMA_signal_6285, new_AGEMA_signal_6283}), .b ({new_AGEMA_signal_2081, Midori_rounds_sub_sBox_PRINCE_3_n12}), .clk (clk), .r (Fresh[230]), .c ({new_AGEMA_signal_2157, Midori_rounds_SR_Result[22]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .a ({new_AGEMA_signal_6293, new_AGEMA_signal_6289}), .b ({new_AGEMA_signal_2083, Midori_rounds_sub_sBox_PRINCE_3_n3}), .clk (clk), .r (Fresh[231]), .c ({new_AGEMA_signal_2159, Midori_rounds_SR_Result[20]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .a ({new_AGEMA_signal_6297, new_AGEMA_signal_6295}), .b ({new_AGEMA_signal_2086, Midori_rounds_sub_sBox_PRINCE_4_n12}), .clk (clk), .r (Fresh[232]), .c ({new_AGEMA_signal_2161, Midori_rounds_SR_Result[38]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .a ({new_AGEMA_signal_6305, new_AGEMA_signal_6301}), .b ({new_AGEMA_signal_2088, Midori_rounds_sub_sBox_PRINCE_4_n3}), .clk (clk), .r (Fresh[233]), .c ({new_AGEMA_signal_2163, Midori_rounds_SR_Result[36]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .a ({new_AGEMA_signal_6309, new_AGEMA_signal_6307}), .b ({new_AGEMA_signal_2091, Midori_rounds_sub_sBox_PRINCE_5_n12}), .clk (clk), .r (Fresh[234]), .c ({new_AGEMA_signal_2165, Midori_rounds_SR_Result[58]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .a ({new_AGEMA_signal_6317, new_AGEMA_signal_6313}), .b ({new_AGEMA_signal_2093, Midori_rounds_sub_sBox_PRINCE_5_n3}), .clk (clk), .r (Fresh[235]), .c ({new_AGEMA_signal_2167, Midori_rounds_SR_Result[56]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .a ({new_AGEMA_signal_6321, new_AGEMA_signal_6319}), .b ({new_AGEMA_signal_2096, Midori_rounds_sub_sBox_PRINCE_6_n12}), .clk (clk), .r (Fresh[236]), .c ({new_AGEMA_signal_2169, Midori_rounds_SR_Result[30]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .a ({new_AGEMA_signal_6329, new_AGEMA_signal_6325}), .b ({new_AGEMA_signal_2098, Midori_rounds_sub_sBox_PRINCE_6_n3}), .clk (clk), .r (Fresh[237]), .c ({new_AGEMA_signal_2171, Midori_rounds_SR_Result[28]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .a ({new_AGEMA_signal_6333, new_AGEMA_signal_6331}), .b ({new_AGEMA_signal_2101, Midori_rounds_sub_sBox_PRINCE_7_n12}), .clk (clk), .r (Fresh[238]), .c ({new_AGEMA_signal_2173, Midori_rounds_SR_Result[2]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .a ({new_AGEMA_signal_6341, new_AGEMA_signal_6337}), .b ({new_AGEMA_signal_2103, Midori_rounds_sub_sBox_PRINCE_7_n3}), .clk (clk), .r (Fresh[239]), .c ({new_AGEMA_signal_2175, Midori_rounds_SR_Result[0]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .a ({new_AGEMA_signal_6345, new_AGEMA_signal_6343}), .b ({new_AGEMA_signal_2106, Midori_rounds_sub_sBox_PRINCE_8_n12}), .clk (clk), .r (Fresh[240]), .c ({new_AGEMA_signal_2177, Midori_rounds_SR_Result[14]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .a ({new_AGEMA_signal_6353, new_AGEMA_signal_6349}), .b ({new_AGEMA_signal_2108, Midori_rounds_sub_sBox_PRINCE_8_n3}), .clk (clk), .r (Fresh[241]), .c ({new_AGEMA_signal_2179, Midori_rounds_SR_Result[12]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .a ({new_AGEMA_signal_6357, new_AGEMA_signal_6355}), .b ({new_AGEMA_signal_2111, Midori_rounds_sub_sBox_PRINCE_9_n12}), .clk (clk), .r (Fresh[242]), .c ({new_AGEMA_signal_2181, Midori_rounds_SR_Result[18]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .a ({new_AGEMA_signal_6365, new_AGEMA_signal_6361}), .b ({new_AGEMA_signal_2113, Midori_rounds_sub_sBox_PRINCE_9_n3}), .clk (clk), .r (Fresh[243]), .c ({new_AGEMA_signal_2183, Midori_rounds_SR_Result[16]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .a ({new_AGEMA_signal_6369, new_AGEMA_signal_6367}), .b ({new_AGEMA_signal_2116, Midori_rounds_sub_sBox_PRINCE_10_n12}), .clk (clk), .r (Fresh[244]), .c ({new_AGEMA_signal_2185, Midori_rounds_SR_Result[54]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .a ({new_AGEMA_signal_6377, new_AGEMA_signal_6373}), .b ({new_AGEMA_signal_2118, Midori_rounds_sub_sBox_PRINCE_10_n3}), .clk (clk), .r (Fresh[245]), .c ({new_AGEMA_signal_2187, Midori_rounds_SR_Result[52]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .a ({new_AGEMA_signal_6381, new_AGEMA_signal_6379}), .b ({new_AGEMA_signal_2121, Midori_rounds_sub_sBox_PRINCE_11_n12}), .clk (clk), .r (Fresh[246]), .c ({new_AGEMA_signal_2189, Midori_rounds_SR_Result[42]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .a ({new_AGEMA_signal_6389, new_AGEMA_signal_6385}), .b ({new_AGEMA_signal_2123, Midori_rounds_sub_sBox_PRINCE_11_n3}), .clk (clk), .r (Fresh[247]), .c ({new_AGEMA_signal_2191, Midori_rounds_SR_Result[40]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6391}), .b ({new_AGEMA_signal_2126, Midori_rounds_sub_sBox_PRINCE_12_n12}), .clk (clk), .r (Fresh[248]), .c ({new_AGEMA_signal_2193, Midori_rounds_SR_Result[26]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .a ({new_AGEMA_signal_6401, new_AGEMA_signal_6397}), .b ({new_AGEMA_signal_2128, Midori_rounds_sub_sBox_PRINCE_12_n3}), .clk (clk), .r (Fresh[249]), .c ({new_AGEMA_signal_2195, Midori_rounds_SR_Result[24]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .a ({new_AGEMA_signal_6405, new_AGEMA_signal_6403}), .b ({new_AGEMA_signal_2131, Midori_rounds_sub_sBox_PRINCE_13_n12}), .clk (clk), .r (Fresh[250]), .c ({new_AGEMA_signal_2197, Midori_rounds_SR_Result[6]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .a ({new_AGEMA_signal_6413, new_AGEMA_signal_6409}), .b ({new_AGEMA_signal_2133, Midori_rounds_sub_sBox_PRINCE_13_n3}), .clk (clk), .r (Fresh[251]), .c ({new_AGEMA_signal_2199, Midori_rounds_SR_Result[4]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .a ({new_AGEMA_signal_6417, new_AGEMA_signal_6415}), .b ({new_AGEMA_signal_2136, Midori_rounds_sub_sBox_PRINCE_14_n12}), .clk (clk), .r (Fresh[252]), .c ({new_AGEMA_signal_2201, Midori_rounds_SR_Result[34]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .a ({new_AGEMA_signal_6425, new_AGEMA_signal_6421}), .b ({new_AGEMA_signal_2138, Midori_rounds_sub_sBox_PRINCE_14_n3}), .clk (clk), .r (Fresh[253]), .c ({new_AGEMA_signal_2203, Midori_rounds_SR_Result[32]}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .a ({new_AGEMA_signal_6429, new_AGEMA_signal_6427}), .b ({new_AGEMA_signal_2141, Midori_rounds_sub_sBox_PRINCE_15_n12}), .clk (clk), .r (Fresh[254]), .c ({new_AGEMA_signal_2205, Midori_rounds_SR_Result[62]}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .a ({new_AGEMA_signal_6437, new_AGEMA_signal_6433}), .b ({new_AGEMA_signal_2143, Midori_rounds_sub_sBox_PRINCE_15_n3}), .clk (clk), .r (Fresh[255]), .c ({new_AGEMA_signal_2207, Midori_rounds_SR_Result[60]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_0_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2175, Midori_rounds_SR_Result[0]}), .a ({new_AGEMA_signal_2563, Midori_rounds_sub_ResultXORkey[0]}), .c ({new_AGEMA_signal_2619, Midori_rounds_mul_input[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_2_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2173, Midori_rounds_SR_Result[2]}), .a ({new_AGEMA_signal_2303, Midori_rounds_sub_ResultXORkey[2]}), .c ({new_AGEMA_signal_2321, Midori_rounds_mul_input[2]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_4_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2199, Midori_rounds_SR_Result[4]}), .a ({new_AGEMA_signal_2557, Midori_rounds_sub_ResultXORkey[4]}), .c ({new_AGEMA_signal_2620, Midori_rounds_mul_input[4]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_6_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2197, Midori_rounds_SR_Result[6]}), .a ({new_AGEMA_signal_2274, Midori_rounds_sub_ResultXORkey[6]}), .c ({new_AGEMA_signal_2324, Midori_rounds_mul_input[6]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_8_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2155, Midori_rounds_SR_Result[8]}), .a ({new_AGEMA_signal_2492, Midori_rounds_sub_ResultXORkey[8]}), .c ({new_AGEMA_signal_2613, Midori_rounds_mul_input[8]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_10_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2153, Midori_rounds_SR_Result[10]}), .a ({new_AGEMA_signal_2319, Midori_rounds_sub_ResultXORkey[10]}), .c ({new_AGEMA_signal_2327, Midori_rounds_mul_input[10]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_12_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2179, Midori_rounds_SR_Result[12]}), .a ({new_AGEMA_signal_2562, Midori_rounds_sub_ResultXORkey[12]}), .c ({new_AGEMA_signal_2621, Midori_rounds_mul_input[12]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_14_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2177, Midori_rounds_SR_Result[14]}), .a ({new_AGEMA_signal_2316, Midori_rounds_sub_ResultXORkey[14]}), .c ({new_AGEMA_signal_2330, Midori_rounds_mul_input[14]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_16_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2183, Midori_rounds_SR_Result[16]}), .a ({new_AGEMA_signal_2561, Midori_rounds_sub_ResultXORkey[16]}), .c ({new_AGEMA_signal_2622, Midori_rounds_mul_input[16]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_18_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2181, Midori_rounds_SR_Result[18]}), .a ({new_AGEMA_signal_2313, Midori_rounds_sub_ResultXORkey[18]}), .c ({new_AGEMA_signal_2333, Midori_rounds_mul_input[18]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_20_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2159, Midori_rounds_SR_Result[20]}), .a ({new_AGEMA_signal_2495, Midori_rounds_sub_ResultXORkey[20]}), .c ({new_AGEMA_signal_2614, Midori_rounds_mul_input[20]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_22_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2157, Midori_rounds_SR_Result[22]}), .a ({new_AGEMA_signal_2309, Midori_rounds_sub_ResultXORkey[22]}), .c ({new_AGEMA_signal_2336, Midori_rounds_mul_input[22]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_24_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2195, Midori_rounds_SR_Result[24]}), .a ({new_AGEMA_signal_2560, Midori_rounds_sub_ResultXORkey[24]}), .c ({new_AGEMA_signal_2623, Midori_rounds_mul_input[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_26_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2193, Midori_rounds_SR_Result[26]}), .a ({new_AGEMA_signal_2306, Midori_rounds_sub_ResultXORkey[26]}), .c ({new_AGEMA_signal_2339, Midori_rounds_mul_input[26]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_28_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2171, Midori_rounds_SR_Result[28]}), .a ({new_AGEMA_signal_2617, Midori_rounds_sub_ResultXORkey[28]}), .c ({new_AGEMA_signal_2630, Midori_rounds_mul_input[28]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_30_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2169, Midori_rounds_SR_Result[30]}), .a ({new_AGEMA_signal_2302, Midori_rounds_sub_ResultXORkey[30]}), .c ({new_AGEMA_signal_2342, Midori_rounds_mul_input[30]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_32_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2203, Midori_rounds_SR_Result[32]}), .a ({new_AGEMA_signal_2559, Midori_rounds_sub_ResultXORkey[32]}), .c ({new_AGEMA_signal_2624, Midori_rounds_mul_input[32]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_34_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2201, Midori_rounds_SR_Result[34]}), .a ({new_AGEMA_signal_2299, Midori_rounds_sub_ResultXORkey[34]}), .c ({new_AGEMA_signal_2345, Midori_rounds_mul_input[34]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_36_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2163, Midori_rounds_SR_Result[36]}), .a ({new_AGEMA_signal_2494, Midori_rounds_sub_ResultXORkey[36]}), .c ({new_AGEMA_signal_2615, Midori_rounds_mul_input[36]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_38_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2161, Midori_rounds_SR_Result[38]}), .a ({new_AGEMA_signal_2296, Midori_rounds_sub_ResultXORkey[38]}), .c ({new_AGEMA_signal_2348, Midori_rounds_mul_input[38]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_40_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2191, Midori_rounds_SR_Result[40]}), .a ({new_AGEMA_signal_2558, Midori_rounds_sub_ResultXORkey[40]}), .c ({new_AGEMA_signal_2625, Midori_rounds_mul_input[40]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_42_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2189, Midori_rounds_SR_Result[42]}), .a ({new_AGEMA_signal_2292, Midori_rounds_sub_ResultXORkey[42]}), .c ({new_AGEMA_signal_2351, Midori_rounds_mul_input[42]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_44_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2151, Midori_rounds_SR_Result[44]}), .a ({new_AGEMA_signal_2493, Midori_rounds_sub_ResultXORkey[44]}), .c ({new_AGEMA_signal_2616, Midori_rounds_mul_input[44]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_46_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2149, Midori_rounds_SR_Result[46]}), .a ({new_AGEMA_signal_2289, Midori_rounds_sub_ResultXORkey[46]}), .c ({new_AGEMA_signal_2354, Midori_rounds_mul_input[46]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_48_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2147, Midori_rounds_SR_Result[48]}), .a ({new_AGEMA_signal_2629, Midori_rounds_sub_ResultXORkey[48]}), .c ({new_AGEMA_signal_2637, Midori_rounds_mul_input[48]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_50_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2145, Midori_rounds_SR_Result[50]}), .a ({new_AGEMA_signal_2286, Midori_rounds_sub_ResultXORkey[50]}), .c ({new_AGEMA_signal_2357, Midori_rounds_mul_input[50]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_52_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2187, Midori_rounds_SR_Result[52]}), .a ({new_AGEMA_signal_2556, Midori_rounds_sub_ResultXORkey[52]}), .c ({new_AGEMA_signal_2626, Midori_rounds_mul_input[52]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_54_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2185, Midori_rounds_SR_Result[54]}), .a ({new_AGEMA_signal_2283, Midori_rounds_sub_ResultXORkey[54]}), .c ({new_AGEMA_signal_2360, Midori_rounds_mul_input[54]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_56_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2167, Midori_rounds_SR_Result[56]}), .a ({new_AGEMA_signal_2555, Midori_rounds_sub_ResultXORkey[56]}), .c ({new_AGEMA_signal_2627, Midori_rounds_mul_input[56]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_58_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2165, Midori_rounds_SR_Result[58]}), .a ({new_AGEMA_signal_2280, Midori_rounds_sub_ResultXORkey[58]}), .c ({new_AGEMA_signal_2363, Midori_rounds_mul_input[58]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_60_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2207, Midori_rounds_SR_Result[60]}), .a ({new_AGEMA_signal_2554, Midori_rounds_sub_ResultXORkey[60]}), .c ({new_AGEMA_signal_2628, Midori_rounds_mul_input[60]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_input_Inst_mux_inst_62_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2205, Midori_rounds_SR_Result[62]}), .a ({new_AGEMA_signal_2276, Midori_rounds_sub_ResultXORkey[62]}), .c ({new_AGEMA_signal_2366, Midori_rounds_mul_input[62]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U23 ( .a ({new_AGEMA_signal_2628, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_2662, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_2668, Midori_rounds_SR_Inv_Result[20]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U21 ( .a ({new_AGEMA_signal_2357, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_2369, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_2394, Midori_rounds_SR_Inv_Result[42]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U19 ( .a ({new_AGEMA_signal_2637, Midori_rounds_mul_input[48]}), .b ({new_AGEMA_signal_2631, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_2661, Midori_rounds_SR_Inv_Result[40]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U16 ( .a ({new_AGEMA_signal_2360, Midori_rounds_mul_input[54]}), .b ({new_AGEMA_signal_2369, Midori_rounds_mul_MC1_n5}), .c ({new_AGEMA_signal_2397, Midori_rounds_SR_Inv_Result[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U15 ( .a ({new_AGEMA_signal_2366, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_2363, Midori_rounds_mul_input[58]}), .c ({new_AGEMA_signal_2369, Midori_rounds_mul_MC1_n5}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U11 ( .a ({new_AGEMA_signal_2363, Midori_rounds_mul_input[58]}), .b ({new_AGEMA_signal_2373, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_2400, Midori_rounds_SR_Inv_Result[62]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U8 ( .a ({new_AGEMA_signal_2627, Midori_rounds_mul_input[56]}), .b ({new_AGEMA_signal_2662, Midori_rounds_mul_MC1_n7}), .c ({new_AGEMA_signal_2669, Midori_rounds_SR_Inv_Result[60]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U7 ( .a ({new_AGEMA_signal_2626, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_2637, Midori_rounds_mul_input[48]}), .c ({new_AGEMA_signal_2662, Midori_rounds_mul_MC1_n7}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U4 ( .a ({new_AGEMA_signal_2366, Midori_rounds_mul_input[62]}), .b ({new_AGEMA_signal_2373, Midori_rounds_mul_MC1_n1}), .c ({new_AGEMA_signal_2403, Midori_rounds_SR_Inv_Result[22]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U3 ( .a ({new_AGEMA_signal_2357, Midori_rounds_mul_input[50]}), .b ({new_AGEMA_signal_2360, Midori_rounds_mul_input[54]}), .c ({new_AGEMA_signal_2373, Midori_rounds_mul_MC1_n1}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U2 ( .a ({new_AGEMA_signal_2626, Midori_rounds_mul_input[52]}), .b ({new_AGEMA_signal_2631, Midori_rounds_mul_MC1_n3}), .c ({new_AGEMA_signal_2638, Midori_rounds_SR_Inv_Result[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC1_U1 ( .a ({new_AGEMA_signal_2628, Midori_rounds_mul_input[60]}), .b ({new_AGEMA_signal_2627, Midori_rounds_mul_input[56]}), .c ({new_AGEMA_signal_2631, Midori_rounds_mul_MC1_n3}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U23 ( .a ({new_AGEMA_signal_2616, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_2632, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_2639, Midori_rounds_SR_Inv_Result[44]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U21 ( .a ({new_AGEMA_signal_2345, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_2375, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_2406, Midori_rounds_SR_Inv_Result[18]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U19 ( .a ({new_AGEMA_signal_2624, Midori_rounds_mul_input[32]}), .b ({new_AGEMA_signal_2633, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_2640, Midori_rounds_SR_Inv_Result[16]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U16 ( .a ({new_AGEMA_signal_2348, Midori_rounds_mul_input[38]}), .b ({new_AGEMA_signal_2375, Midori_rounds_mul_MC2_n5}), .c ({new_AGEMA_signal_2409, Midori_rounds_SR_Inv_Result[58]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U15 ( .a ({new_AGEMA_signal_2354, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_2351, Midori_rounds_mul_input[42]}), .c ({new_AGEMA_signal_2375, Midori_rounds_mul_MC2_n5}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U11 ( .a ({new_AGEMA_signal_2351, Midori_rounds_mul_input[42]}), .b ({new_AGEMA_signal_2379, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_2412, Midori_rounds_SR_Inv_Result[6]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U8 ( .a ({new_AGEMA_signal_2625, Midori_rounds_mul_input[40]}), .b ({new_AGEMA_signal_2632, Midori_rounds_mul_MC2_n7}), .c ({new_AGEMA_signal_2641, Midori_rounds_SR_Inv_Result[4]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U7 ( .a ({new_AGEMA_signal_2615, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_2624, Midori_rounds_mul_input[32]}), .c ({new_AGEMA_signal_2632, Midori_rounds_mul_MC2_n7}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U4 ( .a ({new_AGEMA_signal_2354, Midori_rounds_mul_input[46]}), .b ({new_AGEMA_signal_2379, Midori_rounds_mul_MC2_n1}), .c ({new_AGEMA_signal_2415, Midori_rounds_SR_Inv_Result[46]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U3 ( .a ({new_AGEMA_signal_2345, Midori_rounds_mul_input[34]}), .b ({new_AGEMA_signal_2348, Midori_rounds_mul_input[38]}), .c ({new_AGEMA_signal_2379, Midori_rounds_mul_MC2_n1}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U2 ( .a ({new_AGEMA_signal_2615, Midori_rounds_mul_input[36]}), .b ({new_AGEMA_signal_2633, Midori_rounds_mul_MC2_n3}), .c ({new_AGEMA_signal_2642, Midori_rounds_SR_Inv_Result[56]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC2_U1 ( .a ({new_AGEMA_signal_2616, Midori_rounds_mul_input[44]}), .b ({new_AGEMA_signal_2625, Midori_rounds_mul_input[40]}), .c ({new_AGEMA_signal_2633, Midori_rounds_mul_MC2_n3}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U23 ( .a ({new_AGEMA_signal_2630, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_2634, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_2643, Midori_rounds_SR_Inv_Result[48]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U21 ( .a ({new_AGEMA_signal_2333, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_2381, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_2418, Midori_rounds_SR_Inv_Result[14]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U19 ( .a ({new_AGEMA_signal_2622, Midori_rounds_mul_input[16]}), .b ({new_AGEMA_signal_2645, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_2663, Midori_rounds_SR_Inv_Result[12]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U16 ( .a ({new_AGEMA_signal_2336, Midori_rounds_mul_input[22]}), .b ({new_AGEMA_signal_2381, Midori_rounds_mul_MC3_n5}), .c ({new_AGEMA_signal_2421, Midori_rounds_SR_Inv_Result[38]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U15 ( .a ({new_AGEMA_signal_2342, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_2339, Midori_rounds_mul_input[26]}), .c ({new_AGEMA_signal_2381, Midori_rounds_mul_MC3_n5}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U11 ( .a ({new_AGEMA_signal_2339, Midori_rounds_mul_input[26]}), .b ({new_AGEMA_signal_2385, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_2424, Midori_rounds_SR_Inv_Result[26]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U8 ( .a ({new_AGEMA_signal_2623, Midori_rounds_mul_input[24]}), .b ({new_AGEMA_signal_2634, Midori_rounds_mul_MC3_n7}), .c ({new_AGEMA_signal_2644, Midori_rounds_SR_Inv_Result[24]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U7 ( .a ({new_AGEMA_signal_2614, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_2622, Midori_rounds_mul_input[16]}), .c ({new_AGEMA_signal_2634, Midori_rounds_mul_MC3_n7}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U4 ( .a ({new_AGEMA_signal_2342, Midori_rounds_mul_input[30]}), .b ({new_AGEMA_signal_2385, Midori_rounds_mul_MC3_n1}), .c ({new_AGEMA_signal_2427, Midori_rounds_SR_Inv_Result[50]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U3 ( .a ({new_AGEMA_signal_2333, Midori_rounds_mul_input[18]}), .b ({new_AGEMA_signal_2336, Midori_rounds_mul_input[22]}), .c ({new_AGEMA_signal_2385, Midori_rounds_mul_MC3_n1}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U2 ( .a ({new_AGEMA_signal_2614, Midori_rounds_mul_input[20]}), .b ({new_AGEMA_signal_2645, Midori_rounds_mul_MC3_n3}), .c ({new_AGEMA_signal_2664, Midori_rounds_SR_Inv_Result[36]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC3_U1 ( .a ({new_AGEMA_signal_2630, Midori_rounds_mul_input[28]}), .b ({new_AGEMA_signal_2623, Midori_rounds_mul_input[24]}), .c ({new_AGEMA_signal_2645, Midori_rounds_mul_MC3_n3}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U23 ( .a ({new_AGEMA_signal_2621, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_2635, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_2646, Midori_rounds_SR_Inv_Result[8]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U21 ( .a ({new_AGEMA_signal_2321, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_2387, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_2430, Midori_rounds_SR_Inv_Result[54]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U19 ( .a ({new_AGEMA_signal_2619, Midori_rounds_mul_input[0]}), .b ({new_AGEMA_signal_2636, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_2647, Midori_rounds_SR_Inv_Result[52]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U16 ( .a ({new_AGEMA_signal_2324, Midori_rounds_mul_input[6]}), .b ({new_AGEMA_signal_2387, Midori_rounds_mul_MC4_n5}), .c ({new_AGEMA_signal_2433, Midori_rounds_SR_Inv_Result[30]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U15 ( .a ({new_AGEMA_signal_2330, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_2327, Midori_rounds_mul_input[10]}), .c ({new_AGEMA_signal_2387, Midori_rounds_mul_MC4_n5}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U11 ( .a ({new_AGEMA_signal_2327, Midori_rounds_mul_input[10]}), .b ({new_AGEMA_signal_2391, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_2436, Midori_rounds_SR_Inv_Result[34]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U8 ( .a ({new_AGEMA_signal_2613, Midori_rounds_mul_input[8]}), .b ({new_AGEMA_signal_2635, Midori_rounds_mul_MC4_n7}), .c ({new_AGEMA_signal_2648, Midori_rounds_SR_Inv_Result[32]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U7 ( .a ({new_AGEMA_signal_2620, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_2619, Midori_rounds_mul_input[0]}), .c ({new_AGEMA_signal_2635, Midori_rounds_mul_MC4_n7}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U4 ( .a ({new_AGEMA_signal_2330, Midori_rounds_mul_input[14]}), .b ({new_AGEMA_signal_2391, Midori_rounds_mul_MC4_n1}), .c ({new_AGEMA_signal_2439, Midori_rounds_SR_Inv_Result[10]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U3 ( .a ({new_AGEMA_signal_2321, Midori_rounds_mul_input[2]}), .b ({new_AGEMA_signal_2324, Midori_rounds_mul_input[6]}), .c ({new_AGEMA_signal_2391, Midori_rounds_mul_MC4_n1}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U2 ( .a ({new_AGEMA_signal_2620, Midori_rounds_mul_input[4]}), .b ({new_AGEMA_signal_2636, Midori_rounds_mul_MC4_n3}), .c ({new_AGEMA_signal_2649, Midori_rounds_SR_Inv_Result[28]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) Midori_rounds_mul_MC4_U1 ( .a ({new_AGEMA_signal_2621, Midori_rounds_mul_input[12]}), .b ({new_AGEMA_signal_2613, Midori_rounds_mul_input[8]}), .c ({new_AGEMA_signal_2636, Midori_rounds_mul_MC4_n3}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_0_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2660, Midori_rounds_mul_ResultXORkey[0]}), .a ({new_AGEMA_signal_2638, Midori_rounds_SR_Inv_Result[0]}), .c ({new_AGEMA_signal_2670, Midori_rounds_round_Result[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_2_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2474, Midori_rounds_mul_ResultXORkey[2]}), .a ({new_AGEMA_signal_2397, Midori_rounds_SR_Inv_Result[2]}), .c ({new_AGEMA_signal_2507, Midori_rounds_round_Result[2]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_4_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2651, Midori_rounds_mul_ResultXORkey[4]}), .a ({new_AGEMA_signal_2641, Midori_rounds_SR_Inv_Result[4]}), .c ({new_AGEMA_signal_2671, Midori_rounds_round_Result[4]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_6_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2443, Midori_rounds_mul_ResultXORkey[6]}), .a ({new_AGEMA_signal_2412, Midori_rounds_SR_Inv_Result[6]}), .c ({new_AGEMA_signal_2510, Midori_rounds_round_Result[6]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_8_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2650, Midori_rounds_mul_ResultXORkey[8]}), .a ({new_AGEMA_signal_2646, Midori_rounds_SR_Inv_Result[8]}), .c ({new_AGEMA_signal_2672, Midori_rounds_round_Result[8]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_10_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2491, Midori_rounds_mul_ResultXORkey[10]}), .a ({new_AGEMA_signal_2439, Midori_rounds_SR_Inv_Result[10]}), .c ({new_AGEMA_signal_2513, Midori_rounds_round_Result[10]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_12_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2659, Midori_rounds_mul_ResultXORkey[12]}), .a ({new_AGEMA_signal_2663, Midori_rounds_SR_Inv_Result[12]}), .c ({new_AGEMA_signal_2673, Midori_rounds_round_Result[12]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_14_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2488, Midori_rounds_mul_ResultXORkey[14]}), .a ({new_AGEMA_signal_2418, Midori_rounds_SR_Inv_Result[14]}), .c ({new_AGEMA_signal_2516, Midori_rounds_round_Result[14]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_16_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2667, Midori_rounds_mul_ResultXORkey[16]}), .a ({new_AGEMA_signal_2640, Midori_rounds_SR_Inv_Result[16]}), .c ({new_AGEMA_signal_2694, Midori_rounds_round_Result[16]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_18_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2485, Midori_rounds_mul_ResultXORkey[18]}), .a ({new_AGEMA_signal_2406, Midori_rounds_SR_Inv_Result[18]}), .c ({new_AGEMA_signal_2519, Midori_rounds_round_Result[18]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_20_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2666, Midori_rounds_mul_ResultXORkey[20]}), .a ({new_AGEMA_signal_2668, Midori_rounds_SR_Inv_Result[20]}), .c ({new_AGEMA_signal_2695, Midori_rounds_round_Result[20]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_22_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2480, Midori_rounds_mul_ResultXORkey[22]}), .a ({new_AGEMA_signal_2403, Midori_rounds_SR_Inv_Result[22]}), .c ({new_AGEMA_signal_2522, Midori_rounds_round_Result[22]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_24_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2658, Midori_rounds_mul_ResultXORkey[24]}), .a ({new_AGEMA_signal_2644, Midori_rounds_SR_Inv_Result[24]}), .c ({new_AGEMA_signal_2674, Midori_rounds_round_Result[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_26_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2477, Midori_rounds_mul_ResultXORkey[26]}), .a ({new_AGEMA_signal_2424, Midori_rounds_SR_Inv_Result[26]}), .c ({new_AGEMA_signal_2525, Midori_rounds_round_Result[26]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_28_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2657, Midori_rounds_mul_ResultXORkey[28]}), .a ({new_AGEMA_signal_2649, Midori_rounds_SR_Inv_Result[28]}), .c ({new_AGEMA_signal_2675, Midori_rounds_round_Result[28]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_30_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2473, Midori_rounds_mul_ResultXORkey[30]}), .a ({new_AGEMA_signal_2433, Midori_rounds_SR_Inv_Result[30]}), .c ({new_AGEMA_signal_2528, Midori_rounds_round_Result[30]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_32_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2656, Midori_rounds_mul_ResultXORkey[32]}), .a ({new_AGEMA_signal_2648, Midori_rounds_SR_Inv_Result[32]}), .c ({new_AGEMA_signal_2676, Midori_rounds_round_Result[32]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_34_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2470, Midori_rounds_mul_ResultXORkey[34]}), .a ({new_AGEMA_signal_2436, Midori_rounds_SR_Inv_Result[34]}), .c ({new_AGEMA_signal_2531, Midori_rounds_round_Result[34]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_36_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2655, Midori_rounds_mul_ResultXORkey[36]}), .a ({new_AGEMA_signal_2664, Midori_rounds_SR_Inv_Result[36]}), .c ({new_AGEMA_signal_2677, Midori_rounds_round_Result[36]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_38_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2466, Midori_rounds_mul_ResultXORkey[38]}), .a ({new_AGEMA_signal_2421, Midori_rounds_SR_Inv_Result[38]}), .c ({new_AGEMA_signal_2534, Midori_rounds_round_Result[38]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_40_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2654, Midori_rounds_mul_ResultXORkey[40]}), .a ({new_AGEMA_signal_2661, Midori_rounds_SR_Inv_Result[40]}), .c ({new_AGEMA_signal_2678, Midori_rounds_round_Result[40]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_42_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2462, Midori_rounds_mul_ResultXORkey[42]}), .a ({new_AGEMA_signal_2394, Midori_rounds_SR_Inv_Result[42]}), .c ({new_AGEMA_signal_2537, Midori_rounds_round_Result[42]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_44_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2653, Midori_rounds_mul_ResultXORkey[44]}), .a ({new_AGEMA_signal_2639, Midori_rounds_SR_Inv_Result[44]}), .c ({new_AGEMA_signal_2679, Midori_rounds_round_Result[44]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_46_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2458, Midori_rounds_mul_ResultXORkey[46]}), .a ({new_AGEMA_signal_2415, Midori_rounds_SR_Inv_Result[46]}), .c ({new_AGEMA_signal_2540, Midori_rounds_round_Result[46]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_48_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2652, Midori_rounds_mul_ResultXORkey[48]}), .a ({new_AGEMA_signal_2643, Midori_rounds_SR_Inv_Result[48]}), .c ({new_AGEMA_signal_2680, Midori_rounds_round_Result[48]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_50_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2455, Midori_rounds_mul_ResultXORkey[50]}), .a ({new_AGEMA_signal_2427, Midori_rounds_SR_Inv_Result[50]}), .c ({new_AGEMA_signal_2543, Midori_rounds_round_Result[50]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_52_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2665, Midori_rounds_mul_ResultXORkey[52]}), .a ({new_AGEMA_signal_2647, Midori_rounds_SR_Inv_Result[52]}), .c ({new_AGEMA_signal_2696, Midori_rounds_round_Result[52]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_54_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2452, Midori_rounds_mul_ResultXORkey[54]}), .a ({new_AGEMA_signal_2430, Midori_rounds_SR_Inv_Result[54]}), .c ({new_AGEMA_signal_2546, Midori_rounds_round_Result[54]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_56_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2682, Midori_rounds_mul_ResultXORkey[56]}), .a ({new_AGEMA_signal_2642, Midori_rounds_SR_Inv_Result[56]}), .c ({new_AGEMA_signal_2700, Midori_rounds_round_Result[56]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_58_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2449, Midori_rounds_mul_ResultXORkey[58]}), .a ({new_AGEMA_signal_2409, Midori_rounds_SR_Inv_Result[58]}), .c ({new_AGEMA_signal_2549, Midori_rounds_round_Result[58]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_60_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2681, Midori_rounds_mul_ResultXORkey[60]}), .a ({new_AGEMA_signal_2669, Midori_rounds_SR_Inv_Result[60]}), .c ({new_AGEMA_signal_2701, Midori_rounds_round_Result[60]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_Res_Inst_mux_inst_62_U1 ( .s (new_AGEMA_signal_6439), .b ({new_AGEMA_signal_2445, Midori_rounds_mul_ResultXORkey[62]}), .a ({new_AGEMA_signal_2400, Midori_rounds_SR_Inv_Result[62]}), .c ({new_AGEMA_signal_2552, Midori_rounds_round_Result[62]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (new_AGEMA_signal_2961), .Q (DataOut_s0[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (new_AGEMA_signal_2963), .Q (DataOut_s0[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_2965), .Q (DataOut_s0[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (new_AGEMA_signal_2967), .Q (DataOut_s0[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_2969), .Q (DataOut_s0[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (new_AGEMA_signal_2971), .Q (DataOut_s0[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_2973), .Q (DataOut_s0[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (new_AGEMA_signal_2975), .Q (DataOut_s0[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_2977), .Q (DataOut_s0[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (new_AGEMA_signal_2979), .Q (DataOut_s0[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_2981), .Q (DataOut_s0[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (new_AGEMA_signal_2983), .Q (DataOut_s0[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_2985), .Q (DataOut_s0[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (new_AGEMA_signal_2987), .Q (DataOut_s0[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_2989), .Q (DataOut_s0[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (new_AGEMA_signal_2991), .Q (DataOut_s0[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_2993), .Q (DataOut_s0[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (new_AGEMA_signal_2995), .Q (DataOut_s0[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_2997), .Q (DataOut_s0[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (new_AGEMA_signal_2999), .Q (DataOut_s0[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_3001), .Q (DataOut_s0[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (new_AGEMA_signal_3003), .Q (DataOut_s0[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_3005), .Q (DataOut_s0[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (DataOut_s0[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_3009), .Q (DataOut_s0[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (new_AGEMA_signal_3011), .Q (DataOut_s0[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_3013), .Q (DataOut_s0[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (new_AGEMA_signal_3015), .Q (DataOut_s0[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_3017), .Q (DataOut_s0[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (new_AGEMA_signal_3019), .Q (DataOut_s0[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_3021), .Q (DataOut_s0[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (new_AGEMA_signal_3023), .Q (DataOut_s0[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (new_AGEMA_signal_3031), .Q (done) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_3033), .Q (DataOut_s1[9]) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (new_AGEMA_signal_3035), .Q (DataOut_s1[7]) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_3037), .Q (DataOut_s1[63]) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (new_AGEMA_signal_3039), .Q (DataOut_s1[61]) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_3041), .Q (DataOut_s1[5]) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (new_AGEMA_signal_3043), .Q (DataOut_s1[59]) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_3045), .Q (DataOut_s1[57]) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (new_AGEMA_signal_3047), .Q (DataOut_s1[55]) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_3049), .Q (DataOut_s1[53]) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (new_AGEMA_signal_3051), .Q (DataOut_s1[51]) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_3053), .Q (DataOut_s1[49]) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (new_AGEMA_signal_3055), .Q (DataOut_s1[47]) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_3057), .Q (DataOut_s1[45]) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (new_AGEMA_signal_3059), .Q (DataOut_s1[43]) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_3061), .Q (DataOut_s1[41]) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (new_AGEMA_signal_3063), .Q (DataOut_s1[3]) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (clk), .D (new_AGEMA_signal_3065), .Q (DataOut_s1[39]) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (clk), .D (new_AGEMA_signal_3067), .Q (DataOut_s1[37]) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (clk), .D (new_AGEMA_signal_3069), .Q (DataOut_s1[35]) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (clk), .D (new_AGEMA_signal_3071), .Q (DataOut_s1[33]) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (clk), .D (new_AGEMA_signal_3073), .Q (DataOut_s1[31]) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (clk), .D (new_AGEMA_signal_3075), .Q (DataOut_s1[29]) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (clk), .D (new_AGEMA_signal_3077), .Q (DataOut_s1[27]) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (clk), .D (new_AGEMA_signal_3079), .Q (DataOut_s1[25]) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (clk), .D (new_AGEMA_signal_3081), .Q (DataOut_s1[23]) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (clk), .D (new_AGEMA_signal_3083), .Q (DataOut_s1[21]) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (clk), .D (new_AGEMA_signal_3085), .Q (DataOut_s1[1]) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (clk), .D (new_AGEMA_signal_3087), .Q (DataOut_s1[19]) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (clk), .D (new_AGEMA_signal_3089), .Q (DataOut_s1[17]) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (clk), .D (new_AGEMA_signal_3091), .Q (DataOut_s1[15]) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (clk), .D (new_AGEMA_signal_3093), .Q (DataOut_s1[13]) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (clk), .D (new_AGEMA_signal_3095), .Q (DataOut_s1[11]) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_4715) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_4723) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_4747) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_4771) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_4795) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_4818), .Q (new_AGEMA_signal_4819) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_4843) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_4866), .Q (new_AGEMA_signal_4867) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_4890), .Q (new_AGEMA_signal_4891) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_4899) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_4907) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_4914), .Q (new_AGEMA_signal_4915) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_4923) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_4931) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_4938), .Q (new_AGEMA_signal_4939) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_4946), .Q (new_AGEMA_signal_4947) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_4955) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_4962), .Q (new_AGEMA_signal_4963) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_4970), .Q (new_AGEMA_signal_4971) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_4979) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_4987) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_4994), .Q (new_AGEMA_signal_4995) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_5003) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_5010), .Q (new_AGEMA_signal_5011) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_5018), .Q (new_AGEMA_signal_5019) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_5027) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_5035) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_5042), .Q (new_AGEMA_signal_5043) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_5051) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_5059) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_5066), .Q (new_AGEMA_signal_5067) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_5075) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_5082), .Q (new_AGEMA_signal_5083) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_5090), .Q (new_AGEMA_signal_5091) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_5099) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_5106), .Q (new_AGEMA_signal_5107) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_5114), .Q (new_AGEMA_signal_5115) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_5123) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_5131) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_5138), .Q (new_AGEMA_signal_5139) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_5147) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_5154), .Q (new_AGEMA_signal_5155) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_5162), .Q (new_AGEMA_signal_5163) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_5171) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_5179) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_5186), .Q (new_AGEMA_signal_5187) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_5195) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_5203) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_5210), .Q (new_AGEMA_signal_5211) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_5219) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_5226), .Q (new_AGEMA_signal_5227) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_5234), .Q (new_AGEMA_signal_5235) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_5243) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_5251) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_5258), .Q (new_AGEMA_signal_5259) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_5267) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_5275) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_5282), .Q (new_AGEMA_signal_5283) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_5291) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_5298), .Q (new_AGEMA_signal_5299) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_5306), .Q (new_AGEMA_signal_5307) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_5314), .Q (new_AGEMA_signal_5315) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_5323) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_5330), .Q (new_AGEMA_signal_5331) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_5339) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_5347) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_5354), .Q (new_AGEMA_signal_5355) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_5363) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_5370), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_5378), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_5386), .Q (new_AGEMA_signal_5387) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_5394), .Q (new_AGEMA_signal_5395) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_5411) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_5419) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_5434), .Q (new_AGEMA_signal_5435) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_5443) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_5450), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_5458), .Q (new_AGEMA_signal_5459) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_5466), .Q (new_AGEMA_signal_5467) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_5474), .Q (new_AGEMA_signal_5475) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_5482), .Q (new_AGEMA_signal_5483) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_5491) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_5499) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_5507) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_5514), .Q (new_AGEMA_signal_5515) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_5523) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_5530), .Q (new_AGEMA_signal_5531) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_5538), .Q (new_AGEMA_signal_5539) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_5546), .Q (new_AGEMA_signal_5547) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_5554), .Q (new_AGEMA_signal_5555) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_5563) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_5570), .Q (new_AGEMA_signal_5571) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_5579) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_5586), .Q (new_AGEMA_signal_5587) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_5594), .Q (new_AGEMA_signal_5595) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_5603) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_5610), .Q (new_AGEMA_signal_5611) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_5618), .Q (new_AGEMA_signal_5619) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_5627) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_5635) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_5643) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_5651) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_5658), .Q (new_AGEMA_signal_5659) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_5666), .Q (new_AGEMA_signal_5667) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_5674), .Q (new_AGEMA_signal_5675) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_5682), .Q (new_AGEMA_signal_5683) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_5690), .Q (new_AGEMA_signal_5691) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_5699) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_5707) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_5714), .Q (new_AGEMA_signal_5715) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_5723) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_5730), .Q (new_AGEMA_signal_5731) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_5861) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_5909) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_5957) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_6005) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_6053) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_6101) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_6149) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_6197) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_6245) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_6439) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_6447) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_6455) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_6463) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_6471) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_6472), .Q (new_AGEMA_signal_6473) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_6474), .Q (new_AGEMA_signal_6475) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_6477) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_6478), .Q (new_AGEMA_signal_6479) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_6481) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_6483) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_6485) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_6487) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_6489) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_6490), .Q (new_AGEMA_signal_6491) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_6493) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_6495) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_6497) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_6498), .Q (new_AGEMA_signal_6499) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_6502), .Q (new_AGEMA_signal_6503) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_6507) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_6509) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_6511) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_6513) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_6514), .Q (new_AGEMA_signal_6515) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_6517) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_6519) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_6520), .Q (new_AGEMA_signal_6521) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_6522), .Q (new_AGEMA_signal_6523) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_6525) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_6526), .Q (new_AGEMA_signal_6527) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_6529) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_6530), .Q (new_AGEMA_signal_6531) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_6533) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_6535) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_6537) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_6538), .Q (new_AGEMA_signal_6539) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_6541) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_6543) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_6545) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_6546), .Q (new_AGEMA_signal_6547) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_6550), .Q (new_AGEMA_signal_6551) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_6553) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_6554), .Q (new_AGEMA_signal_6555) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_6556), .Q (new_AGEMA_signal_6557) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_6559) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_6561) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_6562), .Q (new_AGEMA_signal_6563) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_6564), .Q (new_AGEMA_signal_6565) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_6566), .Q (new_AGEMA_signal_6567) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_6568), .Q (new_AGEMA_signal_6569) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_6570), .Q (new_AGEMA_signal_6571) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_6572), .Q (new_AGEMA_signal_6573) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_6574), .Q (new_AGEMA_signal_6575) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_6577) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_6578), .Q (new_AGEMA_signal_6579) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_6580), .Q (new_AGEMA_signal_6581) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_6582), .Q (new_AGEMA_signal_6583) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_6584), .Q (new_AGEMA_signal_6585) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_6586), .Q (new_AGEMA_signal_6587) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_6588), .Q (new_AGEMA_signal_6589) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_6590), .Q (new_AGEMA_signal_6591) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_6592), .Q (new_AGEMA_signal_6593) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_6594), .Q (new_AGEMA_signal_6595) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_6597) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_6598), .Q (new_AGEMA_signal_6599) ) ;

    /* register cells */
    DFF_X1 controller_roundCounter_count_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6447), .Q (round_Signal[0]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6455), .Q (round_Signal[1]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6463), .Q (round_Signal[2]), .QN () ) ;
    DFF_X1 controller_roundCounter_count_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_6471), .Q (round_Signal[3]), .QN () ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_0_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2683, Midori_rounds_roundResult_Reg_SFF_0_DQ}), .Q ({new_AGEMA_signal_1661, Midori_rounds_roundReg_out[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_1_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6475, new_AGEMA_signal_6473}), .Q ({new_AGEMA_signal_2064, Midori_rounds_roundReg_out[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_2_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2566, Midori_rounds_roundResult_Reg_SFF_2_DQ}), .Q ({new_AGEMA_signal_1664, Midori_rounds_roundReg_out[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_3_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6479, new_AGEMA_signal_6477}), .Q ({new_AGEMA_signal_1662, Midori_rounds_roundReg_out[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_4_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2684, Midori_rounds_roundResult_Reg_SFF_4_DQ}), .Q ({new_AGEMA_signal_1669, Midori_rounds_roundReg_out[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_5_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6483, new_AGEMA_signal_6481}), .Q ({new_AGEMA_signal_2069, Midori_rounds_roundReg_out[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_6_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2569, Midori_rounds_roundResult_Reg_SFF_6_DQ}), .Q ({new_AGEMA_signal_1672, Midori_rounds_roundReg_out[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_7_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6487, new_AGEMA_signal_6485}), .Q ({new_AGEMA_signal_1670, Midori_rounds_roundReg_out[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_8_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2685, Midori_rounds_roundResult_Reg_SFF_8_DQ}), .Q ({new_AGEMA_signal_1677, Midori_rounds_roundReg_out[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_9_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6491, new_AGEMA_signal_6489}), .Q ({new_AGEMA_signal_2074, Midori_rounds_roundReg_out[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_10_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2572, Midori_rounds_roundResult_Reg_SFF_10_DQ}), .Q ({new_AGEMA_signal_1680, Midori_rounds_roundReg_out[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_11_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6495, new_AGEMA_signal_6493}), .Q ({new_AGEMA_signal_1678, Midori_rounds_roundReg_out[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_12_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2686, Midori_rounds_roundResult_Reg_SFF_12_DQ}), .Q ({new_AGEMA_signal_1685, Midori_rounds_roundReg_out[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_13_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6499, new_AGEMA_signal_6497}), .Q ({new_AGEMA_signal_2079, Midori_rounds_roundReg_out[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_14_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2575, Midori_rounds_roundResult_Reg_SFF_14_DQ}), .Q ({new_AGEMA_signal_1688, Midori_rounds_roundReg_out[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_15_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6503, new_AGEMA_signal_6501}), .Q ({new_AGEMA_signal_1686, Midori_rounds_roundReg_out[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_16_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2697, Midori_rounds_roundResult_Reg_SFF_16_DQ}), .Q ({new_AGEMA_signal_1693, Midori_rounds_roundReg_out[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_17_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6507, new_AGEMA_signal_6505}), .Q ({new_AGEMA_signal_2084, Midori_rounds_roundReg_out[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_18_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2578, Midori_rounds_roundResult_Reg_SFF_18_DQ}), .Q ({new_AGEMA_signal_1696, Midori_rounds_roundReg_out[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_19_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6511, new_AGEMA_signal_6509}), .Q ({new_AGEMA_signal_1694, Midori_rounds_roundReg_out[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_20_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2698, Midori_rounds_roundResult_Reg_SFF_20_DQ}), .Q ({new_AGEMA_signal_1701, Midori_rounds_roundReg_out[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_21_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6515, new_AGEMA_signal_6513}), .Q ({new_AGEMA_signal_2089, Midori_rounds_roundReg_out[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_22_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2581, Midori_rounds_roundResult_Reg_SFF_22_DQ}), .Q ({new_AGEMA_signal_1704, Midori_rounds_roundReg_out[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_23_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6519, new_AGEMA_signal_6517}), .Q ({new_AGEMA_signal_1702, Midori_rounds_roundReg_out[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_24_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2687, Midori_rounds_roundResult_Reg_SFF_24_DQ}), .Q ({new_AGEMA_signal_1709, Midori_rounds_roundReg_out[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_25_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6523, new_AGEMA_signal_6521}), .Q ({new_AGEMA_signal_2094, Midori_rounds_roundReg_out[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_26_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2584, Midori_rounds_roundResult_Reg_SFF_26_DQ}), .Q ({new_AGEMA_signal_1712, Midori_rounds_roundReg_out[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_27_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6527, new_AGEMA_signal_6525}), .Q ({new_AGEMA_signal_1710, Midori_rounds_roundReg_out[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_28_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2688, Midori_rounds_roundResult_Reg_SFF_28_DQ}), .Q ({new_AGEMA_signal_1717, Midori_rounds_roundReg_out[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_29_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6531, new_AGEMA_signal_6529}), .Q ({new_AGEMA_signal_2099, Midori_rounds_roundReg_out[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_30_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2587, Midori_rounds_roundResult_Reg_SFF_30_DQ}), .Q ({new_AGEMA_signal_1720, Midori_rounds_roundReg_out[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_31_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6535, new_AGEMA_signal_6533}), .Q ({new_AGEMA_signal_1718, Midori_rounds_roundReg_out[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_32_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2689, Midori_rounds_roundResult_Reg_SFF_32_DQ}), .Q ({new_AGEMA_signal_1725, Midori_rounds_roundReg_out[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_33_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6539, new_AGEMA_signal_6537}), .Q ({new_AGEMA_signal_2104, Midori_rounds_roundReg_out[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_34_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2590, Midori_rounds_roundResult_Reg_SFF_34_DQ}), .Q ({new_AGEMA_signal_1728, Midori_rounds_roundReg_out[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_35_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6543, new_AGEMA_signal_6541}), .Q ({new_AGEMA_signal_1726, Midori_rounds_roundReg_out[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_36_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2690, Midori_rounds_roundResult_Reg_SFF_36_DQ}), .Q ({new_AGEMA_signal_1733, Midori_rounds_roundReg_out[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_37_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6547, new_AGEMA_signal_6545}), .Q ({new_AGEMA_signal_2109, Midori_rounds_roundReg_out[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_38_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2593, Midori_rounds_roundResult_Reg_SFF_38_DQ}), .Q ({new_AGEMA_signal_1736, Midori_rounds_roundReg_out[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_39_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6551, new_AGEMA_signal_6549}), .Q ({new_AGEMA_signal_1734, Midori_rounds_roundReg_out[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_40_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2691, Midori_rounds_roundResult_Reg_SFF_40_DQ}), .Q ({new_AGEMA_signal_1741, Midori_rounds_roundReg_out[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_41_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6555, new_AGEMA_signal_6553}), .Q ({new_AGEMA_signal_2114, Midori_rounds_roundReg_out[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_42_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2596, Midori_rounds_roundResult_Reg_SFF_42_DQ}), .Q ({new_AGEMA_signal_1744, Midori_rounds_roundReg_out[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_43_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6559, new_AGEMA_signal_6557}), .Q ({new_AGEMA_signal_1742, Midori_rounds_roundReg_out[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_44_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2692, Midori_rounds_roundResult_Reg_SFF_44_DQ}), .Q ({new_AGEMA_signal_1749, Midori_rounds_roundReg_out[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_45_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6563, new_AGEMA_signal_6561}), .Q ({new_AGEMA_signal_2119, Midori_rounds_roundReg_out[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_46_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2599, Midori_rounds_roundResult_Reg_SFF_46_DQ}), .Q ({new_AGEMA_signal_1752, Midori_rounds_roundReg_out[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_47_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6567, new_AGEMA_signal_6565}), .Q ({new_AGEMA_signal_1750, Midori_rounds_roundReg_out[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_48_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2693, Midori_rounds_roundResult_Reg_SFF_48_DQ}), .Q ({new_AGEMA_signal_1757, Midori_rounds_roundReg_out[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_49_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6571, new_AGEMA_signal_6569}), .Q ({new_AGEMA_signal_2124, Midori_rounds_roundReg_out[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_50_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2602, Midori_rounds_roundResult_Reg_SFF_50_DQ}), .Q ({new_AGEMA_signal_1760, Midori_rounds_roundReg_out[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_51_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6575, new_AGEMA_signal_6573}), .Q ({new_AGEMA_signal_1758, Midori_rounds_roundReg_out[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_52_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2699, Midori_rounds_roundResult_Reg_SFF_52_DQ}), .Q ({new_AGEMA_signal_1765, Midori_rounds_roundReg_out[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_53_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6579, new_AGEMA_signal_6577}), .Q ({new_AGEMA_signal_2129, Midori_rounds_roundReg_out[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_54_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2605, Midori_rounds_roundResult_Reg_SFF_54_DQ}), .Q ({new_AGEMA_signal_1768, Midori_rounds_roundReg_out[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_55_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6583, new_AGEMA_signal_6581}), .Q ({new_AGEMA_signal_1766, Midori_rounds_roundReg_out[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_56_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2702, Midori_rounds_roundResult_Reg_SFF_56_DQ}), .Q ({new_AGEMA_signal_1773, Midori_rounds_roundReg_out[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_57_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6587, new_AGEMA_signal_6585}), .Q ({new_AGEMA_signal_2134, Midori_rounds_roundReg_out[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_58_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2608, Midori_rounds_roundResult_Reg_SFF_58_DQ}), .Q ({new_AGEMA_signal_1776, Midori_rounds_roundReg_out[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_59_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6591, new_AGEMA_signal_6589}), .Q ({new_AGEMA_signal_1774, Midori_rounds_roundReg_out[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_60_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2703, Midori_rounds_roundResult_Reg_SFF_60_DQ}), .Q ({new_AGEMA_signal_1781, Midori_rounds_roundReg_out[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_61_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6595, new_AGEMA_signal_6593}), .Q ({new_AGEMA_signal_2139, Midori_rounds_roundReg_out[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_62_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2611, Midori_rounds_roundResult_Reg_SFF_62_DQ}), .Q ({new_AGEMA_signal_1784, Midori_rounds_roundReg_out[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) Midori_rounds_roundResult_Reg_SFF_63_Q_reg_FF_FF ( .clk (clk), .D ({new_AGEMA_signal_6599, new_AGEMA_signal_6597}), .Q ({new_AGEMA_signal_1782, Midori_rounds_roundReg_out[63]}) ) ;
endmodule
