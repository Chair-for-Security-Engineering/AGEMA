/* modified netlist. Source: module sbox in file Designs/AESSbox/Canright/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module sbox_HPC1_ClockGating_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, rst, Y_s0, Y_s1, Y_s2, Y_s3, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input rst ;
    input [399:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    output Synch ;
    wire sbe_n10 ;
    wire sbe_n9 ;
    wire sbe_n8 ;
    wire sbe_n7 ;
    wire sbe_n6 ;
    wire sbe_n5 ;
    wire sbe_n4 ;
    wire sbe_n3 ;
    wire sbe_n12 ;
    wire sbe_n11 ;
    wire sbe_n2 ;
    wire sbe_n1 ;
    wire sbe_n25 ;
    wire sbe_n24 ;
    wire sbe_n23 ;
    wire sbe_n22 ;
    wire sbe_n21 ;
    wire sbe_n20 ;
    wire sbe_n19 ;
    wire sbe_n18 ;
    wire sbe_n17 ;
    wire sbe_n16 ;
    wire sbe_n15 ;
    wire sbe_n14 ;
    wire sbe_D_0_ ;
    wire sbe_D_2_ ;
    wire sbe_D_3_ ;
    wire sbe_D_5_ ;
    wire sbe_D_6_ ;
    wire sbe_C_0_ ;
    wire sbe_C_1_ ;
    wire sbe_C_2_ ;
    wire sbe_C_3_ ;
    wire sbe_C_4_ ;
    wire sbe_C_5_ ;
    wire sbe_C_6_ ;
    wire sbe_C_7_ ;
    wire sbe_Y_0_ ;
    wire sbe_Y_1_ ;
    wire sbe_Y_2_ ;
    wire sbe_Y_4_ ;
    wire sbe_Y_5_ ;
    wire sbe_Y_6_ ;
    wire sbe_B_3_ ;
    wire sbe_B_6_ ;
    wire sbe_sel_in_m7_n8 ;
    wire sbe_sel_in_m6_n8 ;
    wire sbe_sel_in_m5_n8 ;
    wire sbe_sel_in_m4_n8 ;
    wire sbe_sel_in_m3_n8 ;
    wire sbe_sel_in_m2_n8 ;
    wire sbe_sel_in_m1_n8 ;
    wire sbe_sel_in_m0_n8 ;
    wire sbe_inv_n21 ;
    wire sbe_inv_n20 ;
    wire sbe_inv_n19 ;
    wire sbe_inv_n18 ;
    wire sbe_inv_n17 ;
    wire sbe_inv_n16 ;
    wire sbe_inv_n15 ;
    wire sbe_inv_n14 ;
    wire sbe_inv_n13 ;
    wire sbe_inv_n12 ;
    wire sbe_inv_n11 ;
    wire sbe_inv_n10 ;
    wire sbe_inv_n9 ;
    wire sbe_inv_n8 ;
    wire sbe_inv_n7 ;
    wire sbe_inv_n6 ;
    wire sbe_inv_n5 ;
    wire sbe_inv_n4 ;
    wire sbe_inv_n3 ;
    wire sbe_inv_n2 ;
    wire sbe_inv_dd ;
    wire sbe_inv_dh ;
    wire sbe_inv_dl ;
    wire sbe_inv_sd_0_ ;
    wire sbe_inv_sd_1_ ;
    wire sbe_inv_d_0_ ;
    wire sbe_inv_d_1_ ;
    wire sbe_inv_d_2_ ;
    wire sbe_inv_d_3_ ;
    wire sbe_inv_bb ;
    wire sbe_inv_bh ;
    wire sbe_inv_bl ;
    wire sbe_inv_aa ;
    wire sbe_inv_ah ;
    wire sbe_inv_al ;
    wire sbe_inv_sb_0_ ;
    wire sbe_inv_sb_1_ ;
    wire sbe_inv_sa_0_ ;
    wire sbe_inv_sa_1_ ;
    wire sbe_inv_dinv_n4 ;
    wire sbe_inv_dinv_n3 ;
    wire sbe_inv_dinv_n2 ;
    wire sbe_inv_dinv_n1 ;
    wire sbe_inv_dinv_sd ;
    wire sbe_inv_dinv_d_0_ ;
    wire sbe_inv_dinv_d_1_ ;
    wire sbe_inv_dinv_sb ;
    wire sbe_inv_dinv_sa ;
    wire sbe_inv_dinv_pmul_n9 ;
    wire sbe_inv_dinv_pmul_n8 ;
    wire sbe_inv_dinv_pmul_n7 ;
    wire sbe_inv_dinv_qmul_n9 ;
    wire sbe_inv_dinv_qmul_n8 ;
    wire sbe_inv_dinv_qmul_n7 ;
    wire sbe_inv_pmul_p_0_ ;
    wire sbe_inv_pmul_p_1_ ;
    wire sbe_inv_pmul_himul_n9 ;
    wire sbe_inv_pmul_himul_n8 ;
    wire sbe_inv_pmul_himul_n7 ;
    wire sbe_inv_pmul_lomul_n9 ;
    wire sbe_inv_pmul_lomul_n8 ;
    wire sbe_inv_pmul_lomul_n7 ;
    wire sbe_inv_pmul_summul_n9 ;
    wire sbe_inv_pmul_summul_n8 ;
    wire sbe_inv_pmul_summul_n7 ;
    wire sbe_inv_qmul_p_0_ ;
    wire sbe_inv_qmul_p_1_ ;
    wire sbe_inv_qmul_himul_n9 ;
    wire sbe_inv_qmul_himul_n8 ;
    wire sbe_inv_qmul_himul_n7 ;
    wire sbe_inv_qmul_lomul_n9 ;
    wire sbe_inv_qmul_lomul_n8 ;
    wire sbe_inv_qmul_lomul_n7 ;
    wire sbe_inv_qmul_summul_n9 ;
    wire sbe_inv_qmul_summul_n8 ;
    wire sbe_inv_qmul_summul_n7 ;
    wire sbe_sel_out_m7_n8 ;
    wire sbe_sel_out_m6_n8 ;
    wire sbe_sel_out_m5_n8 ;
    wire sbe_sel_out_m4_n8 ;
    wire sbe_sel_out_m3_n8 ;
    wire sbe_sel_out_m2_n8 ;
    wire sbe_sel_out_m1_n8 ;
    wire sbe_sel_out_m0_n8 ;
    wire [7:0] O ;
    wire [6:3] sbe_X ;
    wire [7:0] sbe_Z ;
    wire [3:0] sbe_inv_c ;
    wire [1:0] sbe_inv_pmul_pl ;
    wire [1:0] sbe_inv_pmul_ph ;
    wire [1:0] sbe_inv_qmul_pl ;
    wire [1:0] sbe_inv_qmul_ph ;
    wire new_AGEMA_signal_198 ;
    wire new_AGEMA_signal_199 ;
    wire new_AGEMA_signal_200 ;
    wire new_AGEMA_signal_207 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_212 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_218 ;
    wire new_AGEMA_signal_219 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_225 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire new_AGEMA_signal_544 ;
    wire new_AGEMA_signal_545 ;
    wire new_AGEMA_signal_546 ;
    wire new_AGEMA_signal_547 ;
    wire new_AGEMA_signal_548 ;
    wire new_AGEMA_signal_549 ;
    wire new_AGEMA_signal_550 ;
    wire new_AGEMA_signal_551 ;
    wire new_AGEMA_signal_552 ;
    wire new_AGEMA_signal_553 ;
    wire new_AGEMA_signal_554 ;
    wire new_AGEMA_signal_555 ;
    wire new_AGEMA_signal_556 ;
    wire new_AGEMA_signal_557 ;
    wire new_AGEMA_signal_558 ;
    wire new_AGEMA_signal_559 ;
    wire new_AGEMA_signal_560 ;
    wire new_AGEMA_signal_561 ;
    wire new_AGEMA_signal_562 ;
    wire new_AGEMA_signal_563 ;
    wire new_AGEMA_signal_564 ;
    wire new_AGEMA_signal_565 ;
    wire new_AGEMA_signal_566 ;
    wire new_AGEMA_signal_567 ;
    wire new_AGEMA_signal_568 ;
    wire new_AGEMA_signal_569 ;
    wire new_AGEMA_signal_570 ;
    wire new_AGEMA_signal_571 ;
    wire new_AGEMA_signal_572 ;
    wire new_AGEMA_signal_573 ;
    wire new_AGEMA_signal_574 ;
    wire new_AGEMA_signal_575 ;
    wire new_AGEMA_signal_576 ;
    wire new_AGEMA_signal_577 ;
    wire new_AGEMA_signal_578 ;
    wire new_AGEMA_signal_579 ;
    wire new_AGEMA_signal_580 ;
    wire new_AGEMA_signal_581 ;
    wire new_AGEMA_signal_582 ;
    wire new_AGEMA_signal_583 ;
    wire new_AGEMA_signal_584 ;
    wire new_AGEMA_signal_585 ;
    wire new_AGEMA_signal_586 ;
    wire new_AGEMA_signal_587 ;
    wire new_AGEMA_signal_588 ;
    wire new_AGEMA_signal_589 ;
    wire new_AGEMA_signal_590 ;
    wire new_AGEMA_signal_591 ;
    wire new_AGEMA_signal_592 ;
    wire new_AGEMA_signal_593 ;
    wire new_AGEMA_signal_594 ;
    wire new_AGEMA_signal_595 ;
    wire new_AGEMA_signal_596 ;
    wire new_AGEMA_signal_597 ;
    wire new_AGEMA_signal_598 ;
    wire new_AGEMA_signal_599 ;
    wire new_AGEMA_signal_600 ;
    wire new_AGEMA_signal_601 ;
    wire new_AGEMA_signal_602 ;
    wire new_AGEMA_signal_603 ;
    wire new_AGEMA_signal_604 ;
    wire new_AGEMA_signal_605 ;
    wire new_AGEMA_signal_606 ;
    wire new_AGEMA_signal_607 ;
    wire new_AGEMA_signal_608 ;
    wire new_AGEMA_signal_609 ;
    wire new_AGEMA_signal_610 ;
    wire new_AGEMA_signal_611 ;
    wire new_AGEMA_signal_612 ;
    wire new_AGEMA_signal_613 ;
    wire new_AGEMA_signal_614 ;
    wire new_AGEMA_signal_615 ;
    wire new_AGEMA_signal_616 ;
    wire new_AGEMA_signal_617 ;
    wire new_AGEMA_signal_618 ;
    wire new_AGEMA_signal_619 ;
    wire new_AGEMA_signal_620 ;
    wire new_AGEMA_signal_621 ;
    wire new_AGEMA_signal_622 ;
    wire new_AGEMA_signal_623 ;
    wire new_AGEMA_signal_624 ;
    wire new_AGEMA_signal_625 ;
    wire new_AGEMA_signal_626 ;
    wire new_AGEMA_signal_627 ;
    wire new_AGEMA_signal_628 ;
    wire new_AGEMA_signal_629 ;
    wire new_AGEMA_signal_630 ;
    wire new_AGEMA_signal_631 ;
    wire new_AGEMA_signal_632 ;
    wire new_AGEMA_signal_633 ;
    wire new_AGEMA_signal_634 ;
    wire new_AGEMA_signal_635 ;
    wire new_AGEMA_signal_636 ;
    wire new_AGEMA_signal_637 ;
    wire new_AGEMA_signal_638 ;
    wire new_AGEMA_signal_639 ;
    wire new_AGEMA_signal_640 ;
    wire new_AGEMA_signal_641 ;
    wire new_AGEMA_signal_642 ;
    wire new_AGEMA_signal_643 ;
    wire new_AGEMA_signal_644 ;
    wire new_AGEMA_signal_645 ;
    wire new_AGEMA_signal_646 ;
    wire new_AGEMA_signal_647 ;
    wire new_AGEMA_signal_648 ;
    wire new_AGEMA_signal_649 ;
    wire new_AGEMA_signal_650 ;
    wire new_AGEMA_signal_651 ;
    wire new_AGEMA_signal_652 ;
    wire new_AGEMA_signal_653 ;
    wire new_AGEMA_signal_654 ;
    wire new_AGEMA_signal_655 ;
    wire new_AGEMA_signal_656 ;
    wire new_AGEMA_signal_657 ;
    wire new_AGEMA_signal_658 ;
    wire new_AGEMA_signal_659 ;
    wire new_AGEMA_signal_660 ;
    wire new_AGEMA_signal_661 ;
    wire new_AGEMA_signal_662 ;
    wire new_AGEMA_signal_663 ;
    wire new_AGEMA_signal_664 ;
    wire new_AGEMA_signal_665 ;
    wire new_AGEMA_signal_666 ;
    wire new_AGEMA_signal_667 ;
    wire new_AGEMA_signal_668 ;
    wire new_AGEMA_signal_669 ;
    wire new_AGEMA_signal_670 ;
    wire new_AGEMA_signal_671 ;
    wire new_AGEMA_signal_672 ;
    wire new_AGEMA_signal_673 ;
    wire new_AGEMA_signal_674 ;
    wire new_AGEMA_signal_675 ;
    wire new_AGEMA_signal_676 ;
    wire new_AGEMA_signal_677 ;
    wire new_AGEMA_signal_678 ;
    wire new_AGEMA_signal_679 ;
    wire new_AGEMA_signal_680 ;
    wire new_AGEMA_signal_681 ;
    wire new_AGEMA_signal_682 ;
    wire new_AGEMA_signal_683 ;
    wire new_AGEMA_signal_684 ;
    wire new_AGEMA_signal_685 ;
    wire new_AGEMA_signal_686 ;
    wire new_AGEMA_signal_687 ;
    wire new_AGEMA_signal_688 ;
    wire new_AGEMA_signal_689 ;
    wire new_AGEMA_signal_690 ;
    wire new_AGEMA_signal_691 ;
    wire new_AGEMA_signal_692 ;
    wire new_AGEMA_signal_693 ;
    wire new_AGEMA_signal_694 ;
    wire new_AGEMA_signal_695 ;
    wire new_AGEMA_signal_696 ;
    wire new_AGEMA_signal_697 ;
    wire new_AGEMA_signal_698 ;
    wire new_AGEMA_signal_699 ;
    wire new_AGEMA_signal_700 ;
    wire new_AGEMA_signal_701 ;
    wire new_AGEMA_signal_702 ;
    wire new_AGEMA_signal_703 ;
    wire new_AGEMA_signal_704 ;
    wire new_AGEMA_signal_705 ;
    wire new_AGEMA_signal_706 ;
    wire new_AGEMA_signal_707 ;
    wire new_AGEMA_signal_708 ;
    wire new_AGEMA_signal_709 ;
    wire new_AGEMA_signal_710 ;
    wire new_AGEMA_signal_711 ;
    wire new_AGEMA_signal_712 ;
    wire new_AGEMA_signal_713 ;
    wire new_AGEMA_signal_714 ;
    wire new_AGEMA_signal_715 ;
    wire new_AGEMA_signal_716 ;
    wire new_AGEMA_signal_717 ;
    wire new_AGEMA_signal_718 ;
    wire new_AGEMA_signal_719 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U39 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, sbe_n25}), .c ({new_AGEMA_signal_260, new_AGEMA_signal_259, new_AGEMA_signal_258, sbe_n12}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U38 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, sbe_Y_4_}), .c ({new_AGEMA_signal_284, new_AGEMA_signal_283, new_AGEMA_signal_282, sbe_n24}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U37 ( .a ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, sbe_Y_2_}), .b ({new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, sbe_n10}), .c ({new_AGEMA_signal_263, new_AGEMA_signal_262, new_AGEMA_signal_261, sbe_n23}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U36 ( .a ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_n9}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, sbe_n8}), .c ({new_AGEMA_signal_239, new_AGEMA_signal_238, new_AGEMA_signal_237, sbe_n22}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U35 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_212, new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n11}), .c ({new_AGEMA_signal_221, new_AGEMA_signal_220, new_AGEMA_signal_219, sbe_n21}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U29 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, sbe_n10}), .c ({new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_Y_6_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U28 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_200, new_AGEMA_signal_199, new_AGEMA_signal_198, sbe_Y_5_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U27 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, sbe_n10}), .c ({new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, sbe_Y_4_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U26 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_n9}), .c ({new_AGEMA_signal_245, new_AGEMA_signal_244, new_AGEMA_signal_243, sbe_n10}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U25 ( .a ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, sbe_n8}), .c ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, sbe_Y_2_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U24 ( .a ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_209, new_AGEMA_signal_208, new_AGEMA_signal_207, sbe_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U23 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_236, new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_n7}), .c ({new_AGEMA_signal_248, new_AGEMA_signal_247, new_AGEMA_signal_246, sbe_Y_1_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U22 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_272, new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_B_6_}), .c ({new_AGEMA_signal_287, new_AGEMA_signal_286, new_AGEMA_signal_285, sbe_Y_0_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U8 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, sbe_n25}), .c ({new_AGEMA_signal_272, new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_B_6_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U7 ( .a ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_n9}), .c ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, sbe_n25}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U6 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n2}), .c ({new_AGEMA_signal_230, new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_n9}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U5 ( .a ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n3}), .b ({new_AGEMA_signal_212, new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n11}), .c ({new_AGEMA_signal_275, new_AGEMA_signal_274, new_AGEMA_signal_273, sbe_B_3_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U4 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_236, new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_n7}), .c ({new_AGEMA_signal_254, new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n3}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U3 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n2}), .c ({new_AGEMA_signal_236, new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_n7}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U2 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_212, new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n11}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_U1 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m7_U2 ( .a ({new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_sel_in_m7_n8}), .b ({new_AGEMA_signal_308, new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_Z[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_212, new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n11}), .a ({new_AGEMA_signal_263, new_AGEMA_signal_262, new_AGEMA_signal_261, sbe_n23}), .c ({new_AGEMA_signal_290, new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_sel_in_m7_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m6_U2 ( .a ({new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, sbe_sel_in_m6_n8}), .b ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, sbe_Z[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_266, new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_Y_6_}), .a ({new_AGEMA_signal_272, new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_B_6_}), .c ({new_AGEMA_signal_293, new_AGEMA_signal_292, new_AGEMA_signal_291, sbe_sel_in_m6_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m5_U2 ( .a ({new_AGEMA_signal_296, new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_sel_in_m5_n8}), .b ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_Z[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_200, new_AGEMA_signal_199, new_AGEMA_signal_198, sbe_Y_5_}), .a ({new_AGEMA_signal_260, new_AGEMA_signal_259, new_AGEMA_signal_258, sbe_n12}), .c ({new_AGEMA_signal_296, new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_sel_in_m5_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m4_U2 ( .a ({new_AGEMA_signal_299, new_AGEMA_signal_298, new_AGEMA_signal_297, sbe_sel_in_m4_n8}), .b ({new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, sbe_Z[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, new_AGEMA_signal_267, sbe_Y_4_}), .a ({new_AGEMA_signal_239, new_AGEMA_signal_238, new_AGEMA_signal_237, sbe_n22}), .c ({new_AGEMA_signal_299, new_AGEMA_signal_298, new_AGEMA_signal_297, sbe_sel_in_m4_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m3_U2 ( .a ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_sel_in_m3_n8}), .b ({new_AGEMA_signal_320, new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_Z[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_221, new_AGEMA_signal_220, new_AGEMA_signal_219, sbe_n21}), .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, new_AGEMA_signal_273, sbe_B_3_}), .c ({new_AGEMA_signal_302, new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_sel_in_m3_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m2_U2 ( .a ({new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, sbe_sel_in_m2_n8}), .b ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, new_AGEMA_signal_225, sbe_Y_2_}), .a ({new_AGEMA_signal_218, new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n2}), .c ({new_AGEMA_signal_257, new_AGEMA_signal_256, new_AGEMA_signal_255, sbe_sel_in_m2_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m1_U2 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_280, new_AGEMA_signal_279, sbe_sel_in_m1_n8}), .b ({new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, sbe_Z[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_248, new_AGEMA_signal_247, new_AGEMA_signal_246, sbe_Y_1_}), .a ({new_AGEMA_signal_251, new_AGEMA_signal_250, new_AGEMA_signal_249, sbe_n25}), .c ({new_AGEMA_signal_281, new_AGEMA_signal_280, new_AGEMA_signal_279, sbe_sel_in_m1_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m0_U2 ( .a ({new_AGEMA_signal_323, new_AGEMA_signal_322, new_AGEMA_signal_321, sbe_sel_in_m0_n8}), .b ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_Z[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_in_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_287, new_AGEMA_signal_286, new_AGEMA_signal_285, sbe_Y_0_}), .a ({new_AGEMA_signal_284, new_AGEMA_signal_283, new_AGEMA_signal_282, sbe_n24}), .c ({new_AGEMA_signal_323, new_AGEMA_signal_322, new_AGEMA_signal_321, sbe_sel_in_m0_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U10 ( .a ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_Z[0]}), .b ({new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, sbe_Z[1]}), .c ({new_AGEMA_signal_368, new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_bl}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U9 ( .a ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[2]}), .b ({new_AGEMA_signal_320, new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_Z[3]}), .c ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_bh}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U8 ( .a ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, sbe_inv_sb_0_}), .b ({new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, sbe_inv_sb_1_}), .c ({new_AGEMA_signal_392, new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_bb}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U7 ( .a ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_Z[0]}), .b ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[2]}), .c ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, sbe_inv_sb_0_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U6 ( .a ({new_AGEMA_signal_320, new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_Z[3]}), .b ({new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, sbe_Z[1]}), .c ({new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, sbe_inv_sb_1_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U5 ( .a ({new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, sbe_Z[4]}), .b ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_Z[5]}), .c ({new_AGEMA_signal_344, new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_al}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U4 ( .a ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, sbe_Z[6]}), .b ({new_AGEMA_signal_308, new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_Z[7]}), .c ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, sbe_inv_ah}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U3 ( .a ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, sbe_inv_sa_1_}), .c ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_aa}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U2 ( .a ({new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, sbe_Z[4]}), .b ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, sbe_Z[6]}), .c ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_sa_0_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U1 ( .a ({new_AGEMA_signal_308, new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_Z[7]}), .b ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_Z[5]}), .c ({new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, sbe_inv_sa_1_}) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk ( clk ), .rst ( rst ), .GatedClk ( clk_gated ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U34 ( .a ({new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_n21}), .b ({new_AGEMA_signal_395, new_AGEMA_signal_394, new_AGEMA_signal_393, sbe_inv_n20}), .c ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_c[3]}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U33 ( .a ({new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, sbe_inv_n19}), .b ({new_AGEMA_signal_329, new_AGEMA_signal_328, new_AGEMA_signal_327, sbe_inv_n18}), .c ({new_AGEMA_signal_395, new_AGEMA_signal_394, new_AGEMA_signal_393, sbe_inv_n20}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U32 ( .ina ({new_AGEMA_signal_308, new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_Z[7]}), .inb ({new_AGEMA_signal_320, new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_Z[3]}), .clk ( clk ), .rnd ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .outt ({new_AGEMA_signal_329, new_AGEMA_signal_328, new_AGEMA_signal_327, sbe_inv_n18}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U31 ( .ina ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_sa_0_}), .inb ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, sbe_inv_sb_0_}), .clk ( clk ), .rnd ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .outt ({new_AGEMA_signal_377, new_AGEMA_signal_376, new_AGEMA_signal_375, sbe_inv_n19}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U30 ( .a ({new_AGEMA_signal_404, new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_n17}), .b ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, sbe_inv_n16}), .c ({new_AGEMA_signal_410, new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_n21}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U29 ( .a ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_n15}), .b ({new_AGEMA_signal_380, new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_n14}), .c ({new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, sbe_inv_c[2]}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U28 ( .a ({new_AGEMA_signal_356, new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_n13}), .b ({new_AGEMA_signal_332, new_AGEMA_signal_331, new_AGEMA_signal_330, sbe_inv_n12}), .c ({new_AGEMA_signal_380, new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_n14}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U27 ( .ina ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, sbe_Z[6]}), .inb ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[2]}), .clk ( clk ), .rnd ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .outt ({new_AGEMA_signal_332, new_AGEMA_signal_331, new_AGEMA_signal_330, sbe_inv_n12}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U26 ( .ina ({new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, sbe_inv_sa_1_}), .inb ({new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, sbe_inv_sb_1_}), .clk ( clk ), .rnd ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .outt ({new_AGEMA_signal_356, new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_n13}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U25 ( .a ({new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, sbe_inv_n11}), .b ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, sbe_inv_n16}), .c ({new_AGEMA_signal_398, new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_n15}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U24 ( .ina ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, sbe_inv_ah}), .inb ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_bh}), .clk ( clk ), .rnd ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .outt ({new_AGEMA_signal_359, new_AGEMA_signal_358, new_AGEMA_signal_357, sbe_inv_n16}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U23 ( .a ({new_AGEMA_signal_416, new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_n10}), .b ({new_AGEMA_signal_401, new_AGEMA_signal_400, new_AGEMA_signal_399, sbe_inv_n9}), .c ({new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, sbe_inv_c[1]}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U22 ( .a ({new_AGEMA_signal_383, new_AGEMA_signal_382, new_AGEMA_signal_381, sbe_inv_n8}), .b ({new_AGEMA_signal_335, new_AGEMA_signal_334, new_AGEMA_signal_333, sbe_inv_n7}), .c ({new_AGEMA_signal_401, new_AGEMA_signal_400, new_AGEMA_signal_399, sbe_inv_n9}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U21 ( .ina ({new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, sbe_Z[1]}), .inb ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_Z[5]}), .clk ( clk ), .rnd ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .outt ({new_AGEMA_signal_335, new_AGEMA_signal_334, new_AGEMA_signal_333, sbe_inv_n7}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U20 ( .ina ({new_AGEMA_signal_344, new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_al}), .inb ({new_AGEMA_signal_368, new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_bl}), .clk ( clk ), .rnd ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .outt ({new_AGEMA_signal_383, new_AGEMA_signal_382, new_AGEMA_signal_381, sbe_inv_n8}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U19 ( .a ({new_AGEMA_signal_404, new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_n17}), .b ({new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, sbe_inv_n11}), .c ({new_AGEMA_signal_416, new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_n10}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U18 ( .ina ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_aa}), .inb ({new_AGEMA_signal_392, new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_bb}), .clk ( clk ), .rnd ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .outt ({new_AGEMA_signal_404, new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_n17}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U17 ( .a ({new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, sbe_inv_n11}), .b ({new_AGEMA_signal_419, new_AGEMA_signal_418, new_AGEMA_signal_417, sbe_inv_n6}), .c ({new_AGEMA_signal_428, new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_c[0]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U16 ( .a ({new_AGEMA_signal_365, new_AGEMA_signal_364, new_AGEMA_signal_363, sbe_inv_n5}), .b ({new_AGEMA_signal_407, new_AGEMA_signal_406, new_AGEMA_signal_405, sbe_inv_n4}), .c ({new_AGEMA_signal_419, new_AGEMA_signal_418, new_AGEMA_signal_417, sbe_inv_n6}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U15 ( .a ({new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_inv_n3}), .b ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_n2}), .c ({new_AGEMA_signal_407, new_AGEMA_signal_406, new_AGEMA_signal_405, sbe_inv_n4}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U14 ( .ina ({new_AGEMA_signal_344, new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_al}), .inb ({new_AGEMA_signal_368, new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_bl}), .clk ( clk ), .rnd ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .outt ({new_AGEMA_signal_386, new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_n2}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U13 ( .ina ({new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, sbe_Z[4]}), .inb ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_Z[0]}), .clk ( clk ), .rnd ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .outt ({new_AGEMA_signal_362, new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_inv_n3}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U12 ( .ina ({new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, sbe_inv_sb_1_}), .inb ({new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, sbe_inv_sa_1_}), .clk ( clk ), .rnd ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .outt ({new_AGEMA_signal_365, new_AGEMA_signal_364, new_AGEMA_signal_363, sbe_inv_n5}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U11 ( .ina ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_sa_0_}), .inb ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, sbe_inv_sb_0_}), .clk ( clk ), .rnd ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .outt ({new_AGEMA_signal_389, new_AGEMA_signal_388, new_AGEMA_signal_387, sbe_inv_n11}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U2 ( .a ({new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, sbe_inv_c[2]}), .b ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_c[3]}), .c ({new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, sbe_inv_dinv_sa}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U1 ( .a ({new_AGEMA_signal_428, new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_c[0]}), .b ({new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, sbe_inv_c[1]}), .c ({new_AGEMA_signal_440, new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_dinv_sb}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U9 ( .a ({new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_452, new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_dinv_d_1_}), .c ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, sbe_inv_dinv_sd}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U8 ( .a ({new_AGEMA_signal_431, new_AGEMA_signal_430, new_AGEMA_signal_429, sbe_inv_dinv_n4}), .b ({new_AGEMA_signal_443, new_AGEMA_signal_442, new_AGEMA_signal_441, sbe_inv_dinv_n3}), .c ({new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, sbe_inv_dinv_d_0_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U7 ( .ina ({new_AGEMA_signal_440, new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_dinv_sb}), .inb ({new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, sbe_inv_dinv_sa}), .clk ( clk ), .rnd ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .outt ({new_AGEMA_signal_443, new_AGEMA_signal_442, new_AGEMA_signal_441, sbe_inv_dinv_n3}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U6 ( .ina ({new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, sbe_inv_c[1]}), .inb ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_c[3]}), .clk ( clk ), .rnd ({Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130]}), .outt ({new_AGEMA_signal_431, new_AGEMA_signal_430, new_AGEMA_signal_429, sbe_inv_dinv_n4}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U5 ( .a ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_dinv_n2}), .b ({new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_dinv_n1}), .c ({new_AGEMA_signal_452, new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_dinv_d_1_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U4 ( .ina ({new_AGEMA_signal_428, new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_c[0]}), .inb ({new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, sbe_inv_c[2]}), .clk ( clk ), .rnd ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140]}), .outt ({new_AGEMA_signal_434, new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_dinv_n1}) ) ;
    nor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_U3 ( .ina ({new_AGEMA_signal_440, new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_dinv_sb}), .inb ({new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, sbe_inv_dinv_sa}), .clk ( clk ), .rnd ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .outt ({new_AGEMA_signal_446, new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_dinv_n2}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U39 ( .a ({new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, sbe_inv_d_0_}), .b ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_d_1_}), .c ({new_AGEMA_signal_488, new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_inv_dl}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U38 ( .a ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, sbe_inv_d_2_}), .b ({new_AGEMA_signal_476, new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_inv_d_3_}), .c ({new_AGEMA_signal_491, new_AGEMA_signal_490, new_AGEMA_signal_489, sbe_inv_dh}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U37 ( .a ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, sbe_inv_sd_1_}), .c ({new_AGEMA_signal_524, new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_inv_dd}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U36 ( .a ({new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, sbe_inv_d_0_}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, sbe_inv_d_2_}), .c ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_inv_sd_0_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_U35 ( .a ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_d_1_}), .b ({new_AGEMA_signal_476, new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_inv_d_3_}), .c ({new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, sbe_inv_sd_1_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_pmul_U5 ( .a ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_inv_dinv_pmul_n8}), .c ({new_AGEMA_signal_476, new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_inv_d_3_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_pmul_U4 ( .ina ({new_AGEMA_signal_452, new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_dinv_d_1_}), .inb ({new_AGEMA_signal_425, new_AGEMA_signal_424, new_AGEMA_signal_423, sbe_inv_c[1]}), .clk ( clk ), .rnd ({Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .outt ({new_AGEMA_signal_458, new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_inv_dinv_pmul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_pmul_U3 ( .a ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, sbe_inv_dinv_pmul_n7}), .c ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, sbe_inv_d_2_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_pmul_U2 ( .ina ({new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, sbe_inv_dinv_d_0_}), .inb ({new_AGEMA_signal_428, new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_c[0]}), .clk ( clk ), .rnd ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170]}), .outt ({new_AGEMA_signal_461, new_AGEMA_signal_460, new_AGEMA_signal_459, sbe_inv_dinv_pmul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_pmul_U1 ( .ina ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, sbe_inv_dinv_sd}), .inb ({new_AGEMA_signal_440, new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_dinv_sb}), .clk ( clk ), .rnd ({Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .outt ({new_AGEMA_signal_470, new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_inv_dinv_pmul_n9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_qmul_U5 ( .a ({new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_464, new_AGEMA_signal_463, new_AGEMA_signal_462, sbe_inv_dinv_qmul_n8}), .c ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_d_1_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_qmul_U4 ( .ina ({new_AGEMA_signal_452, new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_dinv_d_1_}), .inb ({new_AGEMA_signal_422, new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_c[3]}), .clk ( clk ), .rnd ({Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190]}), .outt ({new_AGEMA_signal_464, new_AGEMA_signal_463, new_AGEMA_signal_462, sbe_inv_dinv_qmul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_qmul_U3 ( .a ({new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_467, new_AGEMA_signal_466, new_AGEMA_signal_465, sbe_inv_dinv_qmul_n7}), .c ({new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, sbe_inv_d_0_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_qmul_U2 ( .ina ({new_AGEMA_signal_449, new_AGEMA_signal_448, new_AGEMA_signal_447, sbe_inv_dinv_d_0_}), .inb ({new_AGEMA_signal_413, new_AGEMA_signal_412, new_AGEMA_signal_411, sbe_inv_c[2]}), .clk ( clk ), .rnd ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200]}), .outt ({new_AGEMA_signal_467, new_AGEMA_signal_466, new_AGEMA_signal_465, sbe_inv_dinv_qmul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_dinv_qmul_U1 ( .ina ({new_AGEMA_signal_455, new_AGEMA_signal_454, new_AGEMA_signal_453, sbe_inv_dinv_sd}), .inb ({new_AGEMA_signal_437, new_AGEMA_signal_436, new_AGEMA_signal_435, sbe_inv_dinv_sa}), .clk ( clk ), .rnd ({Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .outt ({new_AGEMA_signal_473, new_AGEMA_signal_472, new_AGEMA_signal_471, sbe_inv_dinv_qmul_n9}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    not_masked #(.security_order(3), .pipeline(0)) sbe_U40 ( .a ({new_AGEMA_signal_596, new_AGEMA_signal_595, new_AGEMA_signal_594, sbe_C_2_}), .b ({new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, sbe_n1}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U34 ( .a ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, sbe_C_7_}), .b ({new_AGEMA_signal_644, new_AGEMA_signal_643, new_AGEMA_signal_642, sbe_n17}), .c ({new_AGEMA_signal_659, new_AGEMA_signal_658, new_AGEMA_signal_657, sbe_n16}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U33 ( .a ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_C_4_}), .b ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, sbe_n18}), .c ({new_AGEMA_signal_644, new_AGEMA_signal_643, new_AGEMA_signal_642, sbe_n17}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U32 ( .a ({new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, sbe_C_5_}), .b ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, sbe_C_1_}), .c ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, sbe_n18}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U31 ( .a ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, sbe_C_1_}), .b ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_C_4_}), .c ({new_AGEMA_signal_629, new_AGEMA_signal_628, new_AGEMA_signal_627, sbe_n15}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U30 ( .a ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, sbe_C_6_}), .b ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, sbe_C_1_}), .c ({new_AGEMA_signal_632, new_AGEMA_signal_631, new_AGEMA_signal_630, sbe_n14}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U21 ( .a ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, sbe_n6}), .b ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, sbe_C_1_}), .c ({new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, sbe_X[6]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U20 ( .a ({new_AGEMA_signal_596, new_AGEMA_signal_595, new_AGEMA_signal_594, sbe_C_2_}), .b ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, sbe_n6}), .c ({new_AGEMA_signal_689, new_AGEMA_signal_688, new_AGEMA_signal_687, sbe_X[5]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U19 ( .a ({new_AGEMA_signal_608, new_AGEMA_signal_607, new_AGEMA_signal_606, sbe_D_5_}), .b ({new_AGEMA_signal_647, new_AGEMA_signal_646, new_AGEMA_signal_645, sbe_n20}), .c ({new_AGEMA_signal_662, new_AGEMA_signal_661, new_AGEMA_signal_660, sbe_n6}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U18 ( .a ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, sbe_n5}), .b ({new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, sbe_D_0_}), .c ({new_AGEMA_signal_665, new_AGEMA_signal_664, new_AGEMA_signal_663, sbe_X[3]}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U17 ( .a ({new_AGEMA_signal_647, new_AGEMA_signal_646, new_AGEMA_signal_645, sbe_n20}), .b ({new_AGEMA_signal_611, new_AGEMA_signal_610, new_AGEMA_signal_609, sbe_n4}), .c ({new_AGEMA_signal_668, new_AGEMA_signal_667, new_AGEMA_signal_666, sbe_D_3_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U16 ( .a ({new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, sbe_C_5_}), .b ({new_AGEMA_signal_635, new_AGEMA_signal_634, new_AGEMA_signal_633, sbe_D_6_}), .c ({new_AGEMA_signal_647, new_AGEMA_signal_646, new_AGEMA_signal_645, sbe_n20}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U15 ( .a ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, sbe_C_7_}), .b ({new_AGEMA_signal_620, new_AGEMA_signal_619, new_AGEMA_signal_618, sbe_C_3_}), .c ({new_AGEMA_signal_635, new_AGEMA_signal_634, new_AGEMA_signal_633, sbe_D_6_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U14 ( .a ({new_AGEMA_signal_608, new_AGEMA_signal_607, new_AGEMA_signal_606, sbe_D_5_}), .b ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, sbe_n5}), .c ({new_AGEMA_signal_671, new_AGEMA_signal_670, new_AGEMA_signal_669, sbe_D_2_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U13 ( .a ({new_AGEMA_signal_596, new_AGEMA_signal_595, new_AGEMA_signal_594, sbe_C_2_}), .b ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, sbe_n19}), .c ({new_AGEMA_signal_650, new_AGEMA_signal_649, new_AGEMA_signal_648, sbe_n5}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U12 ( .a ({new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, sbe_C_5_}), .b ({new_AGEMA_signal_620, new_AGEMA_signal_619, new_AGEMA_signal_618, sbe_C_3_}), .c ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, sbe_n19}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U11 ( .a ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, sbe_C_6_}), .b ({new_AGEMA_signal_599, new_AGEMA_signal_598, new_AGEMA_signal_597, sbe_C_0_}), .c ({new_AGEMA_signal_608, new_AGEMA_signal_607, new_AGEMA_signal_606, sbe_D_5_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U10 ( .a ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, sbe_C_1_}), .b ({new_AGEMA_signal_611, new_AGEMA_signal_610, new_AGEMA_signal_609, sbe_n4}), .c ({new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, sbe_D_0_}) ) ;
    xnor_HPC1 #(.security_order(3), .pipeline(0)) sbe_U9 ( .a ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, sbe_C_6_}), .b ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_C_4_}), .c ({new_AGEMA_signal_611, new_AGEMA_signal_610, new_AGEMA_signal_609, sbe_n4}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_U4 ( .a ({new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_551, new_AGEMA_signal_550, new_AGEMA_signal_549, sbe_inv_pmul_ph[1]}), .c ({new_AGEMA_signal_614, new_AGEMA_signal_613, new_AGEMA_signal_612, sbe_C_7_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_U3 ( .a ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, sbe_inv_pmul_ph[0]}), .c ({new_AGEMA_signal_587, new_AGEMA_signal_586, new_AGEMA_signal_585, sbe_C_6_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_U2 ( .a ({new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, sbe_inv_pmul_pl[1]}), .c ({new_AGEMA_signal_617, new_AGEMA_signal_616, new_AGEMA_signal_615, sbe_C_5_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_U1 ( .a ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_560, new_AGEMA_signal_559, new_AGEMA_signal_558, sbe_inv_pmul_pl[0]}), .c ({new_AGEMA_signal_590, new_AGEMA_signal_589, new_AGEMA_signal_588, sbe_C_4_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_himul_U5 ( .a ({new_AGEMA_signal_527, new_AGEMA_signal_526, new_AGEMA_signal_525, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_500, new_AGEMA_signal_499, new_AGEMA_signal_498, sbe_inv_pmul_himul_n8}), .c ({new_AGEMA_signal_551, new_AGEMA_signal_550, new_AGEMA_signal_549, sbe_inv_pmul_ph[1]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_himul_U4 ( .ina ({new_AGEMA_signal_476, new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_inv_d_3_}), .inb ({new_AGEMA_signal_320, new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_Z[3]}), .clk ( clk ), .rnd ({Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220]}), .outt ({new_AGEMA_signal_500, new_AGEMA_signal_499, new_AGEMA_signal_498, sbe_inv_pmul_himul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_himul_U3 ( .a ({new_AGEMA_signal_527, new_AGEMA_signal_526, new_AGEMA_signal_525, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_503, new_AGEMA_signal_502, new_AGEMA_signal_501, sbe_inv_pmul_himul_n7}), .c ({new_AGEMA_signal_554, new_AGEMA_signal_553, new_AGEMA_signal_552, sbe_inv_pmul_ph[0]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_himul_U2 ( .ina ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, sbe_inv_d_2_}), .inb ({new_AGEMA_signal_278, new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[2]}), .clk ( clk ), .rnd ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230]}), .outt ({new_AGEMA_signal_503, new_AGEMA_signal_502, new_AGEMA_signal_501, sbe_inv_pmul_himul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_himul_U1 ( .ina ({new_AGEMA_signal_491, new_AGEMA_signal_490, new_AGEMA_signal_489, sbe_inv_dh}), .inb ({new_AGEMA_signal_338, new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_bh}), .clk ( clk ), .rnd ({Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .outt ({new_AGEMA_signal_527, new_AGEMA_signal_526, new_AGEMA_signal_525, sbe_inv_pmul_himul_n9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_lomul_U5 ( .a ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_inv_pmul_lomul_n8}), .c ({new_AGEMA_signal_557, new_AGEMA_signal_556, new_AGEMA_signal_555, sbe_inv_pmul_pl[1]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_lomul_U4 ( .ina ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_d_1_}), .inb ({new_AGEMA_signal_305, new_AGEMA_signal_304, new_AGEMA_signal_303, sbe_Z[1]}), .clk ( clk ), .rnd ({Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250]}), .outt ({new_AGEMA_signal_506, new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_inv_pmul_lomul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_lomul_U3 ( .a ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_509, new_AGEMA_signal_508, new_AGEMA_signal_507, sbe_inv_pmul_lomul_n7}), .c ({new_AGEMA_signal_560, new_AGEMA_signal_559, new_AGEMA_signal_558, sbe_inv_pmul_pl[0]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_lomul_U2 ( .ina ({new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, sbe_inv_d_0_}), .inb ({new_AGEMA_signal_326, new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_Z[0]}), .clk ( clk ), .rnd ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260]}), .outt ({new_AGEMA_signal_509, new_AGEMA_signal_508, new_AGEMA_signal_507, sbe_inv_pmul_lomul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_lomul_U1 ( .ina ({new_AGEMA_signal_488, new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_inv_dl}), .inb ({new_AGEMA_signal_368, new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_bl}), .clk ( clk ), .rnd ({Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .outt ({new_AGEMA_signal_530, new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_inv_pmul_lomul_n9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_summul_U5 ( .a ({new_AGEMA_signal_536, new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_563, new_AGEMA_signal_562, new_AGEMA_signal_561, sbe_inv_pmul_summul_n8}), .c ({new_AGEMA_signal_593, new_AGEMA_signal_592, new_AGEMA_signal_591, sbe_inv_pmul_p_1_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_summul_U4 ( .ina ({new_AGEMA_signal_524, new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_inv_dd}), .inb ({new_AGEMA_signal_392, new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_bb}), .clk ( clk ), .rnd ({Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280]}), .outt ({new_AGEMA_signal_563, new_AGEMA_signal_562, new_AGEMA_signal_561, sbe_inv_pmul_summul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_summul_U3 ( .a ({new_AGEMA_signal_536, new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_533, new_AGEMA_signal_532, new_AGEMA_signal_531, sbe_inv_pmul_summul_n7}), .c ({new_AGEMA_signal_566, new_AGEMA_signal_565, new_AGEMA_signal_564, sbe_inv_pmul_p_0_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_summul_U2 ( .ina ({new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, sbe_inv_sd_1_}), .inb ({new_AGEMA_signal_341, new_AGEMA_signal_340, new_AGEMA_signal_339, sbe_inv_sb_1_}), .clk ( clk ), .rnd ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290]}), .outt ({new_AGEMA_signal_533, new_AGEMA_signal_532, new_AGEMA_signal_531, sbe_inv_pmul_summul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_pmul_summul_U1 ( .ina ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_inv_sd_0_}), .inb ({new_AGEMA_signal_371, new_AGEMA_signal_370, new_AGEMA_signal_369, sbe_inv_sb_0_}), .clk ( clk ), .rnd ({Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .outt ({new_AGEMA_signal_536, new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_inv_pmul_summul_n9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_U4 ( .a ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_569, new_AGEMA_signal_568, new_AGEMA_signal_567, sbe_inv_qmul_ph[1]}), .c ({new_AGEMA_signal_620, new_AGEMA_signal_619, new_AGEMA_signal_618, sbe_C_3_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_U3 ( .a ({new_AGEMA_signal_584, new_AGEMA_signal_583, new_AGEMA_signal_582, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_572, new_AGEMA_signal_571, new_AGEMA_signal_570, sbe_inv_qmul_ph[0]}), .c ({new_AGEMA_signal_596, new_AGEMA_signal_595, new_AGEMA_signal_594, sbe_C_2_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_U2 ( .a ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, sbe_inv_qmul_pl[1]}), .c ({new_AGEMA_signal_623, new_AGEMA_signal_622, new_AGEMA_signal_621, sbe_C_1_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_U1 ( .a ({new_AGEMA_signal_584, new_AGEMA_signal_583, new_AGEMA_signal_582, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_qmul_pl[0]}), .c ({new_AGEMA_signal_599, new_AGEMA_signal_598, new_AGEMA_signal_597, sbe_C_0_}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_himul_U5 ( .a ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_512, new_AGEMA_signal_511, new_AGEMA_signal_510, sbe_inv_qmul_himul_n8}), .c ({new_AGEMA_signal_569, new_AGEMA_signal_568, new_AGEMA_signal_567, sbe_inv_qmul_ph[1]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_himul_U4 ( .ina ({new_AGEMA_signal_476, new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_inv_d_3_}), .inb ({new_AGEMA_signal_308, new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_Z[7]}), .clk ( clk ), .rnd ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310]}), .outt ({new_AGEMA_signal_512, new_AGEMA_signal_511, new_AGEMA_signal_510, sbe_inv_qmul_himul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_himul_U3 ( .a ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_515, new_AGEMA_signal_514, new_AGEMA_signal_513, sbe_inv_qmul_himul_n7}), .c ({new_AGEMA_signal_572, new_AGEMA_signal_571, new_AGEMA_signal_570, sbe_inv_qmul_ph[0]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_himul_U2 ( .ina ({new_AGEMA_signal_479, new_AGEMA_signal_478, new_AGEMA_signal_477, sbe_inv_d_2_}), .inb ({new_AGEMA_signal_311, new_AGEMA_signal_310, new_AGEMA_signal_309, sbe_Z[6]}), .clk ( clk ), .rnd ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .outt ({new_AGEMA_signal_515, new_AGEMA_signal_514, new_AGEMA_signal_513, sbe_inv_qmul_himul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_himul_U1 ( .ina ({new_AGEMA_signal_491, new_AGEMA_signal_490, new_AGEMA_signal_489, sbe_inv_dh}), .inb ({new_AGEMA_signal_347, new_AGEMA_signal_346, new_AGEMA_signal_345, sbe_inv_ah}), .clk ( clk ), .rnd ({Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .outt ({new_AGEMA_signal_539, new_AGEMA_signal_538, new_AGEMA_signal_537, sbe_inv_qmul_himul_n9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_lomul_U5 ( .a ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_inv_qmul_lomul_n8}), .c ({new_AGEMA_signal_575, new_AGEMA_signal_574, new_AGEMA_signal_573, sbe_inv_qmul_pl[1]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_lomul_U4 ( .ina ({new_AGEMA_signal_482, new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_inv_d_1_}), .inb ({new_AGEMA_signal_314, new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_Z[5]}), .clk ( clk ), .rnd ({Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340]}), .outt ({new_AGEMA_signal_518, new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_inv_qmul_lomul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_lomul_U3 ( .a ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, sbe_inv_qmul_lomul_n7}), .c ({new_AGEMA_signal_578, new_AGEMA_signal_577, new_AGEMA_signal_576, sbe_inv_qmul_pl[0]}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_lomul_U2 ( .ina ({new_AGEMA_signal_485, new_AGEMA_signal_484, new_AGEMA_signal_483, sbe_inv_d_0_}), .inb ({new_AGEMA_signal_317, new_AGEMA_signal_316, new_AGEMA_signal_315, sbe_Z[4]}), .clk ( clk ), .rnd ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350]}), .outt ({new_AGEMA_signal_521, new_AGEMA_signal_520, new_AGEMA_signal_519, sbe_inv_qmul_lomul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_lomul_U1 ( .ina ({new_AGEMA_signal_488, new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_inv_dl}), .inb ({new_AGEMA_signal_344, new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_al}), .clk ( clk ), .rnd ({Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .outt ({new_AGEMA_signal_542, new_AGEMA_signal_541, new_AGEMA_signal_540, sbe_inv_qmul_lomul_n9}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_summul_U5 ( .a ({new_AGEMA_signal_548, new_AGEMA_signal_547, new_AGEMA_signal_546, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_581, new_AGEMA_signal_580, new_AGEMA_signal_579, sbe_inv_qmul_summul_n8}), .c ({new_AGEMA_signal_602, new_AGEMA_signal_601, new_AGEMA_signal_600, sbe_inv_qmul_p_1_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_summul_U4 ( .ina ({new_AGEMA_signal_524, new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_inv_dd}), .inb ({new_AGEMA_signal_374, new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_aa}), .clk ( clk ), .rnd ({Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370]}), .outt ({new_AGEMA_signal_581, new_AGEMA_signal_580, new_AGEMA_signal_579, sbe_inv_qmul_summul_n8}) ) ;
    xor_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_summul_U3 ( .a ({new_AGEMA_signal_548, new_AGEMA_signal_547, new_AGEMA_signal_546, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_545, new_AGEMA_signal_544, new_AGEMA_signal_543, sbe_inv_qmul_summul_n7}), .c ({new_AGEMA_signal_584, new_AGEMA_signal_583, new_AGEMA_signal_582, sbe_inv_qmul_p_0_}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_summul_U2 ( .ina ({new_AGEMA_signal_497, new_AGEMA_signal_496, new_AGEMA_signal_495, sbe_inv_sd_1_}), .inb ({new_AGEMA_signal_353, new_AGEMA_signal_352, new_AGEMA_signal_351, sbe_inv_sa_1_}), .clk ( clk ), .rnd ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380]}), .outt ({new_AGEMA_signal_545, new_AGEMA_signal_544, new_AGEMA_signal_543, sbe_inv_qmul_summul_n7}) ) ;
    nand_HPC1 #(.security_order(3), .pipeline(0)) sbe_inv_qmul_summul_U1 ( .ina ({new_AGEMA_signal_494, new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_inv_sd_0_}), .inb ({new_AGEMA_signal_350, new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_sa_0_}), .clk ( clk ), .rnd ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .outt ({new_AGEMA_signal_548, new_AGEMA_signal_547, new_AGEMA_signal_546, sbe_inv_qmul_summul_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m7_U2 ( .a ({new_AGEMA_signal_653, new_AGEMA_signal_652, new_AGEMA_signal_651, sbe_sel_out_m7_n8}), .b ({new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, O[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_629, new_AGEMA_signal_628, new_AGEMA_signal_627, sbe_n15}), .a ({new_AGEMA_signal_638, new_AGEMA_signal_637, new_AGEMA_signal_636, sbe_n19}), .c ({new_AGEMA_signal_653, new_AGEMA_signal_652, new_AGEMA_signal_651, sbe_sel_out_m7_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m6_U2 ( .a ({new_AGEMA_signal_704, new_AGEMA_signal_703, new_AGEMA_signal_702, sbe_sel_out_m6_n8}), .b ({new_AGEMA_signal_716, new_AGEMA_signal_715, new_AGEMA_signal_714, O[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_686, new_AGEMA_signal_685, new_AGEMA_signal_684, sbe_X[6]}), .a ({new_AGEMA_signal_635, new_AGEMA_signal_634, new_AGEMA_signal_633, sbe_D_6_}), .c ({new_AGEMA_signal_704, new_AGEMA_signal_703, new_AGEMA_signal_702, sbe_sel_out_m6_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m5_U2 ( .a ({new_AGEMA_signal_707, new_AGEMA_signal_706, new_AGEMA_signal_705, sbe_sel_out_m5_n8}), .b ({new_AGEMA_signal_719, new_AGEMA_signal_718, new_AGEMA_signal_717, O[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_689, new_AGEMA_signal_688, new_AGEMA_signal_687, sbe_X[5]}), .a ({new_AGEMA_signal_608, new_AGEMA_signal_607, new_AGEMA_signal_606, sbe_D_5_}), .c ({new_AGEMA_signal_707, new_AGEMA_signal_706, new_AGEMA_signal_705, sbe_sel_out_m5_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m4_U2 ( .a ({new_AGEMA_signal_677, new_AGEMA_signal_676, new_AGEMA_signal_675, sbe_sel_out_m4_n8}), .b ({new_AGEMA_signal_692, new_AGEMA_signal_691, new_AGEMA_signal_690, O[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_632, new_AGEMA_signal_631, new_AGEMA_signal_630, sbe_n14}), .a ({new_AGEMA_signal_647, new_AGEMA_signal_646, new_AGEMA_signal_645, sbe_n20}), .c ({new_AGEMA_signal_677, new_AGEMA_signal_676, new_AGEMA_signal_675, sbe_sel_out_m4_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m3_U2 ( .a ({new_AGEMA_signal_695, new_AGEMA_signal_694, new_AGEMA_signal_693, sbe_sel_out_m3_n8}), .b ({new_AGEMA_signal_710, new_AGEMA_signal_709, new_AGEMA_signal_708, O[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_665, new_AGEMA_signal_664, new_AGEMA_signal_663, sbe_X[3]}), .a ({new_AGEMA_signal_668, new_AGEMA_signal_667, new_AGEMA_signal_666, sbe_D_3_}), .c ({new_AGEMA_signal_695, new_AGEMA_signal_694, new_AGEMA_signal_693, sbe_sel_out_m3_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m2_U2 ( .a ({new_AGEMA_signal_698, new_AGEMA_signal_697, new_AGEMA_signal_696, sbe_sel_out_m2_n8}), .b ({new_AGEMA_signal_713, new_AGEMA_signal_712, new_AGEMA_signal_711, O[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_659, new_AGEMA_signal_658, new_AGEMA_signal_657, sbe_n16}), .a ({new_AGEMA_signal_671, new_AGEMA_signal_670, new_AGEMA_signal_669, sbe_D_2_}), .c ({new_AGEMA_signal_698, new_AGEMA_signal_697, new_AGEMA_signal_696, sbe_sel_out_m2_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m1_U2 ( .a ({new_AGEMA_signal_680, new_AGEMA_signal_679, new_AGEMA_signal_678, sbe_sel_out_m1_n8}), .b ({new_AGEMA_signal_701, new_AGEMA_signal_700, new_AGEMA_signal_699, O[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_626, new_AGEMA_signal_625, new_AGEMA_signal_624, sbe_n18}), .a ({new_AGEMA_signal_644, new_AGEMA_signal_643, new_AGEMA_signal_642, sbe_n17}), .c ({new_AGEMA_signal_680, new_AGEMA_signal_679, new_AGEMA_signal_678, sbe_sel_out_m1_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m0_U2 ( .a ({new_AGEMA_signal_656, new_AGEMA_signal_655, new_AGEMA_signal_654, sbe_sel_out_m0_n8}), .b ({new_AGEMA_signal_683, new_AGEMA_signal_682, new_AGEMA_signal_681, O[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) sbe_sel_out_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_605, new_AGEMA_signal_604, new_AGEMA_signal_603, sbe_n1}), .a ({new_AGEMA_signal_641, new_AGEMA_signal_640, new_AGEMA_signal_639, sbe_D_0_}), .c ({new_AGEMA_signal_656, new_AGEMA_signal_655, new_AGEMA_signal_654, sbe_sel_out_m0_n8}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_7_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_674, new_AGEMA_signal_673, new_AGEMA_signal_672, O[7]}), .Q ({Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_6_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_716, new_AGEMA_signal_715, new_AGEMA_signal_714, O[6]}), .Q ({Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_5_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_719, new_AGEMA_signal_718, new_AGEMA_signal_717, O[5]}), .Q ({Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_4_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_692, new_AGEMA_signal_691, new_AGEMA_signal_690, O[4]}), .Q ({Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_3_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_710, new_AGEMA_signal_709, new_AGEMA_signal_708, O[3]}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_2_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_713, new_AGEMA_signal_712, new_AGEMA_signal_711, O[2]}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_1_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_701, new_AGEMA_signal_700, new_AGEMA_signal_699, O[1]}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) Y_reg_0_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_683, new_AGEMA_signal_682, new_AGEMA_signal_681, O[0]}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
