/* modified netlist. Source: module PRESENT in file /PRESENT_nibble-serial/AGEMA/PRESENT.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module PRESENT_GHPC_ANF_Pipeline_d1 (data_in_s0, key_s0, clk, reset, data_in_s1, key_s1, Fresh, data_out_s0, done, data_out_s1);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input [63:0] data_in_s1 ;
    input [79:0] key_s1 ;
    input [3:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_443 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_867 ;
    wire signal_870 ;
    wire signal_873 ;
    wire signal_876 ;
    wire signal_879 ;
    wire signal_882 ;
    wire signal_885 ;
    wire signal_888 ;
    wire signal_891 ;
    wire signal_894 ;
    wire signal_897 ;
    wire signal_900 ;
    wire signal_903 ;
    wire signal_906 ;
    wire signal_909 ;
    wire signal_912 ;
    wire signal_914 ;
    wire signal_917 ;
    wire signal_920 ;
    wire signal_923 ;
    wire signal_926 ;
    wire signal_929 ;
    wire signal_932 ;
    wire signal_935 ;
    wire signal_938 ;
    wire signal_941 ;
    wire signal_944 ;
    wire signal_947 ;
    wire signal_950 ;
    wire signal_953 ;
    wire signal_956 ;
    wire signal_959 ;
    wire signal_961 ;
    wire signal_964 ;
    wire signal_967 ;
    wire signal_970 ;
    wire signal_973 ;
    wire signal_976 ;
    wire signal_979 ;
    wire signal_982 ;
    wire signal_985 ;
    wire signal_988 ;
    wire signal_991 ;
    wire signal_994 ;
    wire signal_997 ;
    wire signal_1000 ;
    wire signal_1003 ;
    wire signal_1006 ;
    wire signal_1008 ;
    wire signal_1011 ;
    wire signal_1014 ;
    wire signal_1017 ;
    wire signal_1020 ;
    wire signal_1023 ;
    wire signal_1026 ;
    wire signal_1029 ;
    wire signal_1032 ;
    wire signal_1035 ;
    wire signal_1038 ;
    wire signal_1041 ;
    wire signal_1044 ;
    wire signal_1047 ;
    wire signal_1050 ;
    wire signal_1053 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1279 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1310 ;
    wire signal_1312 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;

    /* cells in depth 0 */
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_0 ( .a ({signal_856, signal_474}), .b ({data_out_s1[60], data_out_s0[60]}), .c ({signal_858, signal_485}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_1 ( .a ({signal_859, signal_473}), .b ({data_out_s1[61], data_out_s0[61]}), .c ({signal_861, signal_484}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_2 ( .a ({signal_862, signal_472}), .b ({data_out_s1[62], data_out_s0[62]}), .c ({signal_864, signal_483}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_3 ( .a ({signal_865, signal_471}), .b ({data_out_s1[63], data_out_s0[63]}), .c ({signal_867, signal_482}) ) ;
    NOR2_X1 cell_4 ( .A1 (reset), .A2 (signal_220), .ZN (signal_236) ) ;
    NOR2_X1 cell_5 ( .A1 (signal_221), .A2 (done), .ZN (signal_220) ) ;
    NOR2_X1 cell_6 ( .A1 (reset), .A2 (signal_222), .ZN (signal_233) ) ;
    NOR2_X1 cell_7 ( .A1 (signal_235), .A2 (signal_223), .ZN (signal_222) ) ;
    NOR2_X1 cell_8 ( .A1 (signal_224), .A2 (signal_225), .ZN (signal_223) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_459), .A2 (signal_461), .ZN (signal_225) ) ;
    OR2_X1 cell_10 ( .A1 (signal_226), .A2 (signal_227), .ZN (signal_224) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_462), .A2 (signal_458), .ZN (signal_227) ) ;
    NAND2_X1 cell_12 ( .A1 (signal_460), .A2 (signal_234), .ZN (signal_226) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_237), .A2 (signal_232), .ZN (done) ) ;
    AND2_X1 cell_14 ( .A1 (signal_221), .A2 (signal_232), .ZN (signal_239) ) ;
    AND2_X1 cell_15 ( .A1 (signal_487), .A2 (signal_228), .ZN (signal_221) ) ;
    NOR2_X1 cell_16 ( .A1 (signal_229), .A2 (signal_230), .ZN (signal_228) ) ;
    NAND2_X1 cell_17 ( .A1 (signal_488), .A2 (signal_489), .ZN (signal_230) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_237), .A2 (signal_486), .ZN (signal_229) ) ;
    NOR2_X1 cell_19 ( .A1 (signal_234), .A2 (signal_232), .ZN (signal_219) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_235), .A2 (signal_237), .ZN (signal_217) ) ;
    NOR2_X1 cell_21 ( .A1 (reset), .A2 (signal_217), .ZN (signal_238) ) ;
    INV_X1 cell_22 ( .A (reset), .ZN (signal_231) ) ;
    INV_X1 cell_23 ( .A (signal_238), .ZN (signal_218) ) ;
    NAND2_X1 cell_24 ( .A1 (signal_240), .A2 (signal_241), .ZN (signal_266) ) ;
    NAND2_X1 cell_25 ( .A1 (signal_242), .A2 (signal_461), .ZN (signal_241) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_243), .A2 (signal_265), .ZN (signal_240) ) ;
    NAND2_X1 cell_27 ( .A1 (signal_244), .A2 (signal_462), .ZN (signal_243) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_245), .A2 (signal_246), .ZN (signal_269) ) ;
    NAND2_X1 cell_29 ( .A1 (signal_247), .A2 (signal_462), .ZN (signal_246) ) ;
    MUX2_X1 cell_30 ( .S (signal_263), .A (signal_248), .B (signal_249), .Z (signal_270) ) ;
    NAND2_X1 cell_31 ( .A1 (signal_242), .A2 (signal_250), .ZN (signal_248) ) ;
    NAND2_X1 cell_32 ( .A1 (signal_244), .A2 (signal_265), .ZN (signal_250) ) ;
    NOR2_X1 cell_33 ( .A1 (signal_251), .A2 (signal_247), .ZN (signal_242) ) ;
    NOR2_X1 cell_34 ( .A1 (signal_239), .A2 (signal_262), .ZN (signal_247) ) ;
    INV_X1 cell_35 ( .A (signal_245), .ZN (signal_251) ) ;
    NAND2_X1 cell_36 ( .A1 (signal_244), .A2 (signal_264), .ZN (signal_245) ) ;
    MUX2_X1 cell_37 ( .S (signal_458), .A (signal_252), .B (signal_253), .Z (signal_271) ) ;
    NAND2_X1 cell_38 ( .A1 (signal_254), .A2 (signal_255), .ZN (signal_253) ) ;
    NAND2_X1 cell_39 ( .A1 (signal_244), .A2 (signal_267), .ZN (signal_254) ) ;
    INV_X1 cell_40 ( .A (signal_256), .ZN (signal_244) ) ;
    NOR2_X1 cell_41 ( .A1 (signal_267), .A2 (signal_257), .ZN (signal_252) ) ;
    INV_X1 cell_42 ( .A (signal_258), .ZN (signal_268) ) ;
    MUX2_X1 cell_43 ( .S (signal_267), .A (signal_255), .B (signal_257), .Z (signal_258) ) ;
    NAND2_X1 cell_44 ( .A1 (signal_460), .A2 (signal_249), .ZN (signal_257) ) ;
    NOR2_X1 cell_45 ( .A1 (signal_256), .A2 (signal_259), .ZN (signal_249) ) ;
    NAND2_X1 cell_46 ( .A1 (signal_239), .A2 (signal_231), .ZN (signal_256) ) ;
    NAND2_X1 cell_47 ( .A1 (signal_231), .A2 (signal_260), .ZN (signal_255) ) ;
    NAND2_X1 cell_48 ( .A1 (signal_239), .A2 (signal_261), .ZN (signal_260) ) ;
    NOR2_X1 cell_49 ( .A1 (signal_263), .A2 (signal_259), .ZN (signal_261) ) ;
    OR2_X1 cell_50 ( .A1 (signal_265), .A2 (signal_264), .ZN (signal_259) ) ;
    INV_X1 cell_51 ( .A (signal_231), .ZN (signal_262) ) ;
    INV_X1 cell_54 ( .A (signal_460), .ZN (signal_263) ) ;
    INV_X1 cell_56 ( .A (signal_462), .ZN (signal_264) ) ;
    INV_X1 cell_58 ( .A (signal_459), .ZN (signal_267) ) ;
    INV_X1 cell_60 ( .A (signal_265), .ZN (signal_461) ) ;
    NOR2_X1 cell_62 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_284) ) ;
    XNOR2_X1 cell_63 ( .A (signal_237), .B (signal_489), .ZN (signal_273) ) ;
    NOR2_X1 cell_64 ( .A1 (signal_274), .A2 (signal_275), .ZN (signal_282) ) ;
    XOR2_X1 cell_65 ( .A (signal_488), .B (signal_276), .Z (signal_275) ) ;
    NOR2_X1 cell_66 ( .A1 (signal_274), .A2 (signal_277), .ZN (signal_283) ) ;
    XOR2_X1 cell_67 ( .A (signal_486), .B (signal_278), .Z (signal_277) ) ;
    NAND2_X1 cell_68 ( .A1 (signal_279), .A2 (signal_487), .ZN (signal_278) ) ;
    NOR2_X1 cell_69 ( .A1 (signal_280), .A2 (signal_274), .ZN (signal_285) ) ;
    INV_X1 cell_70 ( .A (signal_238), .ZN (signal_274) ) ;
    XNOR2_X1 cell_71 ( .A (signal_279), .B (signal_487), .ZN (signal_280) ) ;
    NOR2_X1 cell_72 ( .A1 (signal_281), .A2 (signal_276), .ZN (signal_279) ) ;
    NAND2_X1 cell_73 ( .A1 (signal_237), .A2 (signal_489), .ZN (signal_276) ) ;
    INV_X1 cell_80 ( .A (signal_488), .ZN (signal_281) ) ;
    INV_X1 cell_82 ( .A (signal_234), .ZN (signal_237) ) ;
    INV_X1 cell_84 ( .A (signal_235), .ZN (signal_232) ) ;
    INV_X1 cell_86 ( .A (signal_289), .ZN (signal_290) ) ;
    INV_X1 cell_87 ( .A (signal_289), .ZN (signal_291) ) ;
    INV_X1 cell_88 ( .A (signal_218), .ZN (signal_289) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_109 ( .s (signal_218), .b ({data_out_s1[0], data_out_s0[0]}), .a ({signal_882, signal_549}), .c ({signal_1293, signal_561}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_110 ( .s (signal_218), .b ({data_out_s1[1], data_out_s0[1]}), .a ({signal_885, signal_548}), .c ({signal_1294, signal_560}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_111 ( .s (signal_218), .b ({data_out_s1[2], data_out_s0[2]}), .a ({signal_888, signal_547}), .c ({signal_1295, signal_559}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_112 ( .s (signal_218), .b ({data_out_s1[3], data_out_s0[3]}), .a ({signal_891, signal_546}), .c ({signal_1296, signal_558}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_121 ( .s (signal_290), .b ({data_out_s1[4], data_out_s0[4]}), .a ({signal_894, signal_545}), .c ({signal_1322, signal_565}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_122 ( .s (signal_290), .b ({data_out_s1[5], data_out_s0[5]}), .a ({signal_897, signal_544}), .c ({signal_1323, signal_564}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_123 ( .s (signal_290), .b ({data_out_s1[6], data_out_s0[6]}), .a ({signal_900, signal_543}), .c ({signal_1324, signal_563}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_124 ( .s (signal_290), .b ({data_out_s1[7], data_out_s0[7]}), .a ({signal_903, signal_542}), .c ({signal_1325, signal_562}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_133 ( .s (signal_290), .b ({data_out_s1[8], data_out_s0[8]}), .a ({signal_906, signal_541}), .c ({signal_1326, signal_569}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_134 ( .s (signal_290), .b ({data_out_s1[9], data_out_s0[9]}), .a ({signal_909, signal_540}), .c ({signal_1327, signal_568}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_135 ( .s (signal_290), .b ({data_out_s1[10], data_out_s0[10]}), .a ({signal_912, signal_539}), .c ({signal_1328, signal_567}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_136 ( .s (signal_290), .b ({data_out_s1[11], data_out_s0[11]}), .a ({signal_914, signal_538}), .c ({signal_1329, signal_566}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_145 ( .s (signal_290), .b ({data_out_s1[12], data_out_s0[12]}), .a ({signal_917, signal_537}), .c ({signal_1330, signal_573}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_146 ( .s (signal_290), .b ({data_out_s1[13], data_out_s0[13]}), .a ({signal_920, signal_536}), .c ({signal_1331, signal_572}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_147 ( .s (signal_290), .b ({data_out_s1[14], data_out_s0[14]}), .a ({signal_923, signal_535}), .c ({signal_1332, signal_571}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_148 ( .s (signal_290), .b ({data_out_s1[15], data_out_s0[15]}), .a ({signal_926, signal_534}), .c ({signal_1333, signal_570}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_157 ( .s (signal_290), .b ({data_out_s1[16], data_out_s0[16]}), .a ({signal_929, signal_533}), .c ({signal_1334, signal_577}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_158 ( .s (signal_290), .b ({data_out_s1[17], data_out_s0[17]}), .a ({signal_932, signal_532}), .c ({signal_1335, signal_576}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_159 ( .s (signal_290), .b ({data_out_s1[18], data_out_s0[18]}), .a ({signal_935, signal_531}), .c ({signal_1336, signal_575}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_160 ( .s (signal_290), .b ({data_out_s1[19], data_out_s0[19]}), .a ({signal_938, signal_530}), .c ({signal_1337, signal_574}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_169 ( .s (signal_290), .b ({data_out_s1[20], data_out_s0[20]}), .a ({signal_941, signal_529}), .c ({signal_1338, signal_581}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_170 ( .s (signal_290), .b ({data_out_s1[21], data_out_s0[21]}), .a ({signal_944, signal_528}), .c ({signal_1339, signal_580}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_171 ( .s (signal_290), .b ({data_out_s1[22], data_out_s0[22]}), .a ({signal_947, signal_527}), .c ({signal_1340, signal_579}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_172 ( .s (signal_290), .b ({data_out_s1[23], data_out_s0[23]}), .a ({signal_950, signal_526}), .c ({signal_1341, signal_578}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_181 ( .s (signal_290), .b ({data_out_s1[24], data_out_s0[24]}), .a ({signal_953, signal_525}), .c ({signal_1342, signal_585}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_182 ( .s (signal_290), .b ({data_out_s1[25], data_out_s0[25]}), .a ({signal_956, signal_524}), .c ({signal_1343, signal_584}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_183 ( .s (signal_290), .b ({data_out_s1[26], data_out_s0[26]}), .a ({signal_959, signal_523}), .c ({signal_1344, signal_583}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_184 ( .s (signal_290), .b ({data_out_s1[27], data_out_s0[27]}), .a ({signal_961, signal_522}), .c ({signal_1345, signal_582}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_193 ( .s (signal_290), .b ({data_out_s1[28], data_out_s0[28]}), .a ({signal_964, signal_521}), .c ({signal_1346, signal_589}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_194 ( .s (signal_290), .b ({data_out_s1[29], data_out_s0[29]}), .a ({signal_967, signal_520}), .c ({signal_1347, signal_588}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_195 ( .s (signal_290), .b ({data_out_s1[30], data_out_s0[30]}), .a ({signal_970, signal_519}), .c ({signal_1348, signal_587}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_196 ( .s (signal_290), .b ({data_out_s1[31], data_out_s0[31]}), .a ({signal_973, signal_518}), .c ({signal_1349, signal_586}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_205 ( .s (signal_291), .b ({data_out_s1[32], data_out_s0[32]}), .a ({signal_976, signal_517}), .c ({signal_1350, signal_593}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_206 ( .s (signal_291), .b ({data_out_s1[33], data_out_s0[33]}), .a ({signal_979, signal_516}), .c ({signal_1351, signal_592}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_207 ( .s (signal_291), .b ({data_out_s1[34], data_out_s0[34]}), .a ({signal_982, signal_515}), .c ({signal_1352, signal_591}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_208 ( .s (signal_291), .b ({data_out_s1[35], data_out_s0[35]}), .a ({signal_985, signal_514}), .c ({signal_1353, signal_590}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_217 ( .s (signal_291), .b ({data_out_s1[36], data_out_s0[36]}), .a ({signal_988, signal_513}), .c ({signal_1354, signal_597}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_218 ( .s (signal_291), .b ({data_out_s1[37], data_out_s0[37]}), .a ({signal_991, signal_512}), .c ({signal_1355, signal_596}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_219 ( .s (signal_291), .b ({data_out_s1[38], data_out_s0[38]}), .a ({signal_994, signal_511}), .c ({signal_1356, signal_595}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_220 ( .s (signal_291), .b ({data_out_s1[39], data_out_s0[39]}), .a ({signal_997, signal_510}), .c ({signal_1357, signal_594}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_229 ( .s (signal_291), .b ({data_out_s1[40], data_out_s0[40]}), .a ({signal_1000, signal_509}), .c ({signal_1358, signal_601}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_230 ( .s (signal_291), .b ({data_out_s1[41], data_out_s0[41]}), .a ({signal_1003, signal_508}), .c ({signal_1359, signal_600}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_231 ( .s (signal_291), .b ({data_out_s1[42], data_out_s0[42]}), .a ({signal_1006, signal_507}), .c ({signal_1360, signal_599}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_232 ( .s (signal_291), .b ({data_out_s1[43], data_out_s0[43]}), .a ({signal_1008, signal_506}), .c ({signal_1361, signal_598}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_241 ( .s (signal_291), .b ({data_out_s1[44], data_out_s0[44]}), .a ({signal_1011, signal_505}), .c ({signal_1362, signal_605}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_242 ( .s (signal_291), .b ({data_out_s1[45], data_out_s0[45]}), .a ({signal_1014, signal_504}), .c ({signal_1363, signal_604}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_243 ( .s (signal_291), .b ({data_out_s1[46], data_out_s0[46]}), .a ({signal_1017, signal_503}), .c ({signal_1364, signal_603}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_244 ( .s (signal_291), .b ({data_out_s1[47], data_out_s0[47]}), .a ({signal_1020, signal_502}), .c ({signal_1365, signal_602}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_253 ( .s (signal_291), .b ({data_out_s1[48], data_out_s0[48]}), .a ({signal_1023, signal_501}), .c ({signal_1366, signal_609}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_254 ( .s (signal_291), .b ({data_out_s1[49], data_out_s0[49]}), .a ({signal_1026, signal_500}), .c ({signal_1367, signal_608}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_255 ( .s (signal_291), .b ({data_out_s1[50], data_out_s0[50]}), .a ({signal_1029, signal_499}), .c ({signal_1368, signal_607}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_256 ( .s (signal_291), .b ({data_out_s1[51], data_out_s0[51]}), .a ({signal_1032, signal_498}), .c ({signal_1369, signal_606}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_265 ( .s (signal_291), .b ({data_out_s1[52], data_out_s0[52]}), .a ({signal_1035, signal_497}), .c ({signal_1370, signal_613}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_266 ( .s (signal_291), .b ({data_out_s1[53], data_out_s0[53]}), .a ({signal_1038, signal_496}), .c ({signal_1371, signal_612}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_267 ( .s (signal_291), .b ({data_out_s1[54], data_out_s0[54]}), .a ({signal_1041, signal_495}), .c ({signal_1372, signal_611}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_268 ( .s (signal_291), .b ({data_out_s1[55], data_out_s0[55]}), .a ({signal_1044, signal_494}), .c ({signal_1373, signal_610}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_277 ( .s (signal_291), .b ({data_out_s1[56], data_out_s0[56]}), .a ({signal_1047, signal_493}), .c ({signal_1374, signal_617}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_278 ( .s (signal_291), .b ({data_out_s1[57], data_out_s0[57]}), .a ({signal_1050, signal_492}), .c ({signal_1375, signal_616}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_279 ( .s (signal_291), .b ({data_out_s1[58], data_out_s0[58]}), .a ({signal_1053, signal_491}), .c ({signal_1376, signal_615}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_280 ( .s (signal_291), .b ({data_out_s1[59], data_out_s0[59]}), .a ({signal_1055, signal_490}), .c ({signal_1377, signal_614}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_281 ( .s (reset), .b ({data_out_s1[0], data_out_s0[0]}), .a ({data_in_s1[0], data_in_s0[0]}), .c ({signal_870, signal_553}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_282 ( .s (reset), .b ({data_out_s1[4], data_out_s0[4]}), .a ({data_in_s1[1], data_in_s0[1]}), .c ({signal_873, signal_552}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_283 ( .s (reset), .b ({data_out_s1[8], data_out_s0[8]}), .a ({data_in_s1[2], data_in_s0[2]}), .c ({signal_876, signal_551}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_284 ( .s (reset), .b ({data_out_s1[12], data_out_s0[12]}), .a ({data_in_s1[3], data_in_s0[3]}), .c ({signal_879, signal_550}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_285 ( .s (reset), .b ({data_out_s1[16], data_out_s0[16]}), .a ({data_in_s1[4], data_in_s0[4]}), .c ({signal_882, signal_549}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_286 ( .s (reset), .b ({data_out_s1[20], data_out_s0[20]}), .a ({data_in_s1[5], data_in_s0[5]}), .c ({signal_885, signal_548}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_287 ( .s (reset), .b ({data_out_s1[24], data_out_s0[24]}), .a ({data_in_s1[6], data_in_s0[6]}), .c ({signal_888, signal_547}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_288 ( .s (reset), .b ({data_out_s1[28], data_out_s0[28]}), .a ({data_in_s1[7], data_in_s0[7]}), .c ({signal_891, signal_546}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_289 ( .s (reset), .b ({data_out_s1[32], data_out_s0[32]}), .a ({data_in_s1[8], data_in_s0[8]}), .c ({signal_894, signal_545}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_290 ( .s (reset), .b ({data_out_s1[36], data_out_s0[36]}), .a ({data_in_s1[9], data_in_s0[9]}), .c ({signal_897, signal_544}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_291 ( .s (reset), .b ({data_out_s1[40], data_out_s0[40]}), .a ({data_in_s1[10], data_in_s0[10]}), .c ({signal_900, signal_543}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_292 ( .s (reset), .b ({data_out_s1[44], data_out_s0[44]}), .a ({data_in_s1[11], data_in_s0[11]}), .c ({signal_903, signal_542}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_293 ( .s (reset), .b ({data_out_s1[48], data_out_s0[48]}), .a ({data_in_s1[12], data_in_s0[12]}), .c ({signal_906, signal_541}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_294 ( .s (reset), .b ({data_out_s1[52], data_out_s0[52]}), .a ({data_in_s1[13], data_in_s0[13]}), .c ({signal_909, signal_540}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_295 ( .s (reset), .b ({data_out_s1[56], data_out_s0[56]}), .a ({data_in_s1[14], data_in_s0[14]}), .c ({signal_912, signal_539}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_296 ( .s (reset), .b ({data_out_s1[60], data_out_s0[60]}), .a ({data_in_s1[15], data_in_s0[15]}), .c ({signal_914, signal_538}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_297 ( .s (reset), .b ({data_out_s1[1], data_out_s0[1]}), .a ({data_in_s1[16], data_in_s0[16]}), .c ({signal_917, signal_537}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_298 ( .s (reset), .b ({data_out_s1[5], data_out_s0[5]}), .a ({data_in_s1[17], data_in_s0[17]}), .c ({signal_920, signal_536}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_299 ( .s (reset), .b ({data_out_s1[9], data_out_s0[9]}), .a ({data_in_s1[18], data_in_s0[18]}), .c ({signal_923, signal_535}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_300 ( .s (reset), .b ({data_out_s1[13], data_out_s0[13]}), .a ({data_in_s1[19], data_in_s0[19]}), .c ({signal_926, signal_534}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_301 ( .s (reset), .b ({data_out_s1[17], data_out_s0[17]}), .a ({data_in_s1[20], data_in_s0[20]}), .c ({signal_929, signal_533}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_302 ( .s (reset), .b ({data_out_s1[21], data_out_s0[21]}), .a ({data_in_s1[21], data_in_s0[21]}), .c ({signal_932, signal_532}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_303 ( .s (reset), .b ({data_out_s1[25], data_out_s0[25]}), .a ({data_in_s1[22], data_in_s0[22]}), .c ({signal_935, signal_531}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_304 ( .s (reset), .b ({data_out_s1[29], data_out_s0[29]}), .a ({data_in_s1[23], data_in_s0[23]}), .c ({signal_938, signal_530}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_305 ( .s (reset), .b ({data_out_s1[33], data_out_s0[33]}), .a ({data_in_s1[24], data_in_s0[24]}), .c ({signal_941, signal_529}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_306 ( .s (reset), .b ({data_out_s1[37], data_out_s0[37]}), .a ({data_in_s1[25], data_in_s0[25]}), .c ({signal_944, signal_528}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_307 ( .s (reset), .b ({data_out_s1[41], data_out_s0[41]}), .a ({data_in_s1[26], data_in_s0[26]}), .c ({signal_947, signal_527}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_308 ( .s (reset), .b ({data_out_s1[45], data_out_s0[45]}), .a ({data_in_s1[27], data_in_s0[27]}), .c ({signal_950, signal_526}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_309 ( .s (reset), .b ({data_out_s1[49], data_out_s0[49]}), .a ({data_in_s1[28], data_in_s0[28]}), .c ({signal_953, signal_525}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_310 ( .s (reset), .b ({data_out_s1[53], data_out_s0[53]}), .a ({data_in_s1[29], data_in_s0[29]}), .c ({signal_956, signal_524}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_311 ( .s (reset), .b ({data_out_s1[57], data_out_s0[57]}), .a ({data_in_s1[30], data_in_s0[30]}), .c ({signal_959, signal_523}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_312 ( .s (reset), .b ({data_out_s1[61], data_out_s0[61]}), .a ({data_in_s1[31], data_in_s0[31]}), .c ({signal_961, signal_522}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_313 ( .s (reset), .b ({data_out_s1[2], data_out_s0[2]}), .a ({data_in_s1[32], data_in_s0[32]}), .c ({signal_964, signal_521}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_314 ( .s (reset), .b ({data_out_s1[6], data_out_s0[6]}), .a ({data_in_s1[33], data_in_s0[33]}), .c ({signal_967, signal_520}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_315 ( .s (reset), .b ({data_out_s1[10], data_out_s0[10]}), .a ({data_in_s1[34], data_in_s0[34]}), .c ({signal_970, signal_519}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_316 ( .s (reset), .b ({data_out_s1[14], data_out_s0[14]}), .a ({data_in_s1[35], data_in_s0[35]}), .c ({signal_973, signal_518}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_317 ( .s (reset), .b ({data_out_s1[18], data_out_s0[18]}), .a ({data_in_s1[36], data_in_s0[36]}), .c ({signal_976, signal_517}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_318 ( .s (reset), .b ({data_out_s1[22], data_out_s0[22]}), .a ({data_in_s1[37], data_in_s0[37]}), .c ({signal_979, signal_516}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_319 ( .s (reset), .b ({data_out_s1[26], data_out_s0[26]}), .a ({data_in_s1[38], data_in_s0[38]}), .c ({signal_982, signal_515}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_320 ( .s (reset), .b ({data_out_s1[30], data_out_s0[30]}), .a ({data_in_s1[39], data_in_s0[39]}), .c ({signal_985, signal_514}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_321 ( .s (reset), .b ({data_out_s1[34], data_out_s0[34]}), .a ({data_in_s1[40], data_in_s0[40]}), .c ({signal_988, signal_513}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_322 ( .s (reset), .b ({data_out_s1[38], data_out_s0[38]}), .a ({data_in_s1[41], data_in_s0[41]}), .c ({signal_991, signal_512}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_323 ( .s (reset), .b ({data_out_s1[42], data_out_s0[42]}), .a ({data_in_s1[42], data_in_s0[42]}), .c ({signal_994, signal_511}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_324 ( .s (reset), .b ({data_out_s1[46], data_out_s0[46]}), .a ({data_in_s1[43], data_in_s0[43]}), .c ({signal_997, signal_510}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_325 ( .s (reset), .b ({data_out_s1[50], data_out_s0[50]}), .a ({data_in_s1[44], data_in_s0[44]}), .c ({signal_1000, signal_509}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_326 ( .s (reset), .b ({data_out_s1[54], data_out_s0[54]}), .a ({data_in_s1[45], data_in_s0[45]}), .c ({signal_1003, signal_508}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_327 ( .s (reset), .b ({data_out_s1[58], data_out_s0[58]}), .a ({data_in_s1[46], data_in_s0[46]}), .c ({signal_1006, signal_507}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_328 ( .s (reset), .b ({data_out_s1[62], data_out_s0[62]}), .a ({data_in_s1[47], data_in_s0[47]}), .c ({signal_1008, signal_506}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_329 ( .s (reset), .b ({data_out_s1[3], data_out_s0[3]}), .a ({data_in_s1[48], data_in_s0[48]}), .c ({signal_1011, signal_505}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_330 ( .s (reset), .b ({data_out_s1[7], data_out_s0[7]}), .a ({data_in_s1[49], data_in_s0[49]}), .c ({signal_1014, signal_504}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_331 ( .s (reset), .b ({data_out_s1[11], data_out_s0[11]}), .a ({data_in_s1[50], data_in_s0[50]}), .c ({signal_1017, signal_503}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_332 ( .s (reset), .b ({data_out_s1[15], data_out_s0[15]}), .a ({data_in_s1[51], data_in_s0[51]}), .c ({signal_1020, signal_502}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_333 ( .s (reset), .b ({data_out_s1[19], data_out_s0[19]}), .a ({data_in_s1[52], data_in_s0[52]}), .c ({signal_1023, signal_501}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_334 ( .s (reset), .b ({data_out_s1[23], data_out_s0[23]}), .a ({data_in_s1[53], data_in_s0[53]}), .c ({signal_1026, signal_500}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_335 ( .s (reset), .b ({data_out_s1[27], data_out_s0[27]}), .a ({data_in_s1[54], data_in_s0[54]}), .c ({signal_1029, signal_499}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_336 ( .s (reset), .b ({data_out_s1[31], data_out_s0[31]}), .a ({data_in_s1[55], data_in_s0[55]}), .c ({signal_1032, signal_498}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_337 ( .s (reset), .b ({data_out_s1[35], data_out_s0[35]}), .a ({data_in_s1[56], data_in_s0[56]}), .c ({signal_1035, signal_497}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_338 ( .s (reset), .b ({data_out_s1[39], data_out_s0[39]}), .a ({data_in_s1[57], data_in_s0[57]}), .c ({signal_1038, signal_496}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_339 ( .s (reset), .b ({data_out_s1[43], data_out_s0[43]}), .a ({data_in_s1[58], data_in_s0[58]}), .c ({signal_1041, signal_495}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_340 ( .s (reset), .b ({data_out_s1[47], data_out_s0[47]}), .a ({data_in_s1[59], data_in_s0[59]}), .c ({signal_1044, signal_494}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_341 ( .s (reset), .b ({data_out_s1[51], data_out_s0[51]}), .a ({data_in_s1[60], data_in_s0[60]}), .c ({signal_1047, signal_493}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_342 ( .s (reset), .b ({data_out_s1[55], data_out_s0[55]}), .a ({data_in_s1[61], data_in_s0[61]}), .c ({signal_1050, signal_492}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_343 ( .s (reset), .b ({data_out_s1[59], data_out_s0[59]}), .a ({data_in_s1[62], data_in_s0[62]}), .c ({signal_1053, signal_491}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_344 ( .s (reset), .b ({data_out_s1[63], data_out_s0[63]}), .a ({data_in_s1[63], data_in_s0[63]}), .c ({signal_1055, signal_490}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_345 ( .a ({1'b0, signal_458}), .b ({signal_1056, signal_676}), .c ({signal_1057, signal_618}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_346 ( .a ({1'b0, signal_459}), .b ({signal_1058, signal_677}), .c ({signal_1059, signal_619}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_347 ( .a ({1'b0, signal_460}), .b ({signal_1060, signal_678}), .c ({signal_1061, signal_620}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_348 ( .a ({1'b0, signal_461}), .b ({signal_1274, signal_679}), .c ({signal_1275, signal_621}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_349 ( .a ({1'b0, signal_462}), .b ({signal_1062, signal_680}), .c ({signal_1063, signal_622}) ) ;
    INV_X1 cell_350 ( .A (signal_356), .ZN (signal_358) ) ;
    INV_X1 cell_351 ( .A (signal_356), .ZN (signal_357) ) ;
    INV_X1 cell_352 ( .A (signal_218), .ZN (signal_356) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_361 ( .s (signal_357), .b ({signal_856, signal_474}), .a ({signal_1066, signal_775}), .c ({signal_1378, signal_779}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_362 ( .s (signal_357), .b ({signal_859, signal_473}), .a ({signal_1069, signal_774}), .c ({signal_1379, signal_778}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_363 ( .s (signal_357), .b ({signal_862, signal_472}), .a ({signal_1072, signal_773}), .c ({signal_1380, signal_777}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_364 ( .s (signal_357), .b ({signal_865, signal_471}), .a ({signal_1075, signal_772}), .c ({signal_1381, signal_776}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_373 ( .s (signal_357), .b ({signal_1287, signal_477}), .a ({signal_1078, signal_771}), .c ({signal_1382, signal_783}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_374 ( .s (signal_357), .b ({signal_1289, signal_476}), .a ({signal_1081, signal_770}), .c ({signal_1383, signal_782}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_375 ( .s (signal_357), .b ({signal_1291, signal_475}), .a ({signal_1084, signal_769}), .c ({signal_1384, signal_781}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_376 ( .s (signal_357), .b ({signal_1064, signal_695}), .a ({signal_1087, signal_768}), .c ({signal_1385, signal_780}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_385 ( .s (signal_358), .b ({signal_1067, signal_694}), .a ({signal_1090, signal_767}), .c ({signal_1386, signal_787}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_386 ( .s (signal_358), .b ({signal_1070, signal_693}), .a ({signal_1093, signal_766}), .c ({signal_1387, signal_786}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_387 ( .s (signal_358), .b ({signal_1073, signal_692}), .a ({signal_1096, signal_765}), .c ({signal_1388, signal_785}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_388 ( .s (signal_358), .b ({signal_1076, signal_691}), .a ({signal_1099, signal_764}), .c ({signal_1389, signal_784}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_397 ( .s (signal_358), .b ({signal_1079, signal_690}), .a ({signal_1102, signal_763}), .c ({signal_1390, signal_791}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_398 ( .s (signal_358), .b ({signal_1082, signal_689}), .a ({signal_1105, signal_762}), .c ({signal_1391, signal_790}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_399 ( .s (signal_358), .b ({signal_1085, signal_688}), .a ({signal_1108, signal_761}), .c ({signal_1392, signal_789}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_400 ( .s (signal_358), .b ({signal_1088, signal_687}), .a ({signal_1277, signal_760}), .c ({signal_1393, signal_788}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_409 ( .s (signal_218), .b ({signal_1091, signal_686}), .a ({signal_1285, signal_759}), .c ({signal_1297, signal_795}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_410 ( .s (signal_218), .b ({signal_1094, signal_685}), .a ({signal_1279, signal_758}), .c ({signal_1298, signal_794}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_411 ( .s (signal_218), .b ({signal_1097, signal_684}), .a ({signal_1281, signal_757}), .c ({signal_1299, signal_793}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_412 ( .s (signal_218), .b ({signal_1100, signal_683}), .a ({signal_1283, signal_756}), .c ({signal_1300, signal_792}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_421 ( .s (signal_218), .b ({signal_1103, signal_682}), .a ({signal_1111, signal_755}), .c ({signal_1301, signal_799}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_422 ( .s (signal_218), .b ({signal_1106, signal_681}), .a ({signal_1114, signal_754}), .c ({signal_1302, signal_798}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_423 ( .s (signal_218), .b ({signal_1062, signal_680}), .a ({signal_1117, signal_753}), .c ({signal_1303, signal_797}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_424 ( .s (signal_218), .b ({signal_1274, signal_679}), .a ({signal_1120, signal_752}), .c ({signal_1304, signal_796}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_433 ( .s (signal_357), .b ({signal_1060, signal_678}), .a ({signal_1123, signal_751}), .c ({signal_1394, signal_803}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_434 ( .s (signal_357), .b ({signal_1058, signal_677}), .a ({signal_1126, signal_750}), .c ({signal_1395, signal_802}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_435 ( .s (signal_357), .b ({signal_1056, signal_676}), .a ({signal_1129, signal_749}), .c ({signal_1396, signal_801}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_436 ( .s (signal_357), .b ({signal_1109, signal_675}), .a ({signal_1132, signal_748}), .c ({signal_1397, signal_800}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_445 ( .s (signal_357), .b ({signal_1112, signal_674}), .a ({signal_1135, signal_747}), .c ({signal_1398, signal_807}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_446 ( .s (signal_357), .b ({signal_1115, signal_673}), .a ({signal_1138, signal_746}), .c ({signal_1399, signal_806}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_447 ( .s (signal_357), .b ({signal_1118, signal_672}), .a ({signal_1141, signal_745}), .c ({signal_1400, signal_805}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_448 ( .s (signal_357), .b ({signal_1121, signal_671}), .a ({signal_1144, signal_744}), .c ({signal_1401, signal_804}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_457 ( .s (signal_357), .b ({signal_1124, signal_670}), .a ({signal_1147, signal_743}), .c ({signal_1402, signal_811}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_458 ( .s (signal_357), .b ({signal_1127, signal_669}), .a ({signal_1150, signal_742}), .c ({signal_1403, signal_810}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_459 ( .s (signal_357), .b ({signal_1130, signal_668}), .a ({signal_1153, signal_741}), .c ({signal_1404, signal_809}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_460 ( .s (signal_357), .b ({signal_1133, signal_667}), .a ({signal_1156, signal_740}), .c ({signal_1405, signal_808}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_469 ( .s (signal_357), .b ({signal_1136, signal_666}), .a ({signal_1159, signal_739}), .c ({signal_1406, signal_815}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_470 ( .s (signal_357), .b ({signal_1139, signal_665}), .a ({signal_1162, signal_738}), .c ({signal_1407, signal_814}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_471 ( .s (signal_357), .b ({signal_1142, signal_664}), .a ({signal_1165, signal_737}), .c ({signal_1408, signal_813}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_472 ( .s (signal_357), .b ({signal_1145, signal_663}), .a ({signal_1168, signal_736}), .c ({signal_1409, signal_812}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_481 ( .s (signal_357), .b ({signal_1148, signal_662}), .a ({signal_1171, signal_735}), .c ({signal_1410, signal_819}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_482 ( .s (signal_357), .b ({signal_1151, signal_661}), .a ({signal_1174, signal_734}), .c ({signal_1411, signal_818}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_483 ( .s (signal_357), .b ({signal_1154, signal_660}), .a ({signal_1177, signal_733}), .c ({signal_1412, signal_817}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_484 ( .s (signal_357), .b ({signal_1157, signal_659}), .a ({signal_1180, signal_732}), .c ({signal_1413, signal_816}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_493 ( .s (signal_357), .b ({signal_1160, signal_658}), .a ({signal_1183, signal_731}), .c ({signal_1414, signal_823}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_494 ( .s (signal_357), .b ({signal_1163, signal_657}), .a ({signal_1186, signal_730}), .c ({signal_1415, signal_822}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_495 ( .s (signal_357), .b ({signal_1166, signal_656}), .a ({signal_1189, signal_729}), .c ({signal_1416, signal_821}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_496 ( .s (signal_357), .b ({signal_1169, signal_655}), .a ({signal_1192, signal_728}), .c ({signal_1417, signal_820}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_505 ( .s (signal_357), .b ({signal_1172, signal_654}), .a ({signal_1195, signal_727}), .c ({signal_1418, signal_827}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_506 ( .s (signal_357), .b ({signal_1175, signal_653}), .a ({signal_1198, signal_726}), .c ({signal_1419, signal_826}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_507 ( .s (signal_357), .b ({signal_1178, signal_652}), .a ({signal_1201, signal_725}), .c ({signal_1420, signal_825}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_508 ( .s (signal_357), .b ({signal_1181, signal_651}), .a ({signal_1204, signal_724}), .c ({signal_1421, signal_824}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_517 ( .s (signal_358), .b ({signal_1184, signal_650}), .a ({signal_1207, signal_723}), .c ({signal_1422, signal_831}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_518 ( .s (signal_358), .b ({signal_1187, signal_649}), .a ({signal_1210, signal_722}), .c ({signal_1423, signal_830}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_519 ( .s (signal_358), .b ({signal_1190, signal_648}), .a ({signal_1213, signal_721}), .c ({signal_1424, signal_829}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_520 ( .s (signal_358), .b ({signal_1193, signal_647}), .a ({signal_1216, signal_720}), .c ({signal_1425, signal_828}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_529 ( .s (signal_358), .b ({signal_1196, signal_646}), .a ({signal_1219, signal_719}), .c ({signal_1426, signal_835}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_530 ( .s (signal_358), .b ({signal_1199, signal_645}), .a ({signal_1222, signal_718}), .c ({signal_1427, signal_834}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_531 ( .s (signal_358), .b ({signal_1202, signal_644}), .a ({signal_1225, signal_717}), .c ({signal_1428, signal_833}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_532 ( .s (signal_358), .b ({signal_1205, signal_643}), .a ({signal_1228, signal_716}), .c ({signal_1429, signal_832}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_541 ( .s (signal_358), .b ({signal_1208, signal_642}), .a ({signal_1231, signal_715}), .c ({signal_1430, signal_839}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_542 ( .s (signal_358), .b ({signal_1211, signal_641}), .a ({signal_1234, signal_714}), .c ({signal_1431, signal_838}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_543 ( .s (signal_358), .b ({signal_1214, signal_640}), .a ({signal_1237, signal_713}), .c ({signal_1432, signal_837}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_544 ( .s (signal_358), .b ({signal_1217, signal_639}), .a ({signal_1240, signal_712}), .c ({signal_1433, signal_836}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_553 ( .s (signal_358), .b ({signal_1220, signal_638}), .a ({signal_1243, signal_711}), .c ({signal_1434, signal_843}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_554 ( .s (signal_358), .b ({signal_1223, signal_637}), .a ({signal_1246, signal_710}), .c ({signal_1435, signal_842}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_555 ( .s (signal_358), .b ({signal_1226, signal_636}), .a ({signal_1249, signal_709}), .c ({signal_1436, signal_841}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_556 ( .s (signal_358), .b ({signal_1229, signal_635}), .a ({signal_1252, signal_708}), .c ({signal_1437, signal_840}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_565 ( .s (signal_358), .b ({signal_1232, signal_634}), .a ({signal_1255, signal_707}), .c ({signal_1438, signal_847}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_566 ( .s (signal_358), .b ({signal_1235, signal_633}), .a ({signal_1258, signal_706}), .c ({signal_1439, signal_846}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_567 ( .s (signal_358), .b ({signal_1238, signal_632}), .a ({signal_1261, signal_705}), .c ({signal_1440, signal_845}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_568 ( .s (signal_358), .b ({signal_1241, signal_631}), .a ({signal_1264, signal_704}), .c ({signal_1441, signal_844}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_577 ( .s (signal_358), .b ({signal_1244, signal_630}), .a ({signal_1267, signal_703}), .c ({signal_1442, signal_851}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_578 ( .s (signal_358), .b ({signal_1247, signal_629}), .a ({signal_1269, signal_702}), .c ({signal_1443, signal_850}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_579 ( .s (signal_358), .b ({signal_1250, signal_628}), .a ({signal_1271, signal_701}), .c ({signal_1444, signal_849}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_580 ( .s (signal_358), .b ({signal_1253, signal_627}), .a ({signal_1273, signal_700}), .c ({signal_1445, signal_848}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_593 ( .s (reset), .b ({signal_1064, signal_695}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1066, signal_775}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_594 ( .s (reset), .b ({signal_1067, signal_694}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1069, signal_774}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_595 ( .s (reset), .b ({signal_1070, signal_693}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1072, signal_773}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_596 ( .s (reset), .b ({signal_1073, signal_692}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1075, signal_772}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_597 ( .s (reset), .b ({signal_1076, signal_691}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1078, signal_771}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_598 ( .s (reset), .b ({signal_1079, signal_690}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1081, signal_770}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_599 ( .s (reset), .b ({signal_1082, signal_689}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1084, signal_769}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_600 ( .s (reset), .b ({signal_1085, signal_688}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1087, signal_768}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_601 ( .s (reset), .b ({signal_1088, signal_687}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1090, signal_767}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_602 ( .s (reset), .b ({signal_1091, signal_686}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1093, signal_766}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_603 ( .s (reset), .b ({signal_1094, signal_685}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1096, signal_765}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_604 ( .s (reset), .b ({signal_1097, signal_684}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1099, signal_764}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_605 ( .s (reset), .b ({signal_1100, signal_683}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1102, signal_763}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_606 ( .s (reset), .b ({signal_1103, signal_682}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1105, signal_762}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_607 ( .s (reset), .b ({signal_1106, signal_681}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1108, signal_761}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_608 ( .s (reset), .b ({signal_1063, signal_622}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1277, signal_760}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_609 ( .s (reset), .b ({signal_1275, signal_621}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1285, signal_759}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_610 ( .s (reset), .b ({signal_1061, signal_620}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1279, signal_758}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_611 ( .s (reset), .b ({signal_1059, signal_619}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1281, signal_757}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_612 ( .s (reset), .b ({signal_1057, signal_618}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1283, signal_756}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_613 ( .s (reset), .b ({signal_1109, signal_675}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1111, signal_755}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_614 ( .s (reset), .b ({signal_1112, signal_674}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1114, signal_754}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_615 ( .s (reset), .b ({signal_1115, signal_673}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1117, signal_753}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_616 ( .s (reset), .b ({signal_1118, signal_672}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1120, signal_752}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_617 ( .s (reset), .b ({signal_1121, signal_671}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1123, signal_751}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_618 ( .s (reset), .b ({signal_1124, signal_670}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1126, signal_750}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_619 ( .s (reset), .b ({signal_1127, signal_669}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1129, signal_749}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_620 ( .s (reset), .b ({signal_1130, signal_668}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1132, signal_748}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_621 ( .s (reset), .b ({signal_1133, signal_667}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1135, signal_747}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_622 ( .s (reset), .b ({signal_1136, signal_666}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1138, signal_746}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_623 ( .s (reset), .b ({signal_1139, signal_665}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1141, signal_745}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_624 ( .s (reset), .b ({signal_1142, signal_664}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1144, signal_744}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_625 ( .s (reset), .b ({signal_1145, signal_663}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1147, signal_743}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_626 ( .s (reset), .b ({signal_1148, signal_662}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1150, signal_742}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_627 ( .s (reset), .b ({signal_1151, signal_661}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1153, signal_741}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_628 ( .s (reset), .b ({signal_1154, signal_660}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1156, signal_740}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_629 ( .s (reset), .b ({signal_1157, signal_659}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1159, signal_739}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_630 ( .s (reset), .b ({signal_1160, signal_658}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1162, signal_738}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_631 ( .s (reset), .b ({signal_1163, signal_657}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1165, signal_737}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_632 ( .s (reset), .b ({signal_1166, signal_656}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1168, signal_736}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_633 ( .s (reset), .b ({signal_1169, signal_655}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1171, signal_735}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_634 ( .s (reset), .b ({signal_1172, signal_654}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1174, signal_734}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_635 ( .s (reset), .b ({signal_1175, signal_653}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1177, signal_733}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_636 ( .s (reset), .b ({signal_1178, signal_652}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1180, signal_732}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_637 ( .s (reset), .b ({signal_1181, signal_651}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1183, signal_731}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_638 ( .s (reset), .b ({signal_1184, signal_650}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1186, signal_730}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_639 ( .s (reset), .b ({signal_1187, signal_649}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1189, signal_729}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_640 ( .s (reset), .b ({signal_1190, signal_648}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1192, signal_728}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_641 ( .s (reset), .b ({signal_1193, signal_647}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1195, signal_727}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_642 ( .s (reset), .b ({signal_1196, signal_646}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1198, signal_726}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_643 ( .s (reset), .b ({signal_1199, signal_645}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1201, signal_725}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_644 ( .s (reset), .b ({signal_1202, signal_644}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1204, signal_724}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_645 ( .s (reset), .b ({signal_1205, signal_643}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1207, signal_723}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_646 ( .s (reset), .b ({signal_1208, signal_642}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1210, signal_722}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_647 ( .s (reset), .b ({signal_1211, signal_641}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1213, signal_721}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_648 ( .s (reset), .b ({signal_1214, signal_640}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1216, signal_720}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_649 ( .s (reset), .b ({signal_1217, signal_639}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1219, signal_719}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_650 ( .s (reset), .b ({signal_1220, signal_638}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1222, signal_718}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_651 ( .s (reset), .b ({signal_1223, signal_637}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1225, signal_717}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_652 ( .s (reset), .b ({signal_1226, signal_636}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1228, signal_716}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_653 ( .s (reset), .b ({signal_1229, signal_635}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1231, signal_715}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_654 ( .s (reset), .b ({signal_1232, signal_634}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1234, signal_714}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_655 ( .s (reset), .b ({signal_1235, signal_633}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1237, signal_713}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_656 ( .s (reset), .b ({signal_1238, signal_632}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1240, signal_712}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_657 ( .s (reset), .b ({signal_1241, signal_631}), .a ({key_s1[64], key_s0[64]}), .c ({signal_1243, signal_711}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_658 ( .s (reset), .b ({signal_1244, signal_630}), .a ({key_s1[65], key_s0[65]}), .c ({signal_1246, signal_710}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_659 ( .s (reset), .b ({signal_1247, signal_629}), .a ({key_s1[66], key_s0[66]}), .c ({signal_1249, signal_709}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_660 ( .s (reset), .b ({signal_1250, signal_628}), .a ({key_s1[67], key_s0[67]}), .c ({signal_1252, signal_708}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_661 ( .s (reset), .b ({signal_1253, signal_627}), .a ({key_s1[68], key_s0[68]}), .c ({signal_1255, signal_707}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_662 ( .s (reset), .b ({signal_1256, signal_626}), .a ({key_s1[69], key_s0[69]}), .c ({signal_1258, signal_706}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_663 ( .s (reset), .b ({signal_1259, signal_625}), .a ({key_s1[70], key_s0[70]}), .c ({signal_1261, signal_705}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_664 ( .s (reset), .b ({signal_1262, signal_624}), .a ({key_s1[71], key_s0[71]}), .c ({signal_1264, signal_704}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_665 ( .s (reset), .b ({signal_1265, signal_623}), .a ({key_s1[72], key_s0[72]}), .c ({signal_1267, signal_703}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_666 ( .s (reset), .b ({signal_856, signal_474}), .a ({key_s1[73], key_s0[73]}), .c ({signal_1269, signal_702}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_667 ( .s (reset), .b ({signal_859, signal_473}), .a ({key_s1[74], key_s0[74]}), .c ({signal_1271, signal_701}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_668 ( .s (reset), .b ({signal_862, signal_472}), .a ({key_s1[75], key_s0[75]}), .c ({signal_1273, signal_700}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_696 ( .s (signal_217), .b ({signal_858, signal_485}), .a ({signal_865, signal_471}), .c ({signal_1286, signal_481}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_697 ( .s (signal_217), .b ({signal_861, signal_484}), .a ({signal_1287, signal_477}), .c ({signal_1288, signal_480}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_698 ( .s (signal_217), .b ({signal_864, signal_483}), .a ({signal_1289, signal_476}), .c ({signal_1290, signal_479}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_699 ( .s (signal_217), .b ({signal_867, signal_482}), .a ({signal_1291, signal_475}), .c ({signal_1292, signal_478}) ) ;

    /* cells in depth 1 */
    buf_clk cell_705 ( .C (clk), .D (signal_218), .Q (signal_1458) ) ;
    buf_clk cell_707 ( .C (clk), .D (signal_553), .Q (signal_1460) ) ;
    buf_clk cell_709 ( .C (clk), .D (signal_870), .Q (signal_1462) ) ;
    buf_clk cell_711 ( .C (clk), .D (signal_552), .Q (signal_1464) ) ;
    buf_clk cell_713 ( .C (clk), .D (signal_873), .Q (signal_1466) ) ;
    buf_clk cell_715 ( .C (clk), .D (signal_551), .Q (signal_1468) ) ;
    buf_clk cell_717 ( .C (clk), .D (signal_876), .Q (signal_1470) ) ;
    buf_clk cell_719 ( .C (clk), .D (signal_550), .Q (signal_1472) ) ;
    buf_clk cell_721 ( .C (clk), .D (signal_879), .Q (signal_1474) ) ;
    buf_clk cell_723 ( .C (clk), .D (signal_358), .Q (signal_1476) ) ;
    buf_clk cell_725 ( .C (clk), .D (signal_626), .Q (signal_1478) ) ;
    buf_clk cell_727 ( .C (clk), .D (signal_1256), .Q (signal_1480) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_625), .Q (signal_1482) ) ;
    buf_clk cell_731 ( .C (clk), .D (signal_1259), .Q (signal_1484) ) ;
    buf_clk cell_733 ( .C (clk), .D (signal_624), .Q (signal_1486) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_1262), .Q (signal_1488) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_623), .Q (signal_1490) ) ;
    buf_clk cell_739 ( .C (clk), .D (signal_1265), .Q (signal_1492) ) ;
    buf_clk cell_741 ( .C (clk), .D (reset), .Q (signal_1494) ) ;
    buf_clk cell_743 ( .C (clk), .D (key_s0[76]), .Q (signal_1496) ) ;
    buf_clk cell_745 ( .C (clk), .D (key_s1[76]), .Q (signal_1498) ) ;
    buf_clk cell_747 ( .C (clk), .D (key_s0[77]), .Q (signal_1500) ) ;
    buf_clk cell_749 ( .C (clk), .D (key_s1[77]), .Q (signal_1502) ) ;
    buf_clk cell_751 ( .C (clk), .D (key_s0[78]), .Q (signal_1504) ) ;
    buf_clk cell_753 ( .C (clk), .D (key_s1[78]), .Q (signal_1506) ) ;
    buf_clk cell_755 ( .C (clk), .D (key_s0[79]), .Q (signal_1508) ) ;
    buf_clk cell_757 ( .C (clk), .D (key_s1[79]), .Q (signal_1510) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_481), .Q (signal_1512) ) ;
    buf_clk cell_761 ( .C (clk), .D (signal_1286), .Q (signal_1514) ) ;
    buf_clk cell_763 ( .C (clk), .D (signal_219), .Q (signal_1516) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_485), .Q (signal_1518) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_858), .Q (signal_1520) ) ;
    buf_clk cell_769 ( .C (clk), .D (signal_484), .Q (signal_1522) ) ;
    buf_clk cell_771 ( .C (clk), .D (signal_861), .Q (signal_1524) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_483), .Q (signal_1526) ) ;
    buf_clk cell_775 ( .C (clk), .D (signal_864), .Q (signal_1528) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_482), .Q (signal_1530) ) ;
    buf_clk cell_779 ( .C (clk), .D (signal_867), .Q (signal_1532) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_271), .Q (signal_1534) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_270), .Q (signal_1536) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_269), .Q (signal_1538) ) ;
    buf_clk cell_787 ( .C (clk), .D (signal_268), .Q (signal_1540) ) ;
    buf_clk cell_789 ( .C (clk), .D (signal_266), .Q (signal_1542) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_285), .Q (signal_1544) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_284), .Q (signal_1546) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_283), .Q (signal_1548) ) ;
    buf_clk cell_797 ( .C (clk), .D (signal_282), .Q (signal_1550) ) ;
    buf_clk cell_799 ( .C (clk), .D (signal_236), .Q (signal_1552) ) ;
    buf_clk cell_801 ( .C (clk), .D (signal_233), .Q (signal_1554) ) ;
    buf_clk cell_803 ( .C (clk), .D (signal_558), .Q (signal_1556) ) ;
    buf_clk cell_805 ( .C (clk), .D (signal_1296), .Q (signal_1558) ) ;
    buf_clk cell_807 ( .C (clk), .D (signal_559), .Q (signal_1560) ) ;
    buf_clk cell_809 ( .C (clk), .D (signal_1295), .Q (signal_1562) ) ;
    buf_clk cell_811 ( .C (clk), .D (signal_560), .Q (signal_1564) ) ;
    buf_clk cell_813 ( .C (clk), .D (signal_1294), .Q (signal_1566) ) ;
    buf_clk cell_815 ( .C (clk), .D (signal_561), .Q (signal_1568) ) ;
    buf_clk cell_817 ( .C (clk), .D (signal_1293), .Q (signal_1570) ) ;
    buf_clk cell_819 ( .C (clk), .D (signal_562), .Q (signal_1572) ) ;
    buf_clk cell_821 ( .C (clk), .D (signal_1325), .Q (signal_1574) ) ;
    buf_clk cell_823 ( .C (clk), .D (signal_563), .Q (signal_1576) ) ;
    buf_clk cell_825 ( .C (clk), .D (signal_1324), .Q (signal_1578) ) ;
    buf_clk cell_827 ( .C (clk), .D (signal_564), .Q (signal_1580) ) ;
    buf_clk cell_829 ( .C (clk), .D (signal_1323), .Q (signal_1582) ) ;
    buf_clk cell_831 ( .C (clk), .D (signal_565), .Q (signal_1584) ) ;
    buf_clk cell_833 ( .C (clk), .D (signal_1322), .Q (signal_1586) ) ;
    buf_clk cell_835 ( .C (clk), .D (signal_566), .Q (signal_1588) ) ;
    buf_clk cell_837 ( .C (clk), .D (signal_1329), .Q (signal_1590) ) ;
    buf_clk cell_839 ( .C (clk), .D (signal_567), .Q (signal_1592) ) ;
    buf_clk cell_841 ( .C (clk), .D (signal_1328), .Q (signal_1594) ) ;
    buf_clk cell_843 ( .C (clk), .D (signal_568), .Q (signal_1596) ) ;
    buf_clk cell_845 ( .C (clk), .D (signal_1327), .Q (signal_1598) ) ;
    buf_clk cell_847 ( .C (clk), .D (signal_569), .Q (signal_1600) ) ;
    buf_clk cell_849 ( .C (clk), .D (signal_1326), .Q (signal_1602) ) ;
    buf_clk cell_851 ( .C (clk), .D (signal_570), .Q (signal_1604) ) ;
    buf_clk cell_853 ( .C (clk), .D (signal_1333), .Q (signal_1606) ) ;
    buf_clk cell_855 ( .C (clk), .D (signal_571), .Q (signal_1608) ) ;
    buf_clk cell_857 ( .C (clk), .D (signal_1332), .Q (signal_1610) ) ;
    buf_clk cell_859 ( .C (clk), .D (signal_572), .Q (signal_1612) ) ;
    buf_clk cell_861 ( .C (clk), .D (signal_1331), .Q (signal_1614) ) ;
    buf_clk cell_863 ( .C (clk), .D (signal_573), .Q (signal_1616) ) ;
    buf_clk cell_865 ( .C (clk), .D (signal_1330), .Q (signal_1618) ) ;
    buf_clk cell_867 ( .C (clk), .D (signal_574), .Q (signal_1620) ) ;
    buf_clk cell_869 ( .C (clk), .D (signal_1337), .Q (signal_1622) ) ;
    buf_clk cell_871 ( .C (clk), .D (signal_575), .Q (signal_1624) ) ;
    buf_clk cell_873 ( .C (clk), .D (signal_1336), .Q (signal_1626) ) ;
    buf_clk cell_875 ( .C (clk), .D (signal_576), .Q (signal_1628) ) ;
    buf_clk cell_877 ( .C (clk), .D (signal_1335), .Q (signal_1630) ) ;
    buf_clk cell_879 ( .C (clk), .D (signal_577), .Q (signal_1632) ) ;
    buf_clk cell_881 ( .C (clk), .D (signal_1334), .Q (signal_1634) ) ;
    buf_clk cell_883 ( .C (clk), .D (signal_578), .Q (signal_1636) ) ;
    buf_clk cell_885 ( .C (clk), .D (signal_1341), .Q (signal_1638) ) ;
    buf_clk cell_887 ( .C (clk), .D (signal_579), .Q (signal_1640) ) ;
    buf_clk cell_889 ( .C (clk), .D (signal_1340), .Q (signal_1642) ) ;
    buf_clk cell_891 ( .C (clk), .D (signal_580), .Q (signal_1644) ) ;
    buf_clk cell_893 ( .C (clk), .D (signal_1339), .Q (signal_1646) ) ;
    buf_clk cell_895 ( .C (clk), .D (signal_581), .Q (signal_1648) ) ;
    buf_clk cell_897 ( .C (clk), .D (signal_1338), .Q (signal_1650) ) ;
    buf_clk cell_899 ( .C (clk), .D (signal_582), .Q (signal_1652) ) ;
    buf_clk cell_901 ( .C (clk), .D (signal_1345), .Q (signal_1654) ) ;
    buf_clk cell_903 ( .C (clk), .D (signal_583), .Q (signal_1656) ) ;
    buf_clk cell_905 ( .C (clk), .D (signal_1344), .Q (signal_1658) ) ;
    buf_clk cell_907 ( .C (clk), .D (signal_584), .Q (signal_1660) ) ;
    buf_clk cell_909 ( .C (clk), .D (signal_1343), .Q (signal_1662) ) ;
    buf_clk cell_911 ( .C (clk), .D (signal_585), .Q (signal_1664) ) ;
    buf_clk cell_913 ( .C (clk), .D (signal_1342), .Q (signal_1666) ) ;
    buf_clk cell_915 ( .C (clk), .D (signal_586), .Q (signal_1668) ) ;
    buf_clk cell_917 ( .C (clk), .D (signal_1349), .Q (signal_1670) ) ;
    buf_clk cell_919 ( .C (clk), .D (signal_587), .Q (signal_1672) ) ;
    buf_clk cell_921 ( .C (clk), .D (signal_1348), .Q (signal_1674) ) ;
    buf_clk cell_923 ( .C (clk), .D (signal_588), .Q (signal_1676) ) ;
    buf_clk cell_925 ( .C (clk), .D (signal_1347), .Q (signal_1678) ) ;
    buf_clk cell_927 ( .C (clk), .D (signal_589), .Q (signal_1680) ) ;
    buf_clk cell_929 ( .C (clk), .D (signal_1346), .Q (signal_1682) ) ;
    buf_clk cell_931 ( .C (clk), .D (signal_590), .Q (signal_1684) ) ;
    buf_clk cell_933 ( .C (clk), .D (signal_1353), .Q (signal_1686) ) ;
    buf_clk cell_935 ( .C (clk), .D (signal_591), .Q (signal_1688) ) ;
    buf_clk cell_937 ( .C (clk), .D (signal_1352), .Q (signal_1690) ) ;
    buf_clk cell_939 ( .C (clk), .D (signal_592), .Q (signal_1692) ) ;
    buf_clk cell_941 ( .C (clk), .D (signal_1351), .Q (signal_1694) ) ;
    buf_clk cell_943 ( .C (clk), .D (signal_593), .Q (signal_1696) ) ;
    buf_clk cell_945 ( .C (clk), .D (signal_1350), .Q (signal_1698) ) ;
    buf_clk cell_947 ( .C (clk), .D (signal_594), .Q (signal_1700) ) ;
    buf_clk cell_949 ( .C (clk), .D (signal_1357), .Q (signal_1702) ) ;
    buf_clk cell_951 ( .C (clk), .D (signal_595), .Q (signal_1704) ) ;
    buf_clk cell_953 ( .C (clk), .D (signal_1356), .Q (signal_1706) ) ;
    buf_clk cell_955 ( .C (clk), .D (signal_596), .Q (signal_1708) ) ;
    buf_clk cell_957 ( .C (clk), .D (signal_1355), .Q (signal_1710) ) ;
    buf_clk cell_959 ( .C (clk), .D (signal_597), .Q (signal_1712) ) ;
    buf_clk cell_961 ( .C (clk), .D (signal_1354), .Q (signal_1714) ) ;
    buf_clk cell_963 ( .C (clk), .D (signal_598), .Q (signal_1716) ) ;
    buf_clk cell_965 ( .C (clk), .D (signal_1361), .Q (signal_1718) ) ;
    buf_clk cell_967 ( .C (clk), .D (signal_599), .Q (signal_1720) ) ;
    buf_clk cell_969 ( .C (clk), .D (signal_1360), .Q (signal_1722) ) ;
    buf_clk cell_971 ( .C (clk), .D (signal_600), .Q (signal_1724) ) ;
    buf_clk cell_973 ( .C (clk), .D (signal_1359), .Q (signal_1726) ) ;
    buf_clk cell_975 ( .C (clk), .D (signal_601), .Q (signal_1728) ) ;
    buf_clk cell_977 ( .C (clk), .D (signal_1358), .Q (signal_1730) ) ;
    buf_clk cell_979 ( .C (clk), .D (signal_602), .Q (signal_1732) ) ;
    buf_clk cell_981 ( .C (clk), .D (signal_1365), .Q (signal_1734) ) ;
    buf_clk cell_983 ( .C (clk), .D (signal_603), .Q (signal_1736) ) ;
    buf_clk cell_985 ( .C (clk), .D (signal_1364), .Q (signal_1738) ) ;
    buf_clk cell_987 ( .C (clk), .D (signal_604), .Q (signal_1740) ) ;
    buf_clk cell_989 ( .C (clk), .D (signal_1363), .Q (signal_1742) ) ;
    buf_clk cell_991 ( .C (clk), .D (signal_605), .Q (signal_1744) ) ;
    buf_clk cell_993 ( .C (clk), .D (signal_1362), .Q (signal_1746) ) ;
    buf_clk cell_995 ( .C (clk), .D (signal_606), .Q (signal_1748) ) ;
    buf_clk cell_997 ( .C (clk), .D (signal_1369), .Q (signal_1750) ) ;
    buf_clk cell_999 ( .C (clk), .D (signal_607), .Q (signal_1752) ) ;
    buf_clk cell_1001 ( .C (clk), .D (signal_1368), .Q (signal_1754) ) ;
    buf_clk cell_1003 ( .C (clk), .D (signal_608), .Q (signal_1756) ) ;
    buf_clk cell_1005 ( .C (clk), .D (signal_1367), .Q (signal_1758) ) ;
    buf_clk cell_1007 ( .C (clk), .D (signal_609), .Q (signal_1760) ) ;
    buf_clk cell_1009 ( .C (clk), .D (signal_1366), .Q (signal_1762) ) ;
    buf_clk cell_1011 ( .C (clk), .D (signal_610), .Q (signal_1764) ) ;
    buf_clk cell_1013 ( .C (clk), .D (signal_1373), .Q (signal_1766) ) ;
    buf_clk cell_1015 ( .C (clk), .D (signal_611), .Q (signal_1768) ) ;
    buf_clk cell_1017 ( .C (clk), .D (signal_1372), .Q (signal_1770) ) ;
    buf_clk cell_1019 ( .C (clk), .D (signal_612), .Q (signal_1772) ) ;
    buf_clk cell_1021 ( .C (clk), .D (signal_1371), .Q (signal_1774) ) ;
    buf_clk cell_1023 ( .C (clk), .D (signal_613), .Q (signal_1776) ) ;
    buf_clk cell_1025 ( .C (clk), .D (signal_1370), .Q (signal_1778) ) ;
    buf_clk cell_1027 ( .C (clk), .D (signal_614), .Q (signal_1780) ) ;
    buf_clk cell_1029 ( .C (clk), .D (signal_1377), .Q (signal_1782) ) ;
    buf_clk cell_1031 ( .C (clk), .D (signal_615), .Q (signal_1784) ) ;
    buf_clk cell_1033 ( .C (clk), .D (signal_1376), .Q (signal_1786) ) ;
    buf_clk cell_1035 ( .C (clk), .D (signal_616), .Q (signal_1788) ) ;
    buf_clk cell_1037 ( .C (clk), .D (signal_1375), .Q (signal_1790) ) ;
    buf_clk cell_1039 ( .C (clk), .D (signal_617), .Q (signal_1792) ) ;
    buf_clk cell_1041 ( .C (clk), .D (signal_1374), .Q (signal_1794) ) ;
    buf_clk cell_1043 ( .C (clk), .D (signal_776), .Q (signal_1796) ) ;
    buf_clk cell_1045 ( .C (clk), .D (signal_1381), .Q (signal_1798) ) ;
    buf_clk cell_1047 ( .C (clk), .D (signal_777), .Q (signal_1800) ) ;
    buf_clk cell_1049 ( .C (clk), .D (signal_1380), .Q (signal_1802) ) ;
    buf_clk cell_1051 ( .C (clk), .D (signal_778), .Q (signal_1804) ) ;
    buf_clk cell_1053 ( .C (clk), .D (signal_1379), .Q (signal_1806) ) ;
    buf_clk cell_1055 ( .C (clk), .D (signal_779), .Q (signal_1808) ) ;
    buf_clk cell_1057 ( .C (clk), .D (signal_1378), .Q (signal_1810) ) ;
    buf_clk cell_1059 ( .C (clk), .D (signal_780), .Q (signal_1812) ) ;
    buf_clk cell_1061 ( .C (clk), .D (signal_1385), .Q (signal_1814) ) ;
    buf_clk cell_1063 ( .C (clk), .D (signal_781), .Q (signal_1816) ) ;
    buf_clk cell_1065 ( .C (clk), .D (signal_1384), .Q (signal_1818) ) ;
    buf_clk cell_1067 ( .C (clk), .D (signal_782), .Q (signal_1820) ) ;
    buf_clk cell_1069 ( .C (clk), .D (signal_1383), .Q (signal_1822) ) ;
    buf_clk cell_1071 ( .C (clk), .D (signal_783), .Q (signal_1824) ) ;
    buf_clk cell_1073 ( .C (clk), .D (signal_1382), .Q (signal_1826) ) ;
    buf_clk cell_1075 ( .C (clk), .D (signal_784), .Q (signal_1828) ) ;
    buf_clk cell_1077 ( .C (clk), .D (signal_1389), .Q (signal_1830) ) ;
    buf_clk cell_1079 ( .C (clk), .D (signal_785), .Q (signal_1832) ) ;
    buf_clk cell_1081 ( .C (clk), .D (signal_1388), .Q (signal_1834) ) ;
    buf_clk cell_1083 ( .C (clk), .D (signal_786), .Q (signal_1836) ) ;
    buf_clk cell_1085 ( .C (clk), .D (signal_1387), .Q (signal_1838) ) ;
    buf_clk cell_1087 ( .C (clk), .D (signal_787), .Q (signal_1840) ) ;
    buf_clk cell_1089 ( .C (clk), .D (signal_1386), .Q (signal_1842) ) ;
    buf_clk cell_1091 ( .C (clk), .D (signal_788), .Q (signal_1844) ) ;
    buf_clk cell_1093 ( .C (clk), .D (signal_1393), .Q (signal_1846) ) ;
    buf_clk cell_1095 ( .C (clk), .D (signal_789), .Q (signal_1848) ) ;
    buf_clk cell_1097 ( .C (clk), .D (signal_1392), .Q (signal_1850) ) ;
    buf_clk cell_1099 ( .C (clk), .D (signal_790), .Q (signal_1852) ) ;
    buf_clk cell_1101 ( .C (clk), .D (signal_1391), .Q (signal_1854) ) ;
    buf_clk cell_1103 ( .C (clk), .D (signal_791), .Q (signal_1856) ) ;
    buf_clk cell_1105 ( .C (clk), .D (signal_1390), .Q (signal_1858) ) ;
    buf_clk cell_1107 ( .C (clk), .D (signal_792), .Q (signal_1860) ) ;
    buf_clk cell_1109 ( .C (clk), .D (signal_1300), .Q (signal_1862) ) ;
    buf_clk cell_1111 ( .C (clk), .D (signal_793), .Q (signal_1864) ) ;
    buf_clk cell_1113 ( .C (clk), .D (signal_1299), .Q (signal_1866) ) ;
    buf_clk cell_1115 ( .C (clk), .D (signal_794), .Q (signal_1868) ) ;
    buf_clk cell_1117 ( .C (clk), .D (signal_1298), .Q (signal_1870) ) ;
    buf_clk cell_1119 ( .C (clk), .D (signal_795), .Q (signal_1872) ) ;
    buf_clk cell_1121 ( .C (clk), .D (signal_1297), .Q (signal_1874) ) ;
    buf_clk cell_1123 ( .C (clk), .D (signal_796), .Q (signal_1876) ) ;
    buf_clk cell_1125 ( .C (clk), .D (signal_1304), .Q (signal_1878) ) ;
    buf_clk cell_1127 ( .C (clk), .D (signal_797), .Q (signal_1880) ) ;
    buf_clk cell_1129 ( .C (clk), .D (signal_1303), .Q (signal_1882) ) ;
    buf_clk cell_1131 ( .C (clk), .D (signal_798), .Q (signal_1884) ) ;
    buf_clk cell_1133 ( .C (clk), .D (signal_1302), .Q (signal_1886) ) ;
    buf_clk cell_1135 ( .C (clk), .D (signal_799), .Q (signal_1888) ) ;
    buf_clk cell_1137 ( .C (clk), .D (signal_1301), .Q (signal_1890) ) ;
    buf_clk cell_1139 ( .C (clk), .D (signal_800), .Q (signal_1892) ) ;
    buf_clk cell_1141 ( .C (clk), .D (signal_1397), .Q (signal_1894) ) ;
    buf_clk cell_1143 ( .C (clk), .D (signal_801), .Q (signal_1896) ) ;
    buf_clk cell_1145 ( .C (clk), .D (signal_1396), .Q (signal_1898) ) ;
    buf_clk cell_1147 ( .C (clk), .D (signal_802), .Q (signal_1900) ) ;
    buf_clk cell_1149 ( .C (clk), .D (signal_1395), .Q (signal_1902) ) ;
    buf_clk cell_1151 ( .C (clk), .D (signal_803), .Q (signal_1904) ) ;
    buf_clk cell_1153 ( .C (clk), .D (signal_1394), .Q (signal_1906) ) ;
    buf_clk cell_1155 ( .C (clk), .D (signal_804), .Q (signal_1908) ) ;
    buf_clk cell_1157 ( .C (clk), .D (signal_1401), .Q (signal_1910) ) ;
    buf_clk cell_1159 ( .C (clk), .D (signal_805), .Q (signal_1912) ) ;
    buf_clk cell_1161 ( .C (clk), .D (signal_1400), .Q (signal_1914) ) ;
    buf_clk cell_1163 ( .C (clk), .D (signal_806), .Q (signal_1916) ) ;
    buf_clk cell_1165 ( .C (clk), .D (signal_1399), .Q (signal_1918) ) ;
    buf_clk cell_1167 ( .C (clk), .D (signal_807), .Q (signal_1920) ) ;
    buf_clk cell_1169 ( .C (clk), .D (signal_1398), .Q (signal_1922) ) ;
    buf_clk cell_1171 ( .C (clk), .D (signal_808), .Q (signal_1924) ) ;
    buf_clk cell_1173 ( .C (clk), .D (signal_1405), .Q (signal_1926) ) ;
    buf_clk cell_1175 ( .C (clk), .D (signal_809), .Q (signal_1928) ) ;
    buf_clk cell_1177 ( .C (clk), .D (signal_1404), .Q (signal_1930) ) ;
    buf_clk cell_1179 ( .C (clk), .D (signal_810), .Q (signal_1932) ) ;
    buf_clk cell_1181 ( .C (clk), .D (signal_1403), .Q (signal_1934) ) ;
    buf_clk cell_1183 ( .C (clk), .D (signal_811), .Q (signal_1936) ) ;
    buf_clk cell_1185 ( .C (clk), .D (signal_1402), .Q (signal_1938) ) ;
    buf_clk cell_1187 ( .C (clk), .D (signal_812), .Q (signal_1940) ) ;
    buf_clk cell_1189 ( .C (clk), .D (signal_1409), .Q (signal_1942) ) ;
    buf_clk cell_1191 ( .C (clk), .D (signal_813), .Q (signal_1944) ) ;
    buf_clk cell_1193 ( .C (clk), .D (signal_1408), .Q (signal_1946) ) ;
    buf_clk cell_1195 ( .C (clk), .D (signal_814), .Q (signal_1948) ) ;
    buf_clk cell_1197 ( .C (clk), .D (signal_1407), .Q (signal_1950) ) ;
    buf_clk cell_1199 ( .C (clk), .D (signal_815), .Q (signal_1952) ) ;
    buf_clk cell_1201 ( .C (clk), .D (signal_1406), .Q (signal_1954) ) ;
    buf_clk cell_1203 ( .C (clk), .D (signal_816), .Q (signal_1956) ) ;
    buf_clk cell_1205 ( .C (clk), .D (signal_1413), .Q (signal_1958) ) ;
    buf_clk cell_1207 ( .C (clk), .D (signal_817), .Q (signal_1960) ) ;
    buf_clk cell_1209 ( .C (clk), .D (signal_1412), .Q (signal_1962) ) ;
    buf_clk cell_1211 ( .C (clk), .D (signal_818), .Q (signal_1964) ) ;
    buf_clk cell_1213 ( .C (clk), .D (signal_1411), .Q (signal_1966) ) ;
    buf_clk cell_1215 ( .C (clk), .D (signal_819), .Q (signal_1968) ) ;
    buf_clk cell_1217 ( .C (clk), .D (signal_1410), .Q (signal_1970) ) ;
    buf_clk cell_1219 ( .C (clk), .D (signal_820), .Q (signal_1972) ) ;
    buf_clk cell_1221 ( .C (clk), .D (signal_1417), .Q (signal_1974) ) ;
    buf_clk cell_1223 ( .C (clk), .D (signal_821), .Q (signal_1976) ) ;
    buf_clk cell_1225 ( .C (clk), .D (signal_1416), .Q (signal_1978) ) ;
    buf_clk cell_1227 ( .C (clk), .D (signal_822), .Q (signal_1980) ) ;
    buf_clk cell_1229 ( .C (clk), .D (signal_1415), .Q (signal_1982) ) ;
    buf_clk cell_1231 ( .C (clk), .D (signal_823), .Q (signal_1984) ) ;
    buf_clk cell_1233 ( .C (clk), .D (signal_1414), .Q (signal_1986) ) ;
    buf_clk cell_1235 ( .C (clk), .D (signal_824), .Q (signal_1988) ) ;
    buf_clk cell_1237 ( .C (clk), .D (signal_1421), .Q (signal_1990) ) ;
    buf_clk cell_1239 ( .C (clk), .D (signal_825), .Q (signal_1992) ) ;
    buf_clk cell_1241 ( .C (clk), .D (signal_1420), .Q (signal_1994) ) ;
    buf_clk cell_1243 ( .C (clk), .D (signal_826), .Q (signal_1996) ) ;
    buf_clk cell_1245 ( .C (clk), .D (signal_1419), .Q (signal_1998) ) ;
    buf_clk cell_1247 ( .C (clk), .D (signal_827), .Q (signal_2000) ) ;
    buf_clk cell_1249 ( .C (clk), .D (signal_1418), .Q (signal_2002) ) ;
    buf_clk cell_1251 ( .C (clk), .D (signal_828), .Q (signal_2004) ) ;
    buf_clk cell_1253 ( .C (clk), .D (signal_1425), .Q (signal_2006) ) ;
    buf_clk cell_1255 ( .C (clk), .D (signal_829), .Q (signal_2008) ) ;
    buf_clk cell_1257 ( .C (clk), .D (signal_1424), .Q (signal_2010) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_830), .Q (signal_2012) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_1423), .Q (signal_2014) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_831), .Q (signal_2016) ) ;
    buf_clk cell_1265 ( .C (clk), .D (signal_1422), .Q (signal_2018) ) ;
    buf_clk cell_1267 ( .C (clk), .D (signal_832), .Q (signal_2020) ) ;
    buf_clk cell_1269 ( .C (clk), .D (signal_1429), .Q (signal_2022) ) ;
    buf_clk cell_1271 ( .C (clk), .D (signal_833), .Q (signal_2024) ) ;
    buf_clk cell_1273 ( .C (clk), .D (signal_1428), .Q (signal_2026) ) ;
    buf_clk cell_1275 ( .C (clk), .D (signal_834), .Q (signal_2028) ) ;
    buf_clk cell_1277 ( .C (clk), .D (signal_1427), .Q (signal_2030) ) ;
    buf_clk cell_1279 ( .C (clk), .D (signal_835), .Q (signal_2032) ) ;
    buf_clk cell_1281 ( .C (clk), .D (signal_1426), .Q (signal_2034) ) ;
    buf_clk cell_1283 ( .C (clk), .D (signal_836), .Q (signal_2036) ) ;
    buf_clk cell_1285 ( .C (clk), .D (signal_1433), .Q (signal_2038) ) ;
    buf_clk cell_1287 ( .C (clk), .D (signal_837), .Q (signal_2040) ) ;
    buf_clk cell_1289 ( .C (clk), .D (signal_1432), .Q (signal_2042) ) ;
    buf_clk cell_1291 ( .C (clk), .D (signal_838), .Q (signal_2044) ) ;
    buf_clk cell_1293 ( .C (clk), .D (signal_1431), .Q (signal_2046) ) ;
    buf_clk cell_1295 ( .C (clk), .D (signal_839), .Q (signal_2048) ) ;
    buf_clk cell_1297 ( .C (clk), .D (signal_1430), .Q (signal_2050) ) ;
    buf_clk cell_1299 ( .C (clk), .D (signal_840), .Q (signal_2052) ) ;
    buf_clk cell_1301 ( .C (clk), .D (signal_1437), .Q (signal_2054) ) ;
    buf_clk cell_1303 ( .C (clk), .D (signal_841), .Q (signal_2056) ) ;
    buf_clk cell_1305 ( .C (clk), .D (signal_1436), .Q (signal_2058) ) ;
    buf_clk cell_1307 ( .C (clk), .D (signal_842), .Q (signal_2060) ) ;
    buf_clk cell_1309 ( .C (clk), .D (signal_1435), .Q (signal_2062) ) ;
    buf_clk cell_1311 ( .C (clk), .D (signal_843), .Q (signal_2064) ) ;
    buf_clk cell_1313 ( .C (clk), .D (signal_1434), .Q (signal_2066) ) ;
    buf_clk cell_1315 ( .C (clk), .D (signal_844), .Q (signal_2068) ) ;
    buf_clk cell_1317 ( .C (clk), .D (signal_1441), .Q (signal_2070) ) ;
    buf_clk cell_1319 ( .C (clk), .D (signal_845), .Q (signal_2072) ) ;
    buf_clk cell_1321 ( .C (clk), .D (signal_1440), .Q (signal_2074) ) ;
    buf_clk cell_1323 ( .C (clk), .D (signal_846), .Q (signal_2076) ) ;
    buf_clk cell_1325 ( .C (clk), .D (signal_1439), .Q (signal_2078) ) ;
    buf_clk cell_1327 ( .C (clk), .D (signal_847), .Q (signal_2080) ) ;
    buf_clk cell_1329 ( .C (clk), .D (signal_1438), .Q (signal_2082) ) ;
    buf_clk cell_1331 ( .C (clk), .D (signal_848), .Q (signal_2084) ) ;
    buf_clk cell_1333 ( .C (clk), .D (signal_1445), .Q (signal_2086) ) ;
    buf_clk cell_1335 ( .C (clk), .D (signal_849), .Q (signal_2088) ) ;
    buf_clk cell_1337 ( .C (clk), .D (signal_1444), .Q (signal_2090) ) ;
    buf_clk cell_1339 ( .C (clk), .D (signal_850), .Q (signal_2092) ) ;
    buf_clk cell_1341 ( .C (clk), .D (signal_1443), .Q (signal_2094) ) ;
    buf_clk cell_1343 ( .C (clk), .D (signal_851), .Q (signal_2096) ) ;
    buf_clk cell_1345 ( .C (clk), .D (signal_1442), .Q (signal_2098) ) ;

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_89 ( .s (signal_1459), .b ({signal_1316, signal_466}), .a ({signal_1463, signal_1461}), .c ({signal_1319, signal_557}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_90 ( .s (signal_1459), .b ({signal_1317, signal_465}), .a ({signal_1467, signal_1465}), .c ({signal_1320, signal_556}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_91 ( .s (signal_1459), .b ({signal_1318, signal_464}), .a ({signal_1471, signal_1469}), .c ({signal_1321, signal_555}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_92 ( .s (signal_1459), .b ({signal_1451, signal_463}), .a ({signal_1475, signal_1473}), .c ({signal_1452, signal_554}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_589 ( .s (signal_1477), .b ({signal_1481, signal_1479}), .a ({signal_1310, signal_699}), .c ({signal_1446, signal_855}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_590 ( .s (signal_1477), .b ({signal_1485, signal_1483}), .a ({signal_1312, signal_698}), .c ({signal_1447, signal_854}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_591 ( .s (signal_1477), .b ({signal_1489, signal_1487}), .a ({signal_1314, signal_697}), .c ({signal_1448, signal_853}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_592 ( .s (signal_1477), .b ({signal_1493, signal_1491}), .a ({signal_1450, signal_696}), .c ({signal_1453, signal_852}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_669 ( .s (signal_1495), .b ({signal_1308, signal_470}), .a ({signal_1499, signal_1497}), .c ({signal_1310, signal_699}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_670 ( .s (signal_1495), .b ({signal_1307, signal_469}), .a ({signal_1503, signal_1501}), .c ({signal_1312, signal_698}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_671 ( .s (signal_1495), .b ({signal_1306, signal_468}), .a ({signal_1507, signal_1505}), .c ({signal_1314, signal_697}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_672 ( .s (signal_1495), .b ({signal_1315, signal_467}), .a ({signal_1511, signal_1509}), .c ({signal_1450, signal_696}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_691 ( .a ({signal_1515, signal_1513}), .b ({signal_1305, signal_443}), .c ({signal_1315, signal_467}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_700 ( .s (signal_1517), .b ({signal_1308, signal_470}), .a ({signal_1521, signal_1519}), .c ({signal_1316, signal_466}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_701 ( .s (signal_1517), .b ({signal_1307, signal_469}), .a ({signal_1525, signal_1523}), .c ({signal_1317, signal_465}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_702 ( .s (signal_1517), .b ({signal_1306, signal_468}), .a ({signal_1529, signal_1527}), .c ({signal_1318, signal_464}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_703 ( .s (signal_1517), .b ({signal_1315, signal_467}), .a ({signal_1533, signal_1531}), .c ({signal_1451, signal_463}) ) ;
    PRESENT_step2_ANF #(.low_latency(0), .pipeline(1)) cell_704 ( .in0 ({signal_481, signal_480, signal_479, signal_478}), .in1 ({signal_1286, signal_1288, signal_1290, signal_1292}), .clk (clk), .r ({Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_470, signal_469, signal_468, signal_443}), .out1 ({signal_1308, signal_1307, signal_1306, signal_1305}) ) ;
    buf_clk cell_706 ( .C (clk), .D (signal_1458), .Q (signal_1459) ) ;
    buf_clk cell_708 ( .C (clk), .D (signal_1460), .Q (signal_1461) ) ;
    buf_clk cell_710 ( .C (clk), .D (signal_1462), .Q (signal_1463) ) ;
    buf_clk cell_712 ( .C (clk), .D (signal_1464), .Q (signal_1465) ) ;
    buf_clk cell_714 ( .C (clk), .D (signal_1466), .Q (signal_1467) ) ;
    buf_clk cell_716 ( .C (clk), .D (signal_1468), .Q (signal_1469) ) ;
    buf_clk cell_718 ( .C (clk), .D (signal_1470), .Q (signal_1471) ) ;
    buf_clk cell_720 ( .C (clk), .D (signal_1472), .Q (signal_1473) ) ;
    buf_clk cell_722 ( .C (clk), .D (signal_1474), .Q (signal_1475) ) ;
    buf_clk cell_724 ( .C (clk), .D (signal_1476), .Q (signal_1477) ) ;
    buf_clk cell_726 ( .C (clk), .D (signal_1478), .Q (signal_1479) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_1480), .Q (signal_1481) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_1482), .Q (signal_1483) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_1484), .Q (signal_1485) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_1486), .Q (signal_1487) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_1488), .Q (signal_1489) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_1490), .Q (signal_1491) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_1492), .Q (signal_1493) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_1494), .Q (signal_1495) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_1496), .Q (signal_1497) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_1498), .Q (signal_1499) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_1500), .Q (signal_1501) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_1502), .Q (signal_1503) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_1504), .Q (signal_1505) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_1506), .Q (signal_1507) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_1508), .Q (signal_1509) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_1510), .Q (signal_1511) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_1512), .Q (signal_1513) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_1514), .Q (signal_1515) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_1516), .Q (signal_1517) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_1518), .Q (signal_1519) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_1520), .Q (signal_1521) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_1522), .Q (signal_1523) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_1524), .Q (signal_1525) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_1526), .Q (signal_1527) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_1528), .Q (signal_1529) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_1530), .Q (signal_1531) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_1532), .Q (signal_1533) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_1534), .Q (signal_1535) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_1536), .Q (signal_1537) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_1538), .Q (signal_1539) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_1540), .Q (signal_1541) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_1542), .Q (signal_1543) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_1544), .Q (signal_1545) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_1546), .Q (signal_1547) ) ;
    buf_clk cell_796 ( .C (clk), .D (signal_1548), .Q (signal_1549) ) ;
    buf_clk cell_798 ( .C (clk), .D (signal_1550), .Q (signal_1551) ) ;
    buf_clk cell_800 ( .C (clk), .D (signal_1552), .Q (signal_1553) ) ;
    buf_clk cell_802 ( .C (clk), .D (signal_1554), .Q (signal_1555) ) ;
    buf_clk cell_804 ( .C (clk), .D (signal_1556), .Q (signal_1557) ) ;
    buf_clk cell_806 ( .C (clk), .D (signal_1558), .Q (signal_1559) ) ;
    buf_clk cell_808 ( .C (clk), .D (signal_1560), .Q (signal_1561) ) ;
    buf_clk cell_810 ( .C (clk), .D (signal_1562), .Q (signal_1563) ) ;
    buf_clk cell_812 ( .C (clk), .D (signal_1564), .Q (signal_1565) ) ;
    buf_clk cell_814 ( .C (clk), .D (signal_1566), .Q (signal_1567) ) ;
    buf_clk cell_816 ( .C (clk), .D (signal_1568), .Q (signal_1569) ) ;
    buf_clk cell_818 ( .C (clk), .D (signal_1570), .Q (signal_1571) ) ;
    buf_clk cell_820 ( .C (clk), .D (signal_1572), .Q (signal_1573) ) ;
    buf_clk cell_822 ( .C (clk), .D (signal_1574), .Q (signal_1575) ) ;
    buf_clk cell_824 ( .C (clk), .D (signal_1576), .Q (signal_1577) ) ;
    buf_clk cell_826 ( .C (clk), .D (signal_1578), .Q (signal_1579) ) ;
    buf_clk cell_828 ( .C (clk), .D (signal_1580), .Q (signal_1581) ) ;
    buf_clk cell_830 ( .C (clk), .D (signal_1582), .Q (signal_1583) ) ;
    buf_clk cell_832 ( .C (clk), .D (signal_1584), .Q (signal_1585) ) ;
    buf_clk cell_834 ( .C (clk), .D (signal_1586), .Q (signal_1587) ) ;
    buf_clk cell_836 ( .C (clk), .D (signal_1588), .Q (signal_1589) ) ;
    buf_clk cell_838 ( .C (clk), .D (signal_1590), .Q (signal_1591) ) ;
    buf_clk cell_840 ( .C (clk), .D (signal_1592), .Q (signal_1593) ) ;
    buf_clk cell_842 ( .C (clk), .D (signal_1594), .Q (signal_1595) ) ;
    buf_clk cell_844 ( .C (clk), .D (signal_1596), .Q (signal_1597) ) ;
    buf_clk cell_846 ( .C (clk), .D (signal_1598), .Q (signal_1599) ) ;
    buf_clk cell_848 ( .C (clk), .D (signal_1600), .Q (signal_1601) ) ;
    buf_clk cell_850 ( .C (clk), .D (signal_1602), .Q (signal_1603) ) ;
    buf_clk cell_852 ( .C (clk), .D (signal_1604), .Q (signal_1605) ) ;
    buf_clk cell_854 ( .C (clk), .D (signal_1606), .Q (signal_1607) ) ;
    buf_clk cell_856 ( .C (clk), .D (signal_1608), .Q (signal_1609) ) ;
    buf_clk cell_858 ( .C (clk), .D (signal_1610), .Q (signal_1611) ) ;
    buf_clk cell_860 ( .C (clk), .D (signal_1612), .Q (signal_1613) ) ;
    buf_clk cell_862 ( .C (clk), .D (signal_1614), .Q (signal_1615) ) ;
    buf_clk cell_864 ( .C (clk), .D (signal_1616), .Q (signal_1617) ) ;
    buf_clk cell_866 ( .C (clk), .D (signal_1618), .Q (signal_1619) ) ;
    buf_clk cell_868 ( .C (clk), .D (signal_1620), .Q (signal_1621) ) ;
    buf_clk cell_870 ( .C (clk), .D (signal_1622), .Q (signal_1623) ) ;
    buf_clk cell_872 ( .C (clk), .D (signal_1624), .Q (signal_1625) ) ;
    buf_clk cell_874 ( .C (clk), .D (signal_1626), .Q (signal_1627) ) ;
    buf_clk cell_876 ( .C (clk), .D (signal_1628), .Q (signal_1629) ) ;
    buf_clk cell_878 ( .C (clk), .D (signal_1630), .Q (signal_1631) ) ;
    buf_clk cell_880 ( .C (clk), .D (signal_1632), .Q (signal_1633) ) ;
    buf_clk cell_882 ( .C (clk), .D (signal_1634), .Q (signal_1635) ) ;
    buf_clk cell_884 ( .C (clk), .D (signal_1636), .Q (signal_1637) ) ;
    buf_clk cell_886 ( .C (clk), .D (signal_1638), .Q (signal_1639) ) ;
    buf_clk cell_888 ( .C (clk), .D (signal_1640), .Q (signal_1641) ) ;
    buf_clk cell_890 ( .C (clk), .D (signal_1642), .Q (signal_1643) ) ;
    buf_clk cell_892 ( .C (clk), .D (signal_1644), .Q (signal_1645) ) ;
    buf_clk cell_894 ( .C (clk), .D (signal_1646), .Q (signal_1647) ) ;
    buf_clk cell_896 ( .C (clk), .D (signal_1648), .Q (signal_1649) ) ;
    buf_clk cell_898 ( .C (clk), .D (signal_1650), .Q (signal_1651) ) ;
    buf_clk cell_900 ( .C (clk), .D (signal_1652), .Q (signal_1653) ) ;
    buf_clk cell_902 ( .C (clk), .D (signal_1654), .Q (signal_1655) ) ;
    buf_clk cell_904 ( .C (clk), .D (signal_1656), .Q (signal_1657) ) ;
    buf_clk cell_906 ( .C (clk), .D (signal_1658), .Q (signal_1659) ) ;
    buf_clk cell_908 ( .C (clk), .D (signal_1660), .Q (signal_1661) ) ;
    buf_clk cell_910 ( .C (clk), .D (signal_1662), .Q (signal_1663) ) ;
    buf_clk cell_912 ( .C (clk), .D (signal_1664), .Q (signal_1665) ) ;
    buf_clk cell_914 ( .C (clk), .D (signal_1666), .Q (signal_1667) ) ;
    buf_clk cell_916 ( .C (clk), .D (signal_1668), .Q (signal_1669) ) ;
    buf_clk cell_918 ( .C (clk), .D (signal_1670), .Q (signal_1671) ) ;
    buf_clk cell_920 ( .C (clk), .D (signal_1672), .Q (signal_1673) ) ;
    buf_clk cell_922 ( .C (clk), .D (signal_1674), .Q (signal_1675) ) ;
    buf_clk cell_924 ( .C (clk), .D (signal_1676), .Q (signal_1677) ) ;
    buf_clk cell_926 ( .C (clk), .D (signal_1678), .Q (signal_1679) ) ;
    buf_clk cell_928 ( .C (clk), .D (signal_1680), .Q (signal_1681) ) ;
    buf_clk cell_930 ( .C (clk), .D (signal_1682), .Q (signal_1683) ) ;
    buf_clk cell_932 ( .C (clk), .D (signal_1684), .Q (signal_1685) ) ;
    buf_clk cell_934 ( .C (clk), .D (signal_1686), .Q (signal_1687) ) ;
    buf_clk cell_936 ( .C (clk), .D (signal_1688), .Q (signal_1689) ) ;
    buf_clk cell_938 ( .C (clk), .D (signal_1690), .Q (signal_1691) ) ;
    buf_clk cell_940 ( .C (clk), .D (signal_1692), .Q (signal_1693) ) ;
    buf_clk cell_942 ( .C (clk), .D (signal_1694), .Q (signal_1695) ) ;
    buf_clk cell_944 ( .C (clk), .D (signal_1696), .Q (signal_1697) ) ;
    buf_clk cell_946 ( .C (clk), .D (signal_1698), .Q (signal_1699) ) ;
    buf_clk cell_948 ( .C (clk), .D (signal_1700), .Q (signal_1701) ) ;
    buf_clk cell_950 ( .C (clk), .D (signal_1702), .Q (signal_1703) ) ;
    buf_clk cell_952 ( .C (clk), .D (signal_1704), .Q (signal_1705) ) ;
    buf_clk cell_954 ( .C (clk), .D (signal_1706), .Q (signal_1707) ) ;
    buf_clk cell_956 ( .C (clk), .D (signal_1708), .Q (signal_1709) ) ;
    buf_clk cell_958 ( .C (clk), .D (signal_1710), .Q (signal_1711) ) ;
    buf_clk cell_960 ( .C (clk), .D (signal_1712), .Q (signal_1713) ) ;
    buf_clk cell_962 ( .C (clk), .D (signal_1714), .Q (signal_1715) ) ;
    buf_clk cell_964 ( .C (clk), .D (signal_1716), .Q (signal_1717) ) ;
    buf_clk cell_966 ( .C (clk), .D (signal_1718), .Q (signal_1719) ) ;
    buf_clk cell_968 ( .C (clk), .D (signal_1720), .Q (signal_1721) ) ;
    buf_clk cell_970 ( .C (clk), .D (signal_1722), .Q (signal_1723) ) ;
    buf_clk cell_972 ( .C (clk), .D (signal_1724), .Q (signal_1725) ) ;
    buf_clk cell_974 ( .C (clk), .D (signal_1726), .Q (signal_1727) ) ;
    buf_clk cell_976 ( .C (clk), .D (signal_1728), .Q (signal_1729) ) ;
    buf_clk cell_978 ( .C (clk), .D (signal_1730), .Q (signal_1731) ) ;
    buf_clk cell_980 ( .C (clk), .D (signal_1732), .Q (signal_1733) ) ;
    buf_clk cell_982 ( .C (clk), .D (signal_1734), .Q (signal_1735) ) ;
    buf_clk cell_984 ( .C (clk), .D (signal_1736), .Q (signal_1737) ) ;
    buf_clk cell_986 ( .C (clk), .D (signal_1738), .Q (signal_1739) ) ;
    buf_clk cell_988 ( .C (clk), .D (signal_1740), .Q (signal_1741) ) ;
    buf_clk cell_990 ( .C (clk), .D (signal_1742), .Q (signal_1743) ) ;
    buf_clk cell_992 ( .C (clk), .D (signal_1744), .Q (signal_1745) ) ;
    buf_clk cell_994 ( .C (clk), .D (signal_1746), .Q (signal_1747) ) ;
    buf_clk cell_996 ( .C (clk), .D (signal_1748), .Q (signal_1749) ) ;
    buf_clk cell_998 ( .C (clk), .D (signal_1750), .Q (signal_1751) ) ;
    buf_clk cell_1000 ( .C (clk), .D (signal_1752), .Q (signal_1753) ) ;
    buf_clk cell_1002 ( .C (clk), .D (signal_1754), .Q (signal_1755) ) ;
    buf_clk cell_1004 ( .C (clk), .D (signal_1756), .Q (signal_1757) ) ;
    buf_clk cell_1006 ( .C (clk), .D (signal_1758), .Q (signal_1759) ) ;
    buf_clk cell_1008 ( .C (clk), .D (signal_1760), .Q (signal_1761) ) ;
    buf_clk cell_1010 ( .C (clk), .D (signal_1762), .Q (signal_1763) ) ;
    buf_clk cell_1012 ( .C (clk), .D (signal_1764), .Q (signal_1765) ) ;
    buf_clk cell_1014 ( .C (clk), .D (signal_1766), .Q (signal_1767) ) ;
    buf_clk cell_1016 ( .C (clk), .D (signal_1768), .Q (signal_1769) ) ;
    buf_clk cell_1018 ( .C (clk), .D (signal_1770), .Q (signal_1771) ) ;
    buf_clk cell_1020 ( .C (clk), .D (signal_1772), .Q (signal_1773) ) ;
    buf_clk cell_1022 ( .C (clk), .D (signal_1774), .Q (signal_1775) ) ;
    buf_clk cell_1024 ( .C (clk), .D (signal_1776), .Q (signal_1777) ) ;
    buf_clk cell_1026 ( .C (clk), .D (signal_1778), .Q (signal_1779) ) ;
    buf_clk cell_1028 ( .C (clk), .D (signal_1780), .Q (signal_1781) ) ;
    buf_clk cell_1030 ( .C (clk), .D (signal_1782), .Q (signal_1783) ) ;
    buf_clk cell_1032 ( .C (clk), .D (signal_1784), .Q (signal_1785) ) ;
    buf_clk cell_1034 ( .C (clk), .D (signal_1786), .Q (signal_1787) ) ;
    buf_clk cell_1036 ( .C (clk), .D (signal_1788), .Q (signal_1789) ) ;
    buf_clk cell_1038 ( .C (clk), .D (signal_1790), .Q (signal_1791) ) ;
    buf_clk cell_1040 ( .C (clk), .D (signal_1792), .Q (signal_1793) ) ;
    buf_clk cell_1042 ( .C (clk), .D (signal_1794), .Q (signal_1795) ) ;
    buf_clk cell_1044 ( .C (clk), .D (signal_1796), .Q (signal_1797) ) ;
    buf_clk cell_1046 ( .C (clk), .D (signal_1798), .Q (signal_1799) ) ;
    buf_clk cell_1048 ( .C (clk), .D (signal_1800), .Q (signal_1801) ) ;
    buf_clk cell_1050 ( .C (clk), .D (signal_1802), .Q (signal_1803) ) ;
    buf_clk cell_1052 ( .C (clk), .D (signal_1804), .Q (signal_1805) ) ;
    buf_clk cell_1054 ( .C (clk), .D (signal_1806), .Q (signal_1807) ) ;
    buf_clk cell_1056 ( .C (clk), .D (signal_1808), .Q (signal_1809) ) ;
    buf_clk cell_1058 ( .C (clk), .D (signal_1810), .Q (signal_1811) ) ;
    buf_clk cell_1060 ( .C (clk), .D (signal_1812), .Q (signal_1813) ) ;
    buf_clk cell_1062 ( .C (clk), .D (signal_1814), .Q (signal_1815) ) ;
    buf_clk cell_1064 ( .C (clk), .D (signal_1816), .Q (signal_1817) ) ;
    buf_clk cell_1066 ( .C (clk), .D (signal_1818), .Q (signal_1819) ) ;
    buf_clk cell_1068 ( .C (clk), .D (signal_1820), .Q (signal_1821) ) ;
    buf_clk cell_1070 ( .C (clk), .D (signal_1822), .Q (signal_1823) ) ;
    buf_clk cell_1072 ( .C (clk), .D (signal_1824), .Q (signal_1825) ) ;
    buf_clk cell_1074 ( .C (clk), .D (signal_1826), .Q (signal_1827) ) ;
    buf_clk cell_1076 ( .C (clk), .D (signal_1828), .Q (signal_1829) ) ;
    buf_clk cell_1078 ( .C (clk), .D (signal_1830), .Q (signal_1831) ) ;
    buf_clk cell_1080 ( .C (clk), .D (signal_1832), .Q (signal_1833) ) ;
    buf_clk cell_1082 ( .C (clk), .D (signal_1834), .Q (signal_1835) ) ;
    buf_clk cell_1084 ( .C (clk), .D (signal_1836), .Q (signal_1837) ) ;
    buf_clk cell_1086 ( .C (clk), .D (signal_1838), .Q (signal_1839) ) ;
    buf_clk cell_1088 ( .C (clk), .D (signal_1840), .Q (signal_1841) ) ;
    buf_clk cell_1090 ( .C (clk), .D (signal_1842), .Q (signal_1843) ) ;
    buf_clk cell_1092 ( .C (clk), .D (signal_1844), .Q (signal_1845) ) ;
    buf_clk cell_1094 ( .C (clk), .D (signal_1846), .Q (signal_1847) ) ;
    buf_clk cell_1096 ( .C (clk), .D (signal_1848), .Q (signal_1849) ) ;
    buf_clk cell_1098 ( .C (clk), .D (signal_1850), .Q (signal_1851) ) ;
    buf_clk cell_1100 ( .C (clk), .D (signal_1852), .Q (signal_1853) ) ;
    buf_clk cell_1102 ( .C (clk), .D (signal_1854), .Q (signal_1855) ) ;
    buf_clk cell_1104 ( .C (clk), .D (signal_1856), .Q (signal_1857) ) ;
    buf_clk cell_1106 ( .C (clk), .D (signal_1858), .Q (signal_1859) ) ;
    buf_clk cell_1108 ( .C (clk), .D (signal_1860), .Q (signal_1861) ) ;
    buf_clk cell_1110 ( .C (clk), .D (signal_1862), .Q (signal_1863) ) ;
    buf_clk cell_1112 ( .C (clk), .D (signal_1864), .Q (signal_1865) ) ;
    buf_clk cell_1114 ( .C (clk), .D (signal_1866), .Q (signal_1867) ) ;
    buf_clk cell_1116 ( .C (clk), .D (signal_1868), .Q (signal_1869) ) ;
    buf_clk cell_1118 ( .C (clk), .D (signal_1870), .Q (signal_1871) ) ;
    buf_clk cell_1120 ( .C (clk), .D (signal_1872), .Q (signal_1873) ) ;
    buf_clk cell_1122 ( .C (clk), .D (signal_1874), .Q (signal_1875) ) ;
    buf_clk cell_1124 ( .C (clk), .D (signal_1876), .Q (signal_1877) ) ;
    buf_clk cell_1126 ( .C (clk), .D (signal_1878), .Q (signal_1879) ) ;
    buf_clk cell_1128 ( .C (clk), .D (signal_1880), .Q (signal_1881) ) ;
    buf_clk cell_1130 ( .C (clk), .D (signal_1882), .Q (signal_1883) ) ;
    buf_clk cell_1132 ( .C (clk), .D (signal_1884), .Q (signal_1885) ) ;
    buf_clk cell_1134 ( .C (clk), .D (signal_1886), .Q (signal_1887) ) ;
    buf_clk cell_1136 ( .C (clk), .D (signal_1888), .Q (signal_1889) ) ;
    buf_clk cell_1138 ( .C (clk), .D (signal_1890), .Q (signal_1891) ) ;
    buf_clk cell_1140 ( .C (clk), .D (signal_1892), .Q (signal_1893) ) ;
    buf_clk cell_1142 ( .C (clk), .D (signal_1894), .Q (signal_1895) ) ;
    buf_clk cell_1144 ( .C (clk), .D (signal_1896), .Q (signal_1897) ) ;
    buf_clk cell_1146 ( .C (clk), .D (signal_1898), .Q (signal_1899) ) ;
    buf_clk cell_1148 ( .C (clk), .D (signal_1900), .Q (signal_1901) ) ;
    buf_clk cell_1150 ( .C (clk), .D (signal_1902), .Q (signal_1903) ) ;
    buf_clk cell_1152 ( .C (clk), .D (signal_1904), .Q (signal_1905) ) ;
    buf_clk cell_1154 ( .C (clk), .D (signal_1906), .Q (signal_1907) ) ;
    buf_clk cell_1156 ( .C (clk), .D (signal_1908), .Q (signal_1909) ) ;
    buf_clk cell_1158 ( .C (clk), .D (signal_1910), .Q (signal_1911) ) ;
    buf_clk cell_1160 ( .C (clk), .D (signal_1912), .Q (signal_1913) ) ;
    buf_clk cell_1162 ( .C (clk), .D (signal_1914), .Q (signal_1915) ) ;
    buf_clk cell_1164 ( .C (clk), .D (signal_1916), .Q (signal_1917) ) ;
    buf_clk cell_1166 ( .C (clk), .D (signal_1918), .Q (signal_1919) ) ;
    buf_clk cell_1168 ( .C (clk), .D (signal_1920), .Q (signal_1921) ) ;
    buf_clk cell_1170 ( .C (clk), .D (signal_1922), .Q (signal_1923) ) ;
    buf_clk cell_1172 ( .C (clk), .D (signal_1924), .Q (signal_1925) ) ;
    buf_clk cell_1174 ( .C (clk), .D (signal_1926), .Q (signal_1927) ) ;
    buf_clk cell_1176 ( .C (clk), .D (signal_1928), .Q (signal_1929) ) ;
    buf_clk cell_1178 ( .C (clk), .D (signal_1930), .Q (signal_1931) ) ;
    buf_clk cell_1180 ( .C (clk), .D (signal_1932), .Q (signal_1933) ) ;
    buf_clk cell_1182 ( .C (clk), .D (signal_1934), .Q (signal_1935) ) ;
    buf_clk cell_1184 ( .C (clk), .D (signal_1936), .Q (signal_1937) ) ;
    buf_clk cell_1186 ( .C (clk), .D (signal_1938), .Q (signal_1939) ) ;
    buf_clk cell_1188 ( .C (clk), .D (signal_1940), .Q (signal_1941) ) ;
    buf_clk cell_1190 ( .C (clk), .D (signal_1942), .Q (signal_1943) ) ;
    buf_clk cell_1192 ( .C (clk), .D (signal_1944), .Q (signal_1945) ) ;
    buf_clk cell_1194 ( .C (clk), .D (signal_1946), .Q (signal_1947) ) ;
    buf_clk cell_1196 ( .C (clk), .D (signal_1948), .Q (signal_1949) ) ;
    buf_clk cell_1198 ( .C (clk), .D (signal_1950), .Q (signal_1951) ) ;
    buf_clk cell_1200 ( .C (clk), .D (signal_1952), .Q (signal_1953) ) ;
    buf_clk cell_1202 ( .C (clk), .D (signal_1954), .Q (signal_1955) ) ;
    buf_clk cell_1204 ( .C (clk), .D (signal_1956), .Q (signal_1957) ) ;
    buf_clk cell_1206 ( .C (clk), .D (signal_1958), .Q (signal_1959) ) ;
    buf_clk cell_1208 ( .C (clk), .D (signal_1960), .Q (signal_1961) ) ;
    buf_clk cell_1210 ( .C (clk), .D (signal_1962), .Q (signal_1963) ) ;
    buf_clk cell_1212 ( .C (clk), .D (signal_1964), .Q (signal_1965) ) ;
    buf_clk cell_1214 ( .C (clk), .D (signal_1966), .Q (signal_1967) ) ;
    buf_clk cell_1216 ( .C (clk), .D (signal_1968), .Q (signal_1969) ) ;
    buf_clk cell_1218 ( .C (clk), .D (signal_1970), .Q (signal_1971) ) ;
    buf_clk cell_1220 ( .C (clk), .D (signal_1972), .Q (signal_1973) ) ;
    buf_clk cell_1222 ( .C (clk), .D (signal_1974), .Q (signal_1975) ) ;
    buf_clk cell_1224 ( .C (clk), .D (signal_1976), .Q (signal_1977) ) ;
    buf_clk cell_1226 ( .C (clk), .D (signal_1978), .Q (signal_1979) ) ;
    buf_clk cell_1228 ( .C (clk), .D (signal_1980), .Q (signal_1981) ) ;
    buf_clk cell_1230 ( .C (clk), .D (signal_1982), .Q (signal_1983) ) ;
    buf_clk cell_1232 ( .C (clk), .D (signal_1984), .Q (signal_1985) ) ;
    buf_clk cell_1234 ( .C (clk), .D (signal_1986), .Q (signal_1987) ) ;
    buf_clk cell_1236 ( .C (clk), .D (signal_1988), .Q (signal_1989) ) ;
    buf_clk cell_1238 ( .C (clk), .D (signal_1990), .Q (signal_1991) ) ;
    buf_clk cell_1240 ( .C (clk), .D (signal_1992), .Q (signal_1993) ) ;
    buf_clk cell_1242 ( .C (clk), .D (signal_1994), .Q (signal_1995) ) ;
    buf_clk cell_1244 ( .C (clk), .D (signal_1996), .Q (signal_1997) ) ;
    buf_clk cell_1246 ( .C (clk), .D (signal_1998), .Q (signal_1999) ) ;
    buf_clk cell_1248 ( .C (clk), .D (signal_2000), .Q (signal_2001) ) ;
    buf_clk cell_1250 ( .C (clk), .D (signal_2002), .Q (signal_2003) ) ;
    buf_clk cell_1252 ( .C (clk), .D (signal_2004), .Q (signal_2005) ) ;
    buf_clk cell_1254 ( .C (clk), .D (signal_2006), .Q (signal_2007) ) ;
    buf_clk cell_1256 ( .C (clk), .D (signal_2008), .Q (signal_2009) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_2010), .Q (signal_2011) ) ;
    buf_clk cell_1260 ( .C (clk), .D (signal_2012), .Q (signal_2013) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_2014), .Q (signal_2015) ) ;
    buf_clk cell_1264 ( .C (clk), .D (signal_2016), .Q (signal_2017) ) ;
    buf_clk cell_1266 ( .C (clk), .D (signal_2018), .Q (signal_2019) ) ;
    buf_clk cell_1268 ( .C (clk), .D (signal_2020), .Q (signal_2021) ) ;
    buf_clk cell_1270 ( .C (clk), .D (signal_2022), .Q (signal_2023) ) ;
    buf_clk cell_1272 ( .C (clk), .D (signal_2024), .Q (signal_2025) ) ;
    buf_clk cell_1274 ( .C (clk), .D (signal_2026), .Q (signal_2027) ) ;
    buf_clk cell_1276 ( .C (clk), .D (signal_2028), .Q (signal_2029) ) ;
    buf_clk cell_1278 ( .C (clk), .D (signal_2030), .Q (signal_2031) ) ;
    buf_clk cell_1280 ( .C (clk), .D (signal_2032), .Q (signal_2033) ) ;
    buf_clk cell_1282 ( .C (clk), .D (signal_2034), .Q (signal_2035) ) ;
    buf_clk cell_1284 ( .C (clk), .D (signal_2036), .Q (signal_2037) ) ;
    buf_clk cell_1286 ( .C (clk), .D (signal_2038), .Q (signal_2039) ) ;
    buf_clk cell_1288 ( .C (clk), .D (signal_2040), .Q (signal_2041) ) ;
    buf_clk cell_1290 ( .C (clk), .D (signal_2042), .Q (signal_2043) ) ;
    buf_clk cell_1292 ( .C (clk), .D (signal_2044), .Q (signal_2045) ) ;
    buf_clk cell_1294 ( .C (clk), .D (signal_2046), .Q (signal_2047) ) ;
    buf_clk cell_1296 ( .C (clk), .D (signal_2048), .Q (signal_2049) ) ;
    buf_clk cell_1298 ( .C (clk), .D (signal_2050), .Q (signal_2051) ) ;
    buf_clk cell_1300 ( .C (clk), .D (signal_2052), .Q (signal_2053) ) ;
    buf_clk cell_1302 ( .C (clk), .D (signal_2054), .Q (signal_2055) ) ;
    buf_clk cell_1304 ( .C (clk), .D (signal_2056), .Q (signal_2057) ) ;
    buf_clk cell_1306 ( .C (clk), .D (signal_2058), .Q (signal_2059) ) ;
    buf_clk cell_1308 ( .C (clk), .D (signal_2060), .Q (signal_2061) ) ;
    buf_clk cell_1310 ( .C (clk), .D (signal_2062), .Q (signal_2063) ) ;
    buf_clk cell_1312 ( .C (clk), .D (signal_2064), .Q (signal_2065) ) ;
    buf_clk cell_1314 ( .C (clk), .D (signal_2066), .Q (signal_2067) ) ;
    buf_clk cell_1316 ( .C (clk), .D (signal_2068), .Q (signal_2069) ) ;
    buf_clk cell_1318 ( .C (clk), .D (signal_2070), .Q (signal_2071) ) ;
    buf_clk cell_1320 ( .C (clk), .D (signal_2072), .Q (signal_2073) ) ;
    buf_clk cell_1322 ( .C (clk), .D (signal_2074), .Q (signal_2075) ) ;
    buf_clk cell_1324 ( .C (clk), .D (signal_2076), .Q (signal_2077) ) ;
    buf_clk cell_1326 ( .C (clk), .D (signal_2078), .Q (signal_2079) ) ;
    buf_clk cell_1328 ( .C (clk), .D (signal_2080), .Q (signal_2081) ) ;
    buf_clk cell_1330 ( .C (clk), .D (signal_2082), .Q (signal_2083) ) ;
    buf_clk cell_1332 ( .C (clk), .D (signal_2084), .Q (signal_2085) ) ;
    buf_clk cell_1334 ( .C (clk), .D (signal_2086), .Q (signal_2087) ) ;
    buf_clk cell_1336 ( .C (clk), .D (signal_2088), .Q (signal_2089) ) ;
    buf_clk cell_1338 ( .C (clk), .D (signal_2090), .Q (signal_2091) ) ;
    buf_clk cell_1340 ( .C (clk), .D (signal_2092), .Q (signal_2093) ) ;
    buf_clk cell_1342 ( .C (clk), .D (signal_2094), .Q (signal_2095) ) ;
    buf_clk cell_1344 ( .C (clk), .D (signal_2096), .Q (signal_2097) ) ;
    buf_clk cell_1346 ( .C (clk), .D (signal_2098), .Q (signal_2099) ) ;

    /* register cells */
    DFF_X1 cell_53 ( .CK (clk), .D (signal_1535), .Q (signal_458), .QN () ) ;
    DFF_X1 cell_55 ( .CK (clk), .D (signal_1537), .Q (signal_460), .QN () ) ;
    DFF_X1 cell_57 ( .CK (clk), .D (signal_1539), .Q (signal_462), .QN () ) ;
    DFF_X1 cell_59 ( .CK (clk), .D (signal_1541), .Q (signal_459), .QN () ) ;
    DFF_X1 cell_61 ( .CK (clk), .D (signal_1543), .Q (signal_265), .QN () ) ;
    DFF_X1 cell_75 ( .CK (clk), .D (signal_1545), .Q (signal_487), .QN () ) ;
    DFF_X1 cell_77 ( .CK (clk), .D (signal_1547), .Q (signal_489), .QN () ) ;
    DFF_X1 cell_79 ( .CK (clk), .D (signal_1549), .Q (signal_486), .QN () ) ;
    DFF_X1 cell_81 ( .CK (clk), .D (signal_1551), .Q (signal_488), .QN () ) ;
    DFF_X1 cell_83 ( .CK (clk), .D (signal_1553), .Q (signal_234), .QN () ) ;
    DFF_X1 cell_85 ( .CK (clk), .D (signal_1555), .Q (signal_235), .QN () ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_94 ( .clk (clk), .D ({signal_1319, signal_557}), .Q ({data_out_s1[0], data_out_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_96 ( .clk (clk), .D ({signal_1321, signal_555}), .Q ({data_out_s1[2], data_out_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_98 ( .clk (clk), .D ({signal_1320, signal_556}), .Q ({data_out_s1[1], data_out_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_100 ( .clk (clk), .D ({signal_1452, signal_554}), .Q ({data_out_s1[3], data_out_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_102 ( .clk (clk), .D ({signal_1559, signal_1557}), .Q ({data_out_s1[7], data_out_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_104 ( .clk (clk), .D ({signal_1563, signal_1561}), .Q ({data_out_s1[6], data_out_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_106 ( .clk (clk), .D ({signal_1567, signal_1565}), .Q ({data_out_s1[5], data_out_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_108 ( .clk (clk), .D ({signal_1571, signal_1569}), .Q ({data_out_s1[4], data_out_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_114 ( .clk (clk), .D ({signal_1575, signal_1573}), .Q ({data_out_s1[11], data_out_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_116 ( .clk (clk), .D ({signal_1579, signal_1577}), .Q ({data_out_s1[10], data_out_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_118 ( .clk (clk), .D ({signal_1583, signal_1581}), .Q ({data_out_s1[9], data_out_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_120 ( .clk (clk), .D ({signal_1587, signal_1585}), .Q ({data_out_s1[8], data_out_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_126 ( .clk (clk), .D ({signal_1591, signal_1589}), .Q ({data_out_s1[15], data_out_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_128 ( .clk (clk), .D ({signal_1595, signal_1593}), .Q ({data_out_s1[14], data_out_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_130 ( .clk (clk), .D ({signal_1599, signal_1597}), .Q ({data_out_s1[13], data_out_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_132 ( .clk (clk), .D ({signal_1603, signal_1601}), .Q ({data_out_s1[12], data_out_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_138 ( .clk (clk), .D ({signal_1607, signal_1605}), .Q ({data_out_s1[19], data_out_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_140 ( .clk (clk), .D ({signal_1611, signal_1609}), .Q ({data_out_s1[18], data_out_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_142 ( .clk (clk), .D ({signal_1615, signal_1613}), .Q ({data_out_s1[17], data_out_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_144 ( .clk (clk), .D ({signal_1619, signal_1617}), .Q ({data_out_s1[16], data_out_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_150 ( .clk (clk), .D ({signal_1623, signal_1621}), .Q ({data_out_s1[23], data_out_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_152 ( .clk (clk), .D ({signal_1627, signal_1625}), .Q ({data_out_s1[22], data_out_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_154 ( .clk (clk), .D ({signal_1631, signal_1629}), .Q ({data_out_s1[21], data_out_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_156 ( .clk (clk), .D ({signal_1635, signal_1633}), .Q ({data_out_s1[20], data_out_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_162 ( .clk (clk), .D ({signal_1639, signal_1637}), .Q ({data_out_s1[27], data_out_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_164 ( .clk (clk), .D ({signal_1643, signal_1641}), .Q ({data_out_s1[26], data_out_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_166 ( .clk (clk), .D ({signal_1647, signal_1645}), .Q ({data_out_s1[25], data_out_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_168 ( .clk (clk), .D ({signal_1651, signal_1649}), .Q ({data_out_s1[24], data_out_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_174 ( .clk (clk), .D ({signal_1655, signal_1653}), .Q ({data_out_s1[31], data_out_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_176 ( .clk (clk), .D ({signal_1659, signal_1657}), .Q ({data_out_s1[30], data_out_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_178 ( .clk (clk), .D ({signal_1663, signal_1661}), .Q ({data_out_s1[29], data_out_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_180 ( .clk (clk), .D ({signal_1667, signal_1665}), .Q ({data_out_s1[28], data_out_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_186 ( .clk (clk), .D ({signal_1671, signal_1669}), .Q ({data_out_s1[35], data_out_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_188 ( .clk (clk), .D ({signal_1675, signal_1673}), .Q ({data_out_s1[34], data_out_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_190 ( .clk (clk), .D ({signal_1679, signal_1677}), .Q ({data_out_s1[33], data_out_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_192 ( .clk (clk), .D ({signal_1683, signal_1681}), .Q ({data_out_s1[32], data_out_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_198 ( .clk (clk), .D ({signal_1687, signal_1685}), .Q ({data_out_s1[39], data_out_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_200 ( .clk (clk), .D ({signal_1691, signal_1689}), .Q ({data_out_s1[38], data_out_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_202 ( .clk (clk), .D ({signal_1695, signal_1693}), .Q ({data_out_s1[37], data_out_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_204 ( .clk (clk), .D ({signal_1699, signal_1697}), .Q ({data_out_s1[36], data_out_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_210 ( .clk (clk), .D ({signal_1703, signal_1701}), .Q ({data_out_s1[43], data_out_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_212 ( .clk (clk), .D ({signal_1707, signal_1705}), .Q ({data_out_s1[42], data_out_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_214 ( .clk (clk), .D ({signal_1711, signal_1709}), .Q ({data_out_s1[41], data_out_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_216 ( .clk (clk), .D ({signal_1715, signal_1713}), .Q ({data_out_s1[40], data_out_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_222 ( .clk (clk), .D ({signal_1719, signal_1717}), .Q ({data_out_s1[47], data_out_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_224 ( .clk (clk), .D ({signal_1723, signal_1721}), .Q ({data_out_s1[46], data_out_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_226 ( .clk (clk), .D ({signal_1727, signal_1725}), .Q ({data_out_s1[45], data_out_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_228 ( .clk (clk), .D ({signal_1731, signal_1729}), .Q ({data_out_s1[44], data_out_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_234 ( .clk (clk), .D ({signal_1735, signal_1733}), .Q ({data_out_s1[51], data_out_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_236 ( .clk (clk), .D ({signal_1739, signal_1737}), .Q ({data_out_s1[50], data_out_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_238 ( .clk (clk), .D ({signal_1743, signal_1741}), .Q ({data_out_s1[49], data_out_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_240 ( .clk (clk), .D ({signal_1747, signal_1745}), .Q ({data_out_s1[48], data_out_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_246 ( .clk (clk), .D ({signal_1751, signal_1749}), .Q ({data_out_s1[55], data_out_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_248 ( .clk (clk), .D ({signal_1755, signal_1753}), .Q ({data_out_s1[54], data_out_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_250 ( .clk (clk), .D ({signal_1759, signal_1757}), .Q ({data_out_s1[53], data_out_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_252 ( .clk (clk), .D ({signal_1763, signal_1761}), .Q ({data_out_s1[52], data_out_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_258 ( .clk (clk), .D ({signal_1767, signal_1765}), .Q ({data_out_s1[59], data_out_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_260 ( .clk (clk), .D ({signal_1771, signal_1769}), .Q ({data_out_s1[58], data_out_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_262 ( .clk (clk), .D ({signal_1775, signal_1773}), .Q ({data_out_s1[57], data_out_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_264 ( .clk (clk), .D ({signal_1779, signal_1777}), .Q ({data_out_s1[56], data_out_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_270 ( .clk (clk), .D ({signal_1783, signal_1781}), .Q ({data_out_s1[63], data_out_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_272 ( .clk (clk), .D ({signal_1787, signal_1785}), .Q ({data_out_s1[62], data_out_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_274 ( .clk (clk), .D ({signal_1791, signal_1789}), .Q ({data_out_s1[61], data_out_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_276 ( .clk (clk), .D ({signal_1795, signal_1793}), .Q ({data_out_s1[60], data_out_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_354 ( .clk (clk), .D ({signal_1799, signal_1797}), .Q ({signal_1064, signal_695}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_356 ( .clk (clk), .D ({signal_1803, signal_1801}), .Q ({signal_1291, signal_475}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_358 ( .clk (clk), .D ({signal_1807, signal_1805}), .Q ({signal_1289, signal_476}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_360 ( .clk (clk), .D ({signal_1811, signal_1809}), .Q ({signal_1287, signal_477}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_366 ( .clk (clk), .D ({signal_1815, signal_1813}), .Q ({signal_1076, signal_691}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_368 ( .clk (clk), .D ({signal_1819, signal_1817}), .Q ({signal_1073, signal_692}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_370 ( .clk (clk), .D ({signal_1823, signal_1821}), .Q ({signal_1070, signal_693}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_372 ( .clk (clk), .D ({signal_1827, signal_1825}), .Q ({signal_1067, signal_694}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_378 ( .clk (clk), .D ({signal_1831, signal_1829}), .Q ({signal_1088, signal_687}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_380 ( .clk (clk), .D ({signal_1835, signal_1833}), .Q ({signal_1085, signal_688}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_382 ( .clk (clk), .D ({signal_1839, signal_1837}), .Q ({signal_1082, signal_689}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_384 ( .clk (clk), .D ({signal_1843, signal_1841}), .Q ({signal_1079, signal_690}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_390 ( .clk (clk), .D ({signal_1847, signal_1845}), .Q ({signal_1100, signal_683}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_392 ( .clk (clk), .D ({signal_1851, signal_1849}), .Q ({signal_1097, signal_684}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_394 ( .clk (clk), .D ({signal_1855, signal_1853}), .Q ({signal_1094, signal_685}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_396 ( .clk (clk), .D ({signal_1859, signal_1857}), .Q ({signal_1091, signal_686}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_402 ( .clk (clk), .D ({signal_1863, signal_1861}), .Q ({signal_1274, signal_679}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_404 ( .clk (clk), .D ({signal_1867, signal_1865}), .Q ({signal_1062, signal_680}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_406 ( .clk (clk), .D ({signal_1871, signal_1869}), .Q ({signal_1106, signal_681}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_408 ( .clk (clk), .D ({signal_1875, signal_1873}), .Q ({signal_1103, signal_682}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_414 ( .clk (clk), .D ({signal_1879, signal_1877}), .Q ({signal_1109, signal_675}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_416 ( .clk (clk), .D ({signal_1883, signal_1881}), .Q ({signal_1056, signal_676}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_418 ( .clk (clk), .D ({signal_1887, signal_1885}), .Q ({signal_1058, signal_677}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_420 ( .clk (clk), .D ({signal_1891, signal_1889}), .Q ({signal_1060, signal_678}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_426 ( .clk (clk), .D ({signal_1895, signal_1893}), .Q ({signal_1121, signal_671}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_428 ( .clk (clk), .D ({signal_1899, signal_1897}), .Q ({signal_1118, signal_672}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_430 ( .clk (clk), .D ({signal_1903, signal_1901}), .Q ({signal_1115, signal_673}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_432 ( .clk (clk), .D ({signal_1907, signal_1905}), .Q ({signal_1112, signal_674}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_438 ( .clk (clk), .D ({signal_1911, signal_1909}), .Q ({signal_1133, signal_667}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_440 ( .clk (clk), .D ({signal_1915, signal_1913}), .Q ({signal_1130, signal_668}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_442 ( .clk (clk), .D ({signal_1919, signal_1917}), .Q ({signal_1127, signal_669}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_444 ( .clk (clk), .D ({signal_1923, signal_1921}), .Q ({signal_1124, signal_670}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_450 ( .clk (clk), .D ({signal_1927, signal_1925}), .Q ({signal_1145, signal_663}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_452 ( .clk (clk), .D ({signal_1931, signal_1929}), .Q ({signal_1142, signal_664}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_454 ( .clk (clk), .D ({signal_1935, signal_1933}), .Q ({signal_1139, signal_665}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_456 ( .clk (clk), .D ({signal_1939, signal_1937}), .Q ({signal_1136, signal_666}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_462 ( .clk (clk), .D ({signal_1943, signal_1941}), .Q ({signal_1157, signal_659}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_464 ( .clk (clk), .D ({signal_1947, signal_1945}), .Q ({signal_1154, signal_660}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_466 ( .clk (clk), .D ({signal_1951, signal_1949}), .Q ({signal_1151, signal_661}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_468 ( .clk (clk), .D ({signal_1955, signal_1953}), .Q ({signal_1148, signal_662}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_474 ( .clk (clk), .D ({signal_1959, signal_1957}), .Q ({signal_1169, signal_655}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_476 ( .clk (clk), .D ({signal_1963, signal_1961}), .Q ({signal_1166, signal_656}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_478 ( .clk (clk), .D ({signal_1967, signal_1965}), .Q ({signal_1163, signal_657}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_480 ( .clk (clk), .D ({signal_1971, signal_1969}), .Q ({signal_1160, signal_658}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_486 ( .clk (clk), .D ({signal_1975, signal_1973}), .Q ({signal_1181, signal_651}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_488 ( .clk (clk), .D ({signal_1979, signal_1977}), .Q ({signal_1178, signal_652}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_490 ( .clk (clk), .D ({signal_1983, signal_1981}), .Q ({signal_1175, signal_653}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_492 ( .clk (clk), .D ({signal_1987, signal_1985}), .Q ({signal_1172, signal_654}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_498 ( .clk (clk), .D ({signal_1991, signal_1989}), .Q ({signal_1193, signal_647}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_500 ( .clk (clk), .D ({signal_1995, signal_1993}), .Q ({signal_1190, signal_648}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_502 ( .clk (clk), .D ({signal_1999, signal_1997}), .Q ({signal_1187, signal_649}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_504 ( .clk (clk), .D ({signal_2003, signal_2001}), .Q ({signal_1184, signal_650}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_510 ( .clk (clk), .D ({signal_2007, signal_2005}), .Q ({signal_1205, signal_643}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_512 ( .clk (clk), .D ({signal_2011, signal_2009}), .Q ({signal_1202, signal_644}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_514 ( .clk (clk), .D ({signal_2015, signal_2013}), .Q ({signal_1199, signal_645}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_516 ( .clk (clk), .D ({signal_2019, signal_2017}), .Q ({signal_1196, signal_646}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_522 ( .clk (clk), .D ({signal_2023, signal_2021}), .Q ({signal_1217, signal_639}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_524 ( .clk (clk), .D ({signal_2027, signal_2025}), .Q ({signal_1214, signal_640}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_526 ( .clk (clk), .D ({signal_2031, signal_2029}), .Q ({signal_1211, signal_641}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_528 ( .clk (clk), .D ({signal_2035, signal_2033}), .Q ({signal_1208, signal_642}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_534 ( .clk (clk), .D ({signal_2039, signal_2037}), .Q ({signal_1229, signal_635}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_536 ( .clk (clk), .D ({signal_2043, signal_2041}), .Q ({signal_1226, signal_636}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_538 ( .clk (clk), .D ({signal_2047, signal_2045}), .Q ({signal_1223, signal_637}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_540 ( .clk (clk), .D ({signal_2051, signal_2049}), .Q ({signal_1220, signal_638}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_546 ( .clk (clk), .D ({signal_2055, signal_2053}), .Q ({signal_1241, signal_631}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_548 ( .clk (clk), .D ({signal_2059, signal_2057}), .Q ({signal_1238, signal_632}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_550 ( .clk (clk), .D ({signal_2063, signal_2061}), .Q ({signal_1235, signal_633}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_552 ( .clk (clk), .D ({signal_2067, signal_2065}), .Q ({signal_1232, signal_634}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_558 ( .clk (clk), .D ({signal_2071, signal_2069}), .Q ({signal_1253, signal_627}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_560 ( .clk (clk), .D ({signal_2075, signal_2073}), .Q ({signal_1250, signal_628}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_562 ( .clk (clk), .D ({signal_2079, signal_2077}), .Q ({signal_1247, signal_629}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_564 ( .clk (clk), .D ({signal_2083, signal_2081}), .Q ({signal_1244, signal_630}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_570 ( .clk (clk), .D ({signal_2087, signal_2085}), .Q ({signal_1265, signal_623}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_572 ( .clk (clk), .D ({signal_2091, signal_2089}), .Q ({signal_1262, signal_624}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_574 ( .clk (clk), .D ({signal_2095, signal_2093}), .Q ({signal_1259, signal_625}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_576 ( .clk (clk), .D ({signal_2099, signal_2097}), .Q ({signal_1256, signal_626}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_582 ( .clk (clk), .D ({signal_1453, signal_852}), .Q ({signal_865, signal_471}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_584 ( .clk (clk), .D ({signal_1448, signal_853}), .Q ({signal_862, signal_472}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_586 ( .clk (clk), .D ({signal_1447, signal_854}), .Q ({signal_859, signal_473}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_588 ( .clk (clk), .D ({signal_1446, signal_855}), .Q ({signal_856, signal_474}) ) ;
endmodule
