/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module LED_HPC2_BDDsylvan_Pipeline_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [597:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_356 ;
    wire signal_375 ;
    wire signal_394 ;
    wire signal_413 ;
    wire signal_432 ;
    wire signal_451 ;
    wire signal_470 ;
    wire signal_489 ;
    wire signal_508 ;
    wire signal_527 ;
    wire signal_546 ;
    wire signal_565 ;
    wire signal_584 ;
    wire signal_603 ;
    wire signal_622 ;
    wire signal_641 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1856 ;
    wire signal_1859 ;
    wire signal_1862 ;
    wire signal_1865 ;
    wire signal_1868 ;
    wire signal_1871 ;
    wire signal_1874 ;
    wire signal_1877 ;
    wire signal_1880 ;
    wire signal_1883 ;
    wire signal_1886 ;
    wire signal_1889 ;
    wire signal_1892 ;
    wire signal_1894 ;
    wire signal_1896 ;
    wire signal_1898 ;
    wire signal_1900 ;
    wire signal_1902 ;
    wire signal_1904 ;
    wire signal_1906 ;
    wire signal_1908 ;
    wire signal_1910 ;
    wire signal_1912 ;
    wire signal_1914 ;
    wire signal_1916 ;
    wire signal_1918 ;
    wire signal_1921 ;
    wire signal_1924 ;
    wire signal_1927 ;
    wire signal_1930 ;
    wire signal_1933 ;
    wire signal_1936 ;
    wire signal_1939 ;
    wire signal_1942 ;
    wire signal_1945 ;
    wire signal_1948 ;
    wire signal_1951 ;
    wire signal_1954 ;
    wire signal_1957 ;
    wire signal_1960 ;
    wire signal_1963 ;
    wire signal_1966 ;
    wire signal_1969 ;
    wire signal_1972 ;
    wire signal_1975 ;
    wire signal_1978 ;
    wire signal_1981 ;
    wire signal_1984 ;
    wire signal_1987 ;
    wire signal_1990 ;
    wire signal_1993 ;
    wire signal_1996 ;
    wire signal_1999 ;
    wire signal_2002 ;
    wire signal_2005 ;
    wire signal_2008 ;
    wire signal_2011 ;
    wire signal_2014 ;
    wire signal_2017 ;
    wire signal_2020 ;
    wire signal_2023 ;
    wire signal_2026 ;
    wire signal_2029 ;
    wire signal_2032 ;
    wire signal_2035 ;
    wire signal_2038 ;
    wire signal_2041 ;
    wire signal_2044 ;
    wire signal_2047 ;
    wire signal_2050 ;
    wire signal_2053 ;
    wire signal_2056 ;
    wire signal_2059 ;
    wire signal_2062 ;
    wire signal_2065 ;
    wire signal_2068 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2080 ;
    wire signal_2082 ;
    wire signal_2084 ;
    wire signal_2086 ;
    wire signal_2088 ;
    wire signal_2090 ;
    wire signal_2092 ;
    wire signal_2094 ;
    wire signal_2096 ;
    wire signal_2098 ;
    wire signal_2100 ;
    wire signal_2102 ;
    wire signal_2104 ;
    wire signal_2106 ;
    wire signal_2108 ;
    wire signal_2110 ;
    wire signal_2112 ;
    wire signal_2114 ;
    wire signal_2116 ;
    wire signal_2118 ;
    wire signal_2120 ;
    wire signal_2122 ;
    wire signal_2124 ;
    wire signal_2126 ;
    wire signal_2128 ;
    wire signal_2130 ;
    wire signal_2132 ;
    wire signal_2134 ;
    wire signal_2136 ;
    wire signal_2138 ;
    wire signal_2140 ;
    wire signal_2142 ;
    wire signal_2144 ;
    wire signal_2146 ;
    wire signal_2148 ;
    wire signal_2150 ;
    wire signal_2152 ;
    wire signal_2154 ;
    wire signal_2156 ;
    wire signal_2158 ;
    wire signal_2160 ;
    wire signal_2162 ;
    wire signal_2164 ;
    wire signal_2166 ;
    wire signal_2168 ;
    wire signal_2170 ;
    wire signal_2172 ;
    wire signal_2174 ;
    wire signal_2176 ;
    wire signal_2178 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2992 ;
    wire signal_2994 ;
    wire signal_2996 ;
    wire signal_2998 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3026 ;
    wire signal_3028 ;
    wire signal_3030 ;
    wire signal_3032 ;
    wire signal_3034 ;
    wire signal_3036 ;
    wire signal_3038 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3065 ;
    wire signal_3067 ;
    wire signal_3069 ;
    wire signal_3071 ;
    wire signal_3073 ;
    wire signal_3075 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3112 ;
    wire signal_3114 ;
    wire signal_3116 ;
    wire signal_3118 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3143 ;
    wire signal_3145 ;
    wire signal_3147 ;
    wire signal_3149 ;
    wire signal_3151 ;
    wire signal_3153 ;
    wire signal_3155 ;
    wire signal_3157 ;
    wire signal_3159 ;
    wire signal_3161 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3189 ;
    wire signal_3191 ;
    wire signal_3193 ;
    wire signal_3195 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3215 ;
    wire signal_3217 ;
    wire signal_3219 ;
    wire signal_3221 ;
    wire signal_3223 ;
    wire signal_3225 ;
    wire signal_3227 ;
    wire signal_3229 ;
    wire signal_3231 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3243 ;
    wire signal_3245 ;
    wire signal_3247 ;
    wire signal_3249 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3265 ;
    wire signal_3267 ;
    wire signal_3269 ;
    wire signal_3271 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7759 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7762 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7765 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7768 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7771 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7774 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7777 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7780 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7783 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7786 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7789 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7792 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7795 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7798 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7801 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7804 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7807 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7810 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7813 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7816 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7819 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7822 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7825 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7828 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7831 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7834 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7837 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7840 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;
    wire signal_7973 ;
    wire signal_7974 ;
    wire signal_7975 ;
    wire signal_7976 ;
    wire signal_7977 ;
    wire signal_7978 ;
    wire signal_7979 ;
    wire signal_7980 ;
    wire signal_7981 ;
    wire signal_7982 ;
    wire signal_7983 ;
    wire signal_7984 ;
    wire signal_7985 ;
    wire signal_7986 ;
    wire signal_7987 ;
    wire signal_7988 ;
    wire signal_7989 ;
    wire signal_7990 ;
    wire signal_7991 ;
    wire signal_7992 ;
    wire signal_7993 ;
    wire signal_7994 ;
    wire signal_7995 ;
    wire signal_7996 ;
    wire signal_7997 ;
    wire signal_7998 ;
    wire signal_7999 ;
    wire signal_8000 ;
    wire signal_8001 ;
    wire signal_8002 ;
    wire signal_8003 ;
    wire signal_8004 ;
    wire signal_8005 ;
    wire signal_8006 ;
    wire signal_8007 ;
    wire signal_8008 ;
    wire signal_8009 ;
    wire signal_8010 ;
    wire signal_8011 ;
    wire signal_8012 ;
    wire signal_8013 ;
    wire signal_8014 ;
    wire signal_8015 ;
    wire signal_8016 ;
    wire signal_8017 ;
    wire signal_8018 ;
    wire signal_8019 ;
    wire signal_8020 ;
    wire signal_8021 ;
    wire signal_8022 ;
    wire signal_8023 ;
    wire signal_8024 ;
    wire signal_8025 ;
    wire signal_8026 ;
    wire signal_8027 ;
    wire signal_8028 ;
    wire signal_8029 ;
    wire signal_8030 ;
    wire signal_8031 ;
    wire signal_8032 ;
    wire signal_8033 ;
    wire signal_8034 ;
    wire signal_8035 ;
    wire signal_8036 ;
    wire signal_8037 ;
    wire signal_8038 ;
    wire signal_8039 ;
    wire signal_8040 ;
    wire signal_8041 ;
    wire signal_8042 ;
    wire signal_8043 ;
    wire signal_8044 ;
    wire signal_8045 ;
    wire signal_8046 ;
    wire signal_8047 ;
    wire signal_8048 ;
    wire signal_8049 ;
    wire signal_8050 ;
    wire signal_8051 ;
    wire signal_8052 ;
    wire signal_8053 ;
    wire signal_8054 ;
    wire signal_8055 ;
    wire signal_8056 ;
    wire signal_8057 ;
    wire signal_8058 ;
    wire signal_8059 ;
    wire signal_8060 ;
    wire signal_8061 ;
    wire signal_8062 ;
    wire signal_8063 ;
    wire signal_8064 ;
    wire signal_8065 ;
    wire signal_8066 ;
    wire signal_8067 ;
    wire signal_8068 ;
    wire signal_8069 ;
    wire signal_8070 ;
    wire signal_8071 ;
    wire signal_8072 ;
    wire signal_8073 ;
    wire signal_8074 ;
    wire signal_8075 ;
    wire signal_8076 ;
    wire signal_8077 ;
    wire signal_8078 ;
    wire signal_8079 ;
    wire signal_8080 ;
    wire signal_8081 ;
    wire signal_8082 ;
    wire signal_8083 ;
    wire signal_8084 ;
    wire signal_8085 ;
    wire signal_8086 ;
    wire signal_8087 ;
    wire signal_8088 ;
    wire signal_8089 ;
    wire signal_8090 ;
    wire signal_8091 ;
    wire signal_8092 ;
    wire signal_8093 ;
    wire signal_8094 ;
    wire signal_8095 ;
    wire signal_8096 ;
    wire signal_8097 ;
    wire signal_8098 ;
    wire signal_8099 ;
    wire signal_8100 ;
    wire signal_8101 ;
    wire signal_8102 ;
    wire signal_8103 ;
    wire signal_8104 ;
    wire signal_8105 ;
    wire signal_8106 ;
    wire signal_8107 ;
    wire signal_8108 ;
    wire signal_8109 ;
    wire signal_8110 ;
    wire signal_8111 ;
    wire signal_8112 ;
    wire signal_8113 ;
    wire signal_8114 ;
    wire signal_8115 ;
    wire signal_8116 ;
    wire signal_8117 ;
    wire signal_8118 ;
    wire signal_8119 ;
    wire signal_8120 ;
    wire signal_8121 ;
    wire signal_8122 ;
    wire signal_8123 ;
    wire signal_8124 ;
    wire signal_8125 ;
    wire signal_8126 ;
    wire signal_8127 ;
    wire signal_8128 ;
    wire signal_8129 ;
    wire signal_8130 ;
    wire signal_8131 ;
    wire signal_8132 ;
    wire signal_8133 ;
    wire signal_8134 ;
    wire signal_8135 ;
    wire signal_8136 ;
    wire signal_8137 ;
    wire signal_8138 ;
    wire signal_8139 ;
    wire signal_8140 ;
    wire signal_8141 ;
    wire signal_8142 ;
    wire signal_8143 ;
    wire signal_8144 ;
    wire signal_8145 ;
    wire signal_8146 ;
    wire signal_8147 ;
    wire signal_8148 ;
    wire signal_8149 ;
    wire signal_8150 ;
    wire signal_8151 ;
    wire signal_8152 ;
    wire signal_8153 ;
    wire signal_8154 ;
    wire signal_8155 ;
    wire signal_8156 ;
    wire signal_8157 ;
    wire signal_8158 ;
    wire signal_8159 ;
    wire signal_8160 ;
    wire signal_8161 ;
    wire signal_8162 ;
    wire signal_8163 ;
    wire signal_8164 ;
    wire signal_8165 ;
    wire signal_8166 ;
    wire signal_8167 ;
    wire signal_8168 ;
    wire signal_8169 ;
    wire signal_8170 ;
    wire signal_8171 ;
    wire signal_8172 ;
    wire signal_8173 ;
    wire signal_8174 ;
    wire signal_8175 ;
    wire signal_8176 ;
    wire signal_8177 ;
    wire signal_8178 ;
    wire signal_8179 ;
    wire signal_8180 ;
    wire signal_8181 ;
    wire signal_8182 ;
    wire signal_8183 ;
    wire signal_8184 ;
    wire signal_8185 ;
    wire signal_8186 ;
    wire signal_8187 ;
    wire signal_8188 ;
    wire signal_8189 ;
    wire signal_8190 ;
    wire signal_8191 ;
    wire signal_8192 ;
    wire signal_8193 ;
    wire signal_8194 ;
    wire signal_8195 ;
    wire signal_8196 ;
    wire signal_8197 ;
    wire signal_8198 ;
    wire signal_8199 ;
    wire signal_8200 ;
    wire signal_8201 ;
    wire signal_8202 ;
    wire signal_8203 ;
    wire signal_8204 ;
    wire signal_8205 ;
    wire signal_8206 ;
    wire signal_8207 ;
    wire signal_8208 ;
    wire signal_8209 ;
    wire signal_8210 ;
    wire signal_8211 ;
    wire signal_8212 ;
    wire signal_8213 ;
    wire signal_8214 ;
    wire signal_8215 ;
    wire signal_8216 ;
    wire signal_8217 ;
    wire signal_8218 ;
    wire signal_8219 ;
    wire signal_8220 ;
    wire signal_8221 ;
    wire signal_8222 ;
    wire signal_8223 ;
    wire signal_8224 ;
    wire signal_8225 ;
    wire signal_8226 ;
    wire signal_8227 ;
    wire signal_8228 ;
    wire signal_8229 ;
    wire signal_8230 ;
    wire signal_8231 ;
    wire signal_8232 ;
    wire signal_8233 ;
    wire signal_8234 ;
    wire signal_8235 ;
    wire signal_8236 ;
    wire signal_8237 ;
    wire signal_8238 ;
    wire signal_8239 ;
    wire signal_8240 ;
    wire signal_8241 ;
    wire signal_8242 ;
    wire signal_8243 ;
    wire signal_8244 ;
    wire signal_8245 ;
    wire signal_8246 ;
    wire signal_8247 ;
    wire signal_8248 ;
    wire signal_8249 ;
    wire signal_8250 ;
    wire signal_8251 ;
    wire signal_8252 ;
    wire signal_8253 ;
    wire signal_8254 ;
    wire signal_8255 ;
    wire signal_8256 ;
    wire signal_8257 ;
    wire signal_8258 ;
    wire signal_8259 ;
    wire signal_8260 ;
    wire signal_8261 ;
    wire signal_8262 ;
    wire signal_8263 ;
    wire signal_8264 ;
    wire signal_8265 ;
    wire signal_8266 ;
    wire signal_8267 ;
    wire signal_8268 ;
    wire signal_8269 ;
    wire signal_8270 ;
    wire signal_8271 ;
    wire signal_8272 ;
    wire signal_8273 ;
    wire signal_8274 ;
    wire signal_8275 ;
    wire signal_8276 ;
    wire signal_8277 ;
    wire signal_8278 ;
    wire signal_8279 ;
    wire signal_8280 ;
    wire signal_8281 ;
    wire signal_8282 ;
    wire signal_8283 ;
    wire signal_8284 ;
    wire signal_8285 ;
    wire signal_8286 ;
    wire signal_8287 ;
    wire signal_8288 ;
    wire signal_8289 ;
    wire signal_8290 ;
    wire signal_8291 ;
    wire signal_8292 ;
    wire signal_8293 ;
    wire signal_8294 ;
    wire signal_8295 ;
    wire signal_8296 ;
    wire signal_8297 ;
    wire signal_8298 ;
    wire signal_8299 ;
    wire signal_8300 ;
    wire signal_8301 ;
    wire signal_8302 ;
    wire signal_8303 ;
    wire signal_8304 ;
    wire signal_8305 ;
    wire signal_8306 ;
    wire signal_8307 ;
    wire signal_8308 ;
    wire signal_8309 ;
    wire signal_8310 ;
    wire signal_8311 ;
    wire signal_8312 ;
    wire signal_8313 ;
    wire signal_8314 ;
    wire signal_8315 ;
    wire signal_8316 ;
    wire signal_8317 ;
    wire signal_8318 ;
    wire signal_8319 ;
    wire signal_8320 ;
    wire signal_8321 ;
    wire signal_8322 ;
    wire signal_8323 ;
    wire signal_8324 ;
    wire signal_8325 ;
    wire signal_8326 ;
    wire signal_8327 ;
    wire signal_8328 ;
    wire signal_8329 ;
    wire signal_8330 ;
    wire signal_8331 ;
    wire signal_8332 ;
    wire signal_8333 ;
    wire signal_8334 ;
    wire signal_8335 ;
    wire signal_8336 ;
    wire signal_8337 ;
    wire signal_8338 ;
    wire signal_8339 ;
    wire signal_8340 ;
    wire signal_8341 ;
    wire signal_8342 ;
    wire signal_8343 ;
    wire signal_8344 ;
    wire signal_8345 ;
    wire signal_8346 ;
    wire signal_8347 ;
    wire signal_8348 ;
    wire signal_8349 ;
    wire signal_8350 ;
    wire signal_8351 ;
    wire signal_8352 ;
    wire signal_8353 ;
    wire signal_8354 ;
    wire signal_8355 ;
    wire signal_8356 ;
    wire signal_8357 ;
    wire signal_8358 ;
    wire signal_8359 ;
    wire signal_8360 ;
    wire signal_8361 ;
    wire signal_8362 ;
    wire signal_8363 ;
    wire signal_8364 ;
    wire signal_8365 ;
    wire signal_8366 ;
    wire signal_8367 ;
    wire signal_8368 ;
    wire signal_8369 ;
    wire signal_8370 ;
    wire signal_8371 ;
    wire signal_8372 ;
    wire signal_8373 ;
    wire signal_8374 ;
    wire signal_8375 ;
    wire signal_8376 ;
    wire signal_8377 ;
    wire signal_8378 ;
    wire signal_8379 ;
    wire signal_8380 ;
    wire signal_8381 ;
    wire signal_8382 ;
    wire signal_8383 ;
    wire signal_8384 ;
    wire signal_8385 ;
    wire signal_8386 ;
    wire signal_8387 ;
    wire signal_8388 ;
    wire signal_8389 ;
    wire signal_8390 ;
    wire signal_8391 ;
    wire signal_8392 ;
    wire signal_8393 ;
    wire signal_8394 ;
    wire signal_8395 ;
    wire signal_8396 ;
    wire signal_8397 ;
    wire signal_8398 ;
    wire signal_8399 ;
    wire signal_8400 ;
    wire signal_8401 ;
    wire signal_8402 ;
    wire signal_8403 ;
    wire signal_8404 ;
    wire signal_8405 ;
    wire signal_8406 ;
    wire signal_8407 ;
    wire signal_8408 ;
    wire signal_8409 ;
    wire signal_8410 ;
    wire signal_8411 ;
    wire signal_8412 ;
    wire signal_8413 ;
    wire signal_8414 ;
    wire signal_8415 ;
    wire signal_8416 ;
    wire signal_8417 ;
    wire signal_8418 ;
    wire signal_8419 ;
    wire signal_8420 ;
    wire signal_8421 ;
    wire signal_8422 ;
    wire signal_8423 ;
    wire signal_8424 ;
    wire signal_8425 ;
    wire signal_8426 ;
    wire signal_8427 ;
    wire signal_8428 ;
    wire signal_8429 ;
    wire signal_8430 ;
    wire signal_8431 ;
    wire signal_8432 ;
    wire signal_8433 ;
    wire signal_8434 ;
    wire signal_8435 ;
    wire signal_8436 ;
    wire signal_8437 ;
    wire signal_8438 ;
    wire signal_8439 ;
    wire signal_8440 ;
    wire signal_8441 ;
    wire signal_8442 ;
    wire signal_8443 ;
    wire signal_8444 ;
    wire signal_8445 ;
    wire signal_8446 ;
    wire signal_8447 ;
    wire signal_8448 ;
    wire signal_8449 ;
    wire signal_8450 ;
    wire signal_8451 ;
    wire signal_8452 ;
    wire signal_8453 ;
    wire signal_8454 ;
    wire signal_8455 ;
    wire signal_8456 ;
    wire signal_8457 ;
    wire signal_8458 ;
    wire signal_8459 ;
    wire signal_8460 ;
    wire signal_8461 ;
    wire signal_8462 ;
    wire signal_8463 ;
    wire signal_8464 ;
    wire signal_8465 ;
    wire signal_8466 ;
    wire signal_8467 ;
    wire signal_8468 ;
    wire signal_8469 ;
    wire signal_8470 ;
    wire signal_8471 ;
    wire signal_8472 ;
    wire signal_8473 ;
    wire signal_8474 ;
    wire signal_8475 ;
    wire signal_8476 ;
    wire signal_8477 ;
    wire signal_8478 ;
    wire signal_8479 ;
    wire signal_8480 ;
    wire signal_8481 ;
    wire signal_8482 ;
    wire signal_8483 ;
    wire signal_8484 ;
    wire signal_8485 ;
    wire signal_8486 ;
    wire signal_8487 ;
    wire signal_8488 ;
    wire signal_8489 ;
    wire signal_8490 ;
    wire signal_8491 ;
    wire signal_8492 ;
    wire signal_8493 ;
    wire signal_8494 ;
    wire signal_8495 ;
    wire signal_8496 ;
    wire signal_8497 ;
    wire signal_8498 ;
    wire signal_8499 ;
    wire signal_8500 ;
    wire signal_8501 ;
    wire signal_8502 ;
    wire signal_8503 ;
    wire signal_8504 ;
    wire signal_8505 ;
    wire signal_8506 ;
    wire signal_8507 ;
    wire signal_8508 ;
    wire signal_8509 ;
    wire signal_8510 ;
    wire signal_8511 ;
    wire signal_8512 ;
    wire signal_8513 ;
    wire signal_8514 ;
    wire signal_8515 ;
    wire signal_8516 ;
    wire signal_8517 ;
    wire signal_8518 ;
    wire signal_8519 ;
    wire signal_8520 ;
    wire signal_8521 ;
    wire signal_8522 ;
    wire signal_8523 ;
    wire signal_8524 ;
    wire signal_8525 ;
    wire signal_8526 ;
    wire signal_8527 ;
    wire signal_8528 ;
    wire signal_8529 ;
    wire signal_8530 ;
    wire signal_8531 ;
    wire signal_8532 ;
    wire signal_8533 ;
    wire signal_8534 ;
    wire signal_8535 ;
    wire signal_8536 ;
    wire signal_8537 ;
    wire signal_8538 ;
    wire signal_8539 ;
    wire signal_8540 ;
    wire signal_8541 ;
    wire signal_8542 ;
    wire signal_8543 ;
    wire signal_8544 ;
    wire signal_8545 ;
    wire signal_8546 ;
    wire signal_8547 ;
    wire signal_8548 ;
    wire signal_8549 ;
    wire signal_8550 ;
    wire signal_8551 ;
    wire signal_8552 ;
    wire signal_8553 ;
    wire signal_8554 ;
    wire signal_8555 ;
    wire signal_8556 ;
    wire signal_8557 ;
    wire signal_8558 ;
    wire signal_8559 ;
    wire signal_8560 ;
    wire signal_8561 ;
    wire signal_8562 ;
    wire signal_8563 ;
    wire signal_8564 ;
    wire signal_8565 ;
    wire signal_8566 ;
    wire signal_8567 ;
    wire signal_8568 ;
    wire signal_8569 ;
    wire signal_8570 ;
    wire signal_8571 ;
    wire signal_8572 ;
    wire signal_8573 ;
    wire signal_8574 ;
    wire signal_8575 ;
    wire signal_8576 ;
    wire signal_8577 ;
    wire signal_8578 ;
    wire signal_8579 ;
    wire signal_8580 ;
    wire signal_8581 ;
    wire signal_8582 ;
    wire signal_8583 ;
    wire signal_8584 ;
    wire signal_8585 ;
    wire signal_8586 ;
    wire signal_8587 ;
    wire signal_8588 ;
    wire signal_8589 ;
    wire signal_8590 ;
    wire signal_8591 ;
    wire signal_8592 ;
    wire signal_8593 ;
    wire signal_8594 ;
    wire signal_8595 ;
    wire signal_8596 ;
    wire signal_8597 ;
    wire signal_8598 ;
    wire signal_8599 ;
    wire signal_8600 ;
    wire signal_8601 ;
    wire signal_8602 ;
    wire signal_8603 ;
    wire signal_8604 ;
    wire signal_8605 ;
    wire signal_8606 ;
    wire signal_8607 ;
    wire signal_8608 ;
    wire signal_8609 ;
    wire signal_8610 ;
    wire signal_8611 ;
    wire signal_8612 ;
    wire signal_8613 ;
    wire signal_8614 ;
    wire signal_8615 ;
    wire signal_8616 ;
    wire signal_8617 ;
    wire signal_8618 ;
    wire signal_8619 ;
    wire signal_8620 ;
    wire signal_8621 ;
    wire signal_8622 ;
    wire signal_8623 ;
    wire signal_8624 ;
    wire signal_8625 ;
    wire signal_8626 ;
    wire signal_8627 ;
    wire signal_8628 ;
    wire signal_8629 ;
    wire signal_8630 ;
    wire signal_8631 ;
    wire signal_8632 ;
    wire signal_8633 ;
    wire signal_8634 ;
    wire signal_8635 ;
    wire signal_8636 ;
    wire signal_8637 ;
    wire signal_8638 ;
    wire signal_8639 ;
    wire signal_8640 ;
    wire signal_8641 ;
    wire signal_8642 ;
    wire signal_8643 ;
    wire signal_8644 ;
    wire signal_8645 ;
    wire signal_8646 ;
    wire signal_8647 ;
    wire signal_8648 ;
    wire signal_8649 ;
    wire signal_8650 ;
    wire signal_8651 ;
    wire signal_8652 ;
    wire signal_8653 ;
    wire signal_8654 ;
    wire signal_8655 ;
    wire signal_8656 ;
    wire signal_8657 ;
    wire signal_8658 ;
    wire signal_8659 ;
    wire signal_8660 ;
    wire signal_8661 ;
    wire signal_8662 ;
    wire signal_8663 ;
    wire signal_8664 ;
    wire signal_8665 ;
    wire signal_8666 ;
    wire signal_8667 ;
    wire signal_8668 ;
    wire signal_8669 ;
    wire signal_8670 ;
    wire signal_8671 ;
    wire signal_8672 ;
    wire signal_8673 ;
    wire signal_8674 ;
    wire signal_8675 ;
    wire signal_8676 ;
    wire signal_8677 ;
    wire signal_8678 ;
    wire signal_8679 ;
    wire signal_8680 ;
    wire signal_8681 ;
    wire signal_8682 ;
    wire signal_8683 ;
    wire signal_8684 ;
    wire signal_8685 ;
    wire signal_8686 ;
    wire signal_8687 ;
    wire signal_8688 ;
    wire signal_8689 ;
    wire signal_8690 ;
    wire signal_8691 ;
    wire signal_8692 ;
    wire signal_8693 ;
    wire signal_8694 ;
    wire signal_8695 ;
    wire signal_8696 ;
    wire signal_8697 ;
    wire signal_8698 ;
    wire signal_8699 ;
    wire signal_8700 ;
    wire signal_8701 ;
    wire signal_8702 ;
    wire signal_8703 ;
    wire signal_8704 ;
    wire signal_8705 ;
    wire signal_8706 ;
    wire signal_8707 ;
    wire signal_8708 ;
    wire signal_8709 ;
    wire signal_8710 ;
    wire signal_8711 ;
    wire signal_8712 ;
    wire signal_8713 ;
    wire signal_8714 ;
    wire signal_8715 ;
    wire signal_8716 ;
    wire signal_8717 ;
    wire signal_8718 ;
    wire signal_8719 ;
    wire signal_8720 ;
    wire signal_8721 ;
    wire signal_8722 ;
    wire signal_8723 ;
    wire signal_8724 ;
    wire signal_8725 ;
    wire signal_8726 ;
    wire signal_8727 ;
    wire signal_8728 ;
    wire signal_8729 ;
    wire signal_8730 ;
    wire signal_8731 ;
    wire signal_8732 ;
    wire signal_8733 ;
    wire signal_8734 ;
    wire signal_8735 ;
    wire signal_8736 ;
    wire signal_8737 ;
    wire signal_8738 ;
    wire signal_8739 ;
    wire signal_8740 ;
    wire signal_8741 ;
    wire signal_8742 ;
    wire signal_8743 ;
    wire signal_8744 ;
    wire signal_8745 ;
    wire signal_8746 ;
    wire signal_8747 ;
    wire signal_8748 ;
    wire signal_8749 ;
    wire signal_8750 ;
    wire signal_8751 ;
    wire signal_8752 ;
    wire signal_8753 ;
    wire signal_8754 ;
    wire signal_8755 ;
    wire signal_8756 ;
    wire signal_8757 ;
    wire signal_8758 ;
    wire signal_8759 ;
    wire signal_8760 ;
    wire signal_8761 ;
    wire signal_8762 ;
    wire signal_8763 ;
    wire signal_8764 ;
    wire signal_8765 ;
    wire signal_8766 ;
    wire signal_8767 ;
    wire signal_8768 ;
    wire signal_8769 ;
    wire signal_8770 ;
    wire signal_8771 ;
    wire signal_8772 ;
    wire signal_8773 ;
    wire signal_8774 ;
    wire signal_8775 ;
    wire signal_8776 ;
    wire signal_8777 ;
    wire signal_8778 ;
    wire signal_8779 ;
    wire signal_8780 ;
    wire signal_8781 ;
    wire signal_8782 ;
    wire signal_8783 ;
    wire signal_8784 ;
    wire signal_8785 ;
    wire signal_8786 ;
    wire signal_8787 ;
    wire signal_8788 ;
    wire signal_8789 ;
    wire signal_8790 ;
    wire signal_8791 ;
    wire signal_8792 ;
    wire signal_8793 ;
    wire signal_8794 ;
    wire signal_8795 ;
    wire signal_8796 ;
    wire signal_8797 ;
    wire signal_8798 ;
    wire signal_8799 ;
    wire signal_8800 ;
    wire signal_8801 ;
    wire signal_8802 ;
    wire signal_8803 ;
    wire signal_8804 ;
    wire signal_8805 ;
    wire signal_8806 ;
    wire signal_8807 ;
    wire signal_8808 ;
    wire signal_8809 ;
    wire signal_8810 ;
    wire signal_8811 ;
    wire signal_8812 ;
    wire signal_8813 ;
    wire signal_8814 ;
    wire signal_8815 ;
    wire signal_8816 ;
    wire signal_8817 ;
    wire signal_8818 ;
    wire signal_8819 ;
    wire signal_8820 ;
    wire signal_8821 ;
    wire signal_8822 ;
    wire signal_8823 ;
    wire signal_8824 ;
    wire signal_8825 ;
    wire signal_8826 ;
    wire signal_8827 ;
    wire signal_8828 ;
    wire signal_8829 ;
    wire signal_8830 ;
    wire signal_8831 ;
    wire signal_8832 ;
    wire signal_8833 ;
    wire signal_8834 ;
    wire signal_8835 ;
    wire signal_8836 ;
    wire signal_8837 ;
    wire signal_8838 ;
    wire signal_8839 ;
    wire signal_8840 ;
    wire signal_8841 ;
    wire signal_8842 ;
    wire signal_8843 ;
    wire signal_8844 ;
    wire signal_8845 ;
    wire signal_8846 ;
    wire signal_8847 ;
    wire signal_8848 ;
    wire signal_8849 ;
    wire signal_8850 ;
    wire signal_8851 ;
    wire signal_8852 ;
    wire signal_8853 ;
    wire signal_8854 ;
    wire signal_8855 ;
    wire signal_8856 ;
    wire signal_8857 ;
    wire signal_8858 ;
    wire signal_8859 ;
    wire signal_8860 ;
    wire signal_8861 ;
    wire signal_8862 ;
    wire signal_8863 ;
    wire signal_8864 ;
    wire signal_8865 ;
    wire signal_8866 ;
    wire signal_8867 ;
    wire signal_8868 ;
    wire signal_8869 ;
    wire signal_8870 ;
    wire signal_8871 ;
    wire signal_8872 ;
    wire signal_8873 ;
    wire signal_8874 ;
    wire signal_8875 ;
    wire signal_8876 ;
    wire signal_8877 ;
    wire signal_8878 ;
    wire signal_8879 ;
    wire signal_8880 ;
    wire signal_8881 ;
    wire signal_8882 ;
    wire signal_8883 ;
    wire signal_8884 ;
    wire signal_8885 ;
    wire signal_8886 ;
    wire signal_8887 ;
    wire signal_8888 ;
    wire signal_8889 ;
    wire signal_8890 ;
    wire signal_8891 ;
    wire signal_8892 ;
    wire signal_8893 ;
    wire signal_8894 ;
    wire signal_8895 ;
    wire signal_8896 ;
    wire signal_8897 ;
    wire signal_8898 ;
    wire signal_8899 ;
    wire signal_8900 ;
    wire signal_8901 ;
    wire signal_8902 ;
    wire signal_8903 ;
    wire signal_8904 ;
    wire signal_8905 ;
    wire signal_8906 ;
    wire signal_8907 ;
    wire signal_8908 ;
    wire signal_8909 ;
    wire signal_8910 ;
    wire signal_8911 ;
    wire signal_8912 ;
    wire signal_8913 ;
    wire signal_8914 ;
    wire signal_8915 ;
    wire signal_8916 ;
    wire signal_8917 ;
    wire signal_8918 ;
    wire signal_8919 ;
    wire signal_8920 ;
    wire signal_8921 ;
    wire signal_8922 ;
    wire signal_8923 ;
    wire signal_8924 ;
    wire signal_8925 ;
    wire signal_8926 ;
    wire signal_8927 ;
    wire signal_8928 ;
    wire signal_8929 ;
    wire signal_8930 ;
    wire signal_8931 ;
    wire signal_8932 ;
    wire signal_8933 ;
    wire signal_8934 ;
    wire signal_8935 ;
    wire signal_8936 ;
    wire signal_8937 ;
    wire signal_8938 ;
    wire signal_8939 ;
    wire signal_8940 ;
    wire signal_8941 ;
    wire signal_8942 ;
    wire signal_8943 ;
    wire signal_8944 ;
    wire signal_8945 ;
    wire signal_8946 ;
    wire signal_8947 ;
    wire signal_8948 ;
    wire signal_8949 ;
    wire signal_8950 ;
    wire signal_8951 ;
    wire signal_8952 ;
    wire signal_8953 ;
    wire signal_8954 ;
    wire signal_8955 ;
    wire signal_8956 ;
    wire signal_8957 ;
    wire signal_8958 ;
    wire signal_8959 ;
    wire signal_8960 ;
    wire signal_8961 ;
    wire signal_8962 ;
    wire signal_8963 ;
    wire signal_8964 ;
    wire signal_8965 ;
    wire signal_8966 ;
    wire signal_8967 ;
    wire signal_8968 ;
    wire signal_8969 ;
    wire signal_8970 ;
    wire signal_8971 ;
    wire signal_8972 ;
    wire signal_8973 ;
    wire signal_8974 ;
    wire signal_8975 ;
    wire signal_8976 ;
    wire signal_8977 ;
    wire signal_8978 ;
    wire signal_8979 ;
    wire signal_8980 ;
    wire signal_8981 ;
    wire signal_8982 ;
    wire signal_8983 ;
    wire signal_8984 ;
    wire signal_8985 ;
    wire signal_8986 ;
    wire signal_8987 ;
    wire signal_8988 ;
    wire signal_8989 ;
    wire signal_8990 ;
    wire signal_8991 ;
    wire signal_8992 ;
    wire signal_8993 ;
    wire signal_8994 ;
    wire signal_8995 ;
    wire signal_8996 ;
    wire signal_8997 ;
    wire signal_8998 ;
    wire signal_8999 ;
    wire signal_9000 ;
    wire signal_9001 ;
    wire signal_9002 ;
    wire signal_9003 ;
    wire signal_9004 ;
    wire signal_9005 ;
    wire signal_9006 ;
    wire signal_9007 ;
    wire signal_9008 ;
    wire signal_9009 ;
    wire signal_9010 ;
    wire signal_9011 ;
    wire signal_9012 ;
    wire signal_9013 ;
    wire signal_9014 ;
    wire signal_9015 ;
    wire signal_9016 ;
    wire signal_9017 ;
    wire signal_9018 ;
    wire signal_9019 ;
    wire signal_9020 ;
    wire signal_9021 ;
    wire signal_9022 ;
    wire signal_9023 ;
    wire signal_9024 ;
    wire signal_9025 ;
    wire signal_9026 ;
    wire signal_9027 ;
    wire signal_9028 ;
    wire signal_9029 ;
    wire signal_9030 ;
    wire signal_9031 ;
    wire signal_9032 ;
    wire signal_9033 ;
    wire signal_9034 ;
    wire signal_9035 ;
    wire signal_9036 ;
    wire signal_9037 ;
    wire signal_9038 ;
    wire signal_9039 ;
    wire signal_9040 ;
    wire signal_9041 ;
    wire signal_9042 ;
    wire signal_9043 ;
    wire signal_9044 ;
    wire signal_9045 ;
    wire signal_9046 ;
    wire signal_9047 ;
    wire signal_9048 ;
    wire signal_9049 ;
    wire signal_9050 ;
    wire signal_9051 ;
    wire signal_9052 ;
    wire signal_9053 ;
    wire signal_9054 ;
    wire signal_9055 ;
    wire signal_9056 ;
    wire signal_9057 ;
    wire signal_9058 ;
    wire signal_9059 ;
    wire signal_9060 ;
    wire signal_9061 ;
    wire signal_9062 ;
    wire signal_9063 ;
    wire signal_9064 ;
    wire signal_9065 ;
    wire signal_9066 ;
    wire signal_9067 ;
    wire signal_9068 ;
    wire signal_9069 ;
    wire signal_9070 ;
    wire signal_9071 ;
    wire signal_9072 ;
    wire signal_9073 ;
    wire signal_9074 ;
    wire signal_9075 ;
    wire signal_9076 ;
    wire signal_9077 ;
    wire signal_9078 ;
    wire signal_9079 ;
    wire signal_9080 ;
    wire signal_9081 ;
    wire signal_9082 ;
    wire signal_9083 ;
    wire signal_9084 ;
    wire signal_9085 ;
    wire signal_9086 ;
    wire signal_9087 ;
    wire signal_9088 ;
    wire signal_9089 ;
    wire signal_9090 ;
    wire signal_9091 ;
    wire signal_9092 ;
    wire signal_9093 ;
    wire signal_9094 ;
    wire signal_9095 ;
    wire signal_9096 ;
    wire signal_9097 ;
    wire signal_9098 ;
    wire signal_9099 ;
    wire signal_9100 ;
    wire signal_9101 ;
    wire signal_9102 ;
    wire signal_9103 ;
    wire signal_9104 ;
    wire signal_9105 ;
    wire signal_9106 ;
    wire signal_9107 ;
    wire signal_9108 ;
    wire signal_9109 ;
    wire signal_9110 ;
    wire signal_9111 ;
    wire signal_9112 ;
    wire signal_9113 ;
    wire signal_9114 ;
    wire signal_9115 ;
    wire signal_9116 ;
    wire signal_9117 ;
    wire signal_9118 ;
    wire signal_9119 ;
    wire signal_9120 ;
    wire signal_9121 ;
    wire signal_9122 ;
    wire signal_9123 ;
    wire signal_9124 ;
    wire signal_9125 ;
    wire signal_9126 ;
    wire signal_9127 ;
    wire signal_9128 ;
    wire signal_9129 ;
    wire signal_9130 ;
    wire signal_9131 ;
    wire signal_9132 ;
    wire signal_9133 ;
    wire signal_9134 ;
    wire signal_9135 ;
    wire signal_9136 ;
    wire signal_9137 ;
    wire signal_9138 ;
    wire signal_9139 ;
    wire signal_9140 ;
    wire signal_9141 ;
    wire signal_9142 ;
    wire signal_9143 ;
    wire signal_9144 ;
    wire signal_9145 ;
    wire signal_9146 ;
    wire signal_9147 ;
    wire signal_9148 ;
    wire signal_9149 ;
    wire signal_9150 ;
    wire signal_9151 ;
    wire signal_9152 ;
    wire signal_9153 ;
    wire signal_9154 ;
    wire signal_9155 ;
    wire signal_9156 ;
    wire signal_9157 ;
    wire signal_9158 ;
    wire signal_9159 ;
    wire signal_9160 ;
    wire signal_9161 ;
    wire signal_9162 ;
    wire signal_9163 ;
    wire signal_9164 ;
    wire signal_9165 ;
    wire signal_9166 ;
    wire signal_9167 ;
    wire signal_9168 ;
    wire signal_9169 ;
    wire signal_9170 ;
    wire signal_9171 ;
    wire signal_9172 ;
    wire signal_9173 ;
    wire signal_9174 ;
    wire signal_9175 ;
    wire signal_9176 ;
    wire signal_9177 ;
    wire signal_9178 ;
    wire signal_9179 ;
    wire signal_9180 ;
    wire signal_9181 ;
    wire signal_9182 ;
    wire signal_9183 ;
    wire signal_9184 ;
    wire signal_9185 ;
    wire signal_9186 ;
    wire signal_9187 ;
    wire signal_9188 ;
    wire signal_9189 ;
    wire signal_9190 ;
    wire signal_9191 ;
    wire signal_9192 ;
    wire signal_9193 ;
    wire signal_9194 ;
    wire signal_9195 ;
    wire signal_9196 ;
    wire signal_9197 ;
    wire signal_9198 ;
    wire signal_9199 ;
    wire signal_9200 ;
    wire signal_9201 ;
    wire signal_9202 ;
    wire signal_9203 ;
    wire signal_9204 ;
    wire signal_9205 ;
    wire signal_9206 ;
    wire signal_9207 ;
    wire signal_9208 ;
    wire signal_9209 ;
    wire signal_9210 ;
    wire signal_9211 ;
    wire signal_9212 ;
    wire signal_9213 ;
    wire signal_9214 ;
    wire signal_9215 ;
    wire signal_9216 ;
    wire signal_9217 ;
    wire signal_9218 ;
    wire signal_9219 ;
    wire signal_9220 ;
    wire signal_9221 ;
    wire signal_9222 ;
    wire signal_9223 ;
    wire signal_9224 ;
    wire signal_9225 ;
    wire signal_9226 ;
    wire signal_9227 ;
    wire signal_9228 ;
    wire signal_9229 ;
    wire signal_9230 ;
    wire signal_9231 ;
    wire signal_9232 ;
    wire signal_9233 ;
    wire signal_9234 ;
    wire signal_9235 ;
    wire signal_9236 ;
    wire signal_9237 ;
    wire signal_9238 ;
    wire signal_9239 ;
    wire signal_9240 ;
    wire signal_9241 ;
    wire signal_9242 ;
    wire signal_9243 ;
    wire signal_9244 ;
    wire signal_9245 ;
    wire signal_9246 ;
    wire signal_9247 ;
    wire signal_9248 ;
    wire signal_9249 ;
    wire signal_9250 ;
    wire signal_9251 ;
    wire signal_9252 ;
    wire signal_9253 ;
    wire signal_9254 ;
    wire signal_9255 ;
    wire signal_9256 ;
    wire signal_9257 ;
    wire signal_9258 ;
    wire signal_9259 ;
    wire signal_9260 ;
    wire signal_9261 ;
    wire signal_9262 ;
    wire signal_9263 ;
    wire signal_9264 ;
    wire signal_9265 ;
    wire signal_9266 ;
    wire signal_9267 ;
    wire signal_9268 ;
    wire signal_9269 ;
    wire signal_9270 ;
    wire signal_9271 ;
    wire signal_9272 ;
    wire signal_9273 ;
    wire signal_9274 ;
    wire signal_9275 ;
    wire signal_9276 ;
    wire signal_9277 ;
    wire signal_9278 ;
    wire signal_9279 ;
    wire signal_9280 ;
    wire signal_9281 ;
    wire signal_9282 ;
    wire signal_9283 ;
    wire signal_9284 ;
    wire signal_9285 ;
    wire signal_9286 ;
    wire signal_9287 ;
    wire signal_9288 ;
    wire signal_9289 ;
    wire signal_9290 ;
    wire signal_9291 ;
    wire signal_9292 ;
    wire signal_9293 ;
    wire signal_9294 ;
    wire signal_9295 ;
    wire signal_9296 ;
    wire signal_9297 ;
    wire signal_9298 ;
    wire signal_9299 ;
    wire signal_9300 ;
    wire signal_9301 ;
    wire signal_9302 ;
    wire signal_9303 ;
    wire signal_9304 ;
    wire signal_9305 ;
    wire signal_9306 ;
    wire signal_9307 ;
    wire signal_9308 ;
    wire signal_9309 ;
    wire signal_9310 ;
    wire signal_9311 ;
    wire signal_9312 ;
    wire signal_9313 ;
    wire signal_9314 ;
    wire signal_9315 ;
    wire signal_9316 ;
    wire signal_9317 ;
    wire signal_9318 ;
    wire signal_9319 ;
    wire signal_9320 ;
    wire signal_9321 ;
    wire signal_9322 ;
    wire signal_9323 ;
    wire signal_9324 ;
    wire signal_9325 ;
    wire signal_9326 ;
    wire signal_9327 ;
    wire signal_9328 ;
    wire signal_9329 ;
    wire signal_9330 ;
    wire signal_9331 ;
    wire signal_9332 ;
    wire signal_9333 ;
    wire signal_9334 ;
    wire signal_9335 ;
    wire signal_9336 ;
    wire signal_9337 ;
    wire signal_9338 ;
    wire signal_9339 ;
    wire signal_9340 ;
    wire signal_9341 ;
    wire signal_9342 ;
    wire signal_9343 ;
    wire signal_9344 ;
    wire signal_9345 ;
    wire signal_9346 ;
    wire signal_9347 ;
    wire signal_9348 ;
    wire signal_9349 ;
    wire signal_9350 ;
    wire signal_9351 ;
    wire signal_9352 ;
    wire signal_9353 ;
    wire signal_9354 ;
    wire signal_9355 ;
    wire signal_9356 ;
    wire signal_9357 ;
    wire signal_9358 ;
    wire signal_9359 ;
    wire signal_9360 ;
    wire signal_9361 ;
    wire signal_9362 ;
    wire signal_9363 ;
    wire signal_9364 ;
    wire signal_9365 ;
    wire signal_9366 ;
    wire signal_9367 ;
    wire signal_9368 ;
    wire signal_9369 ;
    wire signal_9370 ;
    wire signal_9371 ;
    wire signal_9372 ;
    wire signal_9373 ;
    wire signal_9374 ;
    wire signal_9375 ;
    wire signal_9376 ;
    wire signal_9377 ;
    wire signal_9378 ;
    wire signal_9379 ;
    wire signal_9380 ;
    wire signal_9381 ;
    wire signal_9382 ;
    wire signal_9383 ;
    wire signal_9384 ;
    wire signal_9385 ;
    wire signal_9386 ;
    wire signal_9387 ;
    wire signal_9388 ;
    wire signal_9389 ;
    wire signal_9390 ;
    wire signal_9391 ;
    wire signal_9392 ;
    wire signal_9393 ;
    wire signal_9394 ;
    wire signal_9395 ;
    wire signal_9396 ;
    wire signal_9397 ;
    wire signal_9398 ;
    wire signal_9399 ;
    wire signal_9400 ;
    wire signal_9401 ;
    wire signal_9402 ;
    wire signal_9403 ;
    wire signal_9404 ;
    wire signal_9405 ;
    wire signal_9406 ;
    wire signal_9407 ;
    wire signal_9408 ;
    wire signal_9409 ;
    wire signal_9410 ;
    wire signal_9411 ;
    wire signal_9412 ;
    wire signal_9413 ;
    wire signal_9414 ;
    wire signal_9415 ;
    wire signal_9416 ;
    wire signal_9417 ;
    wire signal_9418 ;
    wire signal_9419 ;
    wire signal_9420 ;
    wire signal_9421 ;
    wire signal_9422 ;
    wire signal_9423 ;
    wire signal_9424 ;
    wire signal_9425 ;
    wire signal_9426 ;
    wire signal_9427 ;
    wire signal_9428 ;
    wire signal_9429 ;
    wire signal_9430 ;
    wire signal_9431 ;
    wire signal_9432 ;
    wire signal_9433 ;
    wire signal_9434 ;
    wire signal_9435 ;
    wire signal_9436 ;
    wire signal_9437 ;
    wire signal_9438 ;
    wire signal_9439 ;
    wire signal_9440 ;
    wire signal_9441 ;
    wire signal_9442 ;
    wire signal_9443 ;
    wire signal_9444 ;
    wire signal_9445 ;
    wire signal_9446 ;
    wire signal_9447 ;
    wire signal_9448 ;
    wire signal_9449 ;
    wire signal_9450 ;
    wire signal_9451 ;
    wire signal_9452 ;
    wire signal_9453 ;
    wire signal_9454 ;
    wire signal_9455 ;
    wire signal_9456 ;
    wire signal_9457 ;
    wire signal_9458 ;
    wire signal_9459 ;
    wire signal_9460 ;
    wire signal_9461 ;
    wire signal_9462 ;
    wire signal_9463 ;
    wire signal_9464 ;
    wire signal_9465 ;
    wire signal_9466 ;
    wire signal_9467 ;
    wire signal_9468 ;
    wire signal_9469 ;
    wire signal_9470 ;
    wire signal_9471 ;
    wire signal_9472 ;
    wire signal_9473 ;
    wire signal_9474 ;
    wire signal_9475 ;
    wire signal_9476 ;
    wire signal_9477 ;
    wire signal_9478 ;
    wire signal_9479 ;
    wire signal_9480 ;
    wire signal_9481 ;
    wire signal_9482 ;
    wire signal_9483 ;
    wire signal_9484 ;
    wire signal_9485 ;
    wire signal_9486 ;
    wire signal_9487 ;
    wire signal_9488 ;
    wire signal_9489 ;
    wire signal_9490 ;
    wire signal_9491 ;
    wire signal_9492 ;
    wire signal_9493 ;
    wire signal_9494 ;
    wire signal_9495 ;
    wire signal_9496 ;
    wire signal_9497 ;
    wire signal_9498 ;
    wire signal_9499 ;
    wire signal_9500 ;
    wire signal_9501 ;
    wire signal_9502 ;
    wire signal_9503 ;
    wire signal_9504 ;
    wire signal_9505 ;
    wire signal_9506 ;
    wire signal_9507 ;
    wire signal_9508 ;
    wire signal_9509 ;
    wire signal_9510 ;
    wire signal_9511 ;
    wire signal_9512 ;
    wire signal_9513 ;
    wire signal_9514 ;
    wire signal_9515 ;
    wire signal_9516 ;
    wire signal_9517 ;
    wire signal_9518 ;
    wire signal_9519 ;
    wire signal_9520 ;
    wire signal_9521 ;
    wire signal_9522 ;
    wire signal_9523 ;
    wire signal_9524 ;
    wire signal_9525 ;
    wire signal_9526 ;
    wire signal_9527 ;
    wire signal_9528 ;
    wire signal_9529 ;
    wire signal_9530 ;
    wire signal_9531 ;
    wire signal_9532 ;
    wire signal_9533 ;
    wire signal_9534 ;
    wire signal_9535 ;
    wire signal_9536 ;
    wire signal_9537 ;
    wire signal_9538 ;
    wire signal_9539 ;
    wire signal_9540 ;
    wire signal_9541 ;
    wire signal_9542 ;
    wire signal_9543 ;
    wire signal_9544 ;
    wire signal_9545 ;
    wire signal_9546 ;
    wire signal_9547 ;
    wire signal_9548 ;
    wire signal_9549 ;
    wire signal_9550 ;
    wire signal_9551 ;
    wire signal_9552 ;
    wire signal_9553 ;
    wire signal_9554 ;
    wire signal_9555 ;
    wire signal_9556 ;
    wire signal_9557 ;
    wire signal_9558 ;
    wire signal_9559 ;
    wire signal_9560 ;
    wire signal_9561 ;
    wire signal_9562 ;
    wire signal_9563 ;
    wire signal_9564 ;
    wire signal_9565 ;
    wire signal_9566 ;
    wire signal_9567 ;
    wire signal_9568 ;
    wire signal_9569 ;
    wire signal_9570 ;
    wire signal_9571 ;
    wire signal_9572 ;
    wire signal_9573 ;
    wire signal_9574 ;
    wire signal_9575 ;
    wire signal_9576 ;
    wire signal_9577 ;
    wire signal_9578 ;
    wire signal_9579 ;
    wire signal_9580 ;
    wire signal_9581 ;
    wire signal_9582 ;
    wire signal_9583 ;
    wire signal_9584 ;
    wire signal_9585 ;
    wire signal_9586 ;
    wire signal_9587 ;
    wire signal_9588 ;
    wire signal_9589 ;
    wire signal_9590 ;
    wire signal_9591 ;
    wire signal_9592 ;
    wire signal_9593 ;
    wire signal_9594 ;
    wire signal_9595 ;
    wire signal_9596 ;
    wire signal_9597 ;
    wire signal_9598 ;
    wire signal_9599 ;
    wire signal_9600 ;
    wire signal_9601 ;
    wire signal_9602 ;
    wire signal_9603 ;
    wire signal_9604 ;
    wire signal_9605 ;
    wire signal_9606 ;
    wire signal_9607 ;
    wire signal_9608 ;
    wire signal_9609 ;
    wire signal_9610 ;
    wire signal_9611 ;
    wire signal_9612 ;
    wire signal_9613 ;
    wire signal_9614 ;
    wire signal_9615 ;
    wire signal_9616 ;
    wire signal_9617 ;
    wire signal_9618 ;
    wire signal_9619 ;
    wire signal_9620 ;
    wire signal_9621 ;
    wire signal_9622 ;
    wire signal_9623 ;
    wire signal_9624 ;
    wire signal_9625 ;
    wire signal_9626 ;
    wire signal_9627 ;
    wire signal_9628 ;
    wire signal_9629 ;
    wire signal_9630 ;
    wire signal_9631 ;
    wire signal_9632 ;
    wire signal_9633 ;
    wire signal_9634 ;
    wire signal_9635 ;
    wire signal_9636 ;
    wire signal_9637 ;
    wire signal_9638 ;
    wire signal_9639 ;
    wire signal_9640 ;
    wire signal_9641 ;
    wire signal_9642 ;
    wire signal_9643 ;
    wire signal_9644 ;
    wire signal_9645 ;
    wire signal_9646 ;
    wire signal_9647 ;
    wire signal_9648 ;
    wire signal_9649 ;
    wire signal_9650 ;
    wire signal_9651 ;
    wire signal_9652 ;
    wire signal_9653 ;
    wire signal_9654 ;
    wire signal_9655 ;
    wire signal_9656 ;
    wire signal_9657 ;
    wire signal_9658 ;
    wire signal_9659 ;
    wire signal_9660 ;
    wire signal_9661 ;
    wire signal_9662 ;
    wire signal_9663 ;
    wire signal_9664 ;
    wire signal_9665 ;
    wire signal_9666 ;
    wire signal_9667 ;
    wire signal_9668 ;
    wire signal_9669 ;
    wire signal_9670 ;
    wire signal_9671 ;
    wire signal_9672 ;
    wire signal_9673 ;
    wire signal_9674 ;
    wire signal_9675 ;
    wire signal_9676 ;
    wire signal_9677 ;
    wire signal_9678 ;
    wire signal_9679 ;
    wire signal_9680 ;
    wire signal_9681 ;
    wire signal_9682 ;
    wire signal_9683 ;
    wire signal_9684 ;
    wire signal_9685 ;
    wire signal_9686 ;
    wire signal_9687 ;
    wire signal_9688 ;
    wire signal_9689 ;
    wire signal_9690 ;
    wire signal_9691 ;
    wire signal_9692 ;
    wire signal_9693 ;
    wire signal_9694 ;
    wire signal_9695 ;
    wire signal_9696 ;
    wire signal_9697 ;
    wire signal_9698 ;
    wire signal_9699 ;
    wire signal_9700 ;
    wire signal_9701 ;
    wire signal_9702 ;
    wire signal_9703 ;
    wire signal_9704 ;
    wire signal_9705 ;
    wire signal_9706 ;
    wire signal_9707 ;
    wire signal_9708 ;
    wire signal_9709 ;
    wire signal_9710 ;
    wire signal_9711 ;
    wire signal_9712 ;
    wire signal_9713 ;
    wire signal_9714 ;
    wire signal_9715 ;
    wire signal_9716 ;
    wire signal_9717 ;
    wire signal_9718 ;
    wire signal_9719 ;
    wire signal_9720 ;
    wire signal_9721 ;
    wire signal_9722 ;
    wire signal_9723 ;
    wire signal_9724 ;
    wire signal_9725 ;
    wire signal_9726 ;
    wire signal_9727 ;
    wire signal_9728 ;
    wire signal_9729 ;
    wire signal_9730 ;
    wire signal_9731 ;
    wire signal_9732 ;
    wire signal_9733 ;
    wire signal_9734 ;
    wire signal_9735 ;
    wire signal_9736 ;
    wire signal_9737 ;
    wire signal_9738 ;
    wire signal_9739 ;
    wire signal_9740 ;
    wire signal_9741 ;
    wire signal_9742 ;
    wire signal_9743 ;
    wire signal_9744 ;
    wire signal_9745 ;
    wire signal_9746 ;
    wire signal_9747 ;
    wire signal_9748 ;
    wire signal_9749 ;
    wire signal_9750 ;
    wire signal_9751 ;
    wire signal_9752 ;
    wire signal_9753 ;
    wire signal_9754 ;
    wire signal_9755 ;
    wire signal_9756 ;
    wire signal_9757 ;
    wire signal_9758 ;
    wire signal_9759 ;
    wire signal_9760 ;
    wire signal_9761 ;
    wire signal_9762 ;
    wire signal_9763 ;
    wire signal_9764 ;
    wire signal_9765 ;
    wire signal_9766 ;
    wire signal_9767 ;
    wire signal_9768 ;
    wire signal_9769 ;
    wire signal_9770 ;
    wire signal_9771 ;
    wire signal_9772 ;
    wire signal_9773 ;
    wire signal_9774 ;
    wire signal_9775 ;
    wire signal_9776 ;
    wire signal_9777 ;
    wire signal_9778 ;
    wire signal_9779 ;
    wire signal_9780 ;
    wire signal_9781 ;
    wire signal_9782 ;
    wire signal_9783 ;
    wire signal_9784 ;
    wire signal_9785 ;
    wire signal_9786 ;
    wire signal_9787 ;
    wire signal_9788 ;
    wire signal_9789 ;
    wire signal_9790 ;
    wire signal_9791 ;
    wire signal_9792 ;
    wire signal_9793 ;
    wire signal_9794 ;
    wire signal_9795 ;
    wire signal_9796 ;
    wire signal_9797 ;
    wire signal_9798 ;
    wire signal_9799 ;
    wire signal_9800 ;
    wire signal_9801 ;
    wire signal_9802 ;
    wire signal_9803 ;
    wire signal_9804 ;
    wire signal_9805 ;
    wire signal_9806 ;
    wire signal_9807 ;
    wire signal_9808 ;
    wire signal_9809 ;
    wire signal_9810 ;
    wire signal_9811 ;
    wire signal_9812 ;
    wire signal_9813 ;
    wire signal_9814 ;
    wire signal_9815 ;
    wire signal_9816 ;
    wire signal_9817 ;
    wire signal_9818 ;
    wire signal_9819 ;
    wire signal_9820 ;
    wire signal_9821 ;
    wire signal_9822 ;
    wire signal_9823 ;
    wire signal_9824 ;
    wire signal_9825 ;
    wire signal_9826 ;
    wire signal_9827 ;
    wire signal_9828 ;
    wire signal_9829 ;
    wire signal_9830 ;
    wire signal_9831 ;
    wire signal_9832 ;
    wire signal_9833 ;
    wire signal_9834 ;
    wire signal_9835 ;
    wire signal_9836 ;
    wire signal_9837 ;
    wire signal_9838 ;
    wire signal_9839 ;
    wire signal_9840 ;
    wire signal_9841 ;
    wire signal_9842 ;
    wire signal_9843 ;
    wire signal_9844 ;
    wire signal_9845 ;
    wire signal_9846 ;
    wire signal_9847 ;
    wire signal_9848 ;
    wire signal_9849 ;
    wire signal_9850 ;
    wire signal_9851 ;
    wire signal_9852 ;
    wire signal_9853 ;
    wire signal_9854 ;
    wire signal_9855 ;
    wire signal_9856 ;
    wire signal_9857 ;
    wire signal_9858 ;
    wire signal_9859 ;
    wire signal_9860 ;
    wire signal_9861 ;
    wire signal_9862 ;
    wire signal_9863 ;
    wire signal_9864 ;
    wire signal_9865 ;
    wire signal_9866 ;
    wire signal_9867 ;
    wire signal_9868 ;
    wire signal_9869 ;
    wire signal_9870 ;
    wire signal_9871 ;
    wire signal_9872 ;
    wire signal_9873 ;
    wire signal_9874 ;
    wire signal_9875 ;
    wire signal_9876 ;
    wire signal_9877 ;
    wire signal_9878 ;
    wire signal_9879 ;
    wire signal_9880 ;
    wire signal_9881 ;
    wire signal_9882 ;
    wire signal_9883 ;
    wire signal_9884 ;
    wire signal_9885 ;
    wire signal_9886 ;
    wire signal_9887 ;
    wire signal_9888 ;
    wire signal_9889 ;
    wire signal_9890 ;
    wire signal_9891 ;
    wire signal_9892 ;
    wire signal_9893 ;
    wire signal_9894 ;
    wire signal_9895 ;
    wire signal_9896 ;
    wire signal_9897 ;
    wire signal_9898 ;
    wire signal_9899 ;
    wire signal_9900 ;
    wire signal_9901 ;
    wire signal_9902 ;
    wire signal_9903 ;
    wire signal_9904 ;
    wire signal_9905 ;
    wire signal_9906 ;
    wire signal_9907 ;
    wire signal_9908 ;
    wire signal_9909 ;
    wire signal_9910 ;
    wire signal_9911 ;
    wire signal_9912 ;
    wire signal_9913 ;
    wire signal_9914 ;
    wire signal_9915 ;
    wire signal_9916 ;
    wire signal_9917 ;
    wire signal_9918 ;
    wire signal_9919 ;
    wire signal_9920 ;
    wire signal_9921 ;
    wire signal_9922 ;
    wire signal_9923 ;
    wire signal_9924 ;
    wire signal_9925 ;
    wire signal_9926 ;
    wire signal_9927 ;
    wire signal_9928 ;
    wire signal_9929 ;
    wire signal_9930 ;
    wire signal_9931 ;
    wire signal_9932 ;
    wire signal_9933 ;
    wire signal_9934 ;
    wire signal_9935 ;
    wire signal_9936 ;
    wire signal_9937 ;
    wire signal_9938 ;
    wire signal_9939 ;
    wire signal_9940 ;
    wire signal_9941 ;
    wire signal_9942 ;
    wire signal_9943 ;
    wire signal_9944 ;
    wire signal_9945 ;
    wire signal_9946 ;
    wire signal_9947 ;
    wire signal_9948 ;
    wire signal_9949 ;
    wire signal_9950 ;
    wire signal_9951 ;
    wire signal_9952 ;
    wire signal_9953 ;
    wire signal_9954 ;
    wire signal_9955 ;
    wire signal_9956 ;
    wire signal_9957 ;
    wire signal_9958 ;
    wire signal_9959 ;
    wire signal_9960 ;
    wire signal_9961 ;
    wire signal_9962 ;
    wire signal_9963 ;
    wire signal_9964 ;
    wire signal_9965 ;
    wire signal_9966 ;
    wire signal_9967 ;
    wire signal_9968 ;
    wire signal_9969 ;
    wire signal_9970 ;
    wire signal_9971 ;
    wire signal_9972 ;
    wire signal_9973 ;
    wire signal_9974 ;
    wire signal_9975 ;
    wire signal_9976 ;
    wire signal_9977 ;
    wire signal_9978 ;
    wire signal_9979 ;
    wire signal_9980 ;
    wire signal_9981 ;
    wire signal_9982 ;
    wire signal_9983 ;
    wire signal_9984 ;
    wire signal_9985 ;
    wire signal_9986 ;
    wire signal_9987 ;
    wire signal_9988 ;
    wire signal_9989 ;
    wire signal_9990 ;
    wire signal_9991 ;
    wire signal_9992 ;
    wire signal_9993 ;
    wire signal_9994 ;
    wire signal_9995 ;
    wire signal_9996 ;
    wire signal_9997 ;
    wire signal_9998 ;
    wire signal_9999 ;
    wire signal_10000 ;
    wire signal_10001 ;
    wire signal_10002 ;
    wire signal_10003 ;
    wire signal_10004 ;
    wire signal_10005 ;
    wire signal_10006 ;
    wire signal_10007 ;
    wire signal_10008 ;
    wire signal_10009 ;
    wire signal_10010 ;
    wire signal_10011 ;
    wire signal_10012 ;
    wire signal_10013 ;
    wire signal_10014 ;
    wire signal_10015 ;
    wire signal_10016 ;
    wire signal_10017 ;
    wire signal_10018 ;
    wire signal_10019 ;
    wire signal_10020 ;
    wire signal_10021 ;
    wire signal_10022 ;
    wire signal_10023 ;
    wire signal_10024 ;
    wire signal_10025 ;
    wire signal_10026 ;
    wire signal_10027 ;
    wire signal_10028 ;
    wire signal_10029 ;
    wire signal_10030 ;
    wire signal_10031 ;
    wire signal_10032 ;
    wire signal_10033 ;
    wire signal_10034 ;
    wire signal_10035 ;
    wire signal_10036 ;
    wire signal_10037 ;
    wire signal_10038 ;
    wire signal_10039 ;
    wire signal_10040 ;
    wire signal_10041 ;
    wire signal_10042 ;
    wire signal_10043 ;
    wire signal_10044 ;
    wire signal_10045 ;
    wire signal_10046 ;
    wire signal_10047 ;
    wire signal_10048 ;
    wire signal_10049 ;
    wire signal_10050 ;
    wire signal_10051 ;
    wire signal_10052 ;
    wire signal_10053 ;
    wire signal_10054 ;
    wire signal_10055 ;
    wire signal_10056 ;
    wire signal_10057 ;
    wire signal_10058 ;
    wire signal_10059 ;
    wire signal_10060 ;
    wire signal_10061 ;
    wire signal_10062 ;
    wire signal_10063 ;
    wire signal_10064 ;
    wire signal_10065 ;
    wire signal_10066 ;
    wire signal_10067 ;
    wire signal_10068 ;
    wire signal_10069 ;
    wire signal_10070 ;
    wire signal_10071 ;
    wire signal_10072 ;
    wire signal_10073 ;
    wire signal_10074 ;
    wire signal_10075 ;
    wire signal_10076 ;
    wire signal_10077 ;
    wire signal_10078 ;
    wire signal_10079 ;
    wire signal_10080 ;
    wire signal_10081 ;
    wire signal_10082 ;
    wire signal_10083 ;
    wire signal_10084 ;
    wire signal_10085 ;
    wire signal_10086 ;
    wire signal_10087 ;
    wire signal_10088 ;
    wire signal_10089 ;
    wire signal_10090 ;
    wire signal_10091 ;
    wire signal_10092 ;
    wire signal_10093 ;
    wire signal_10094 ;
    wire signal_10095 ;
    wire signal_10096 ;
    wire signal_10097 ;
    wire signal_10098 ;
    wire signal_10099 ;
    wire signal_10100 ;
    wire signal_10101 ;

    /* cells in depth 0 */
    NOR2_X1 cell_0 ( .A1 (signal_875), .A2 (signal_878), .ZN (signal_266) ) ;
    NAND2_X1 cell_1 ( .A1 (signal_879), .A2 (signal_266), .ZN (signal_267) ) ;
    NOR2_X1 cell_2 ( .A1 (signal_874), .A2 (signal_267), .ZN (signal_268) ) ;
    NAND2_X1 cell_3 ( .A1 (signal_876), .A2 (signal_268), .ZN (signal_269) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_877), .A2 (signal_269), .ZN (signal_270) ) ;
    NOR2_X1 cell_5 ( .A1 (OUT_done), .A2 (signal_270), .ZN (signal_271) ) ;
    NOR2_X1 cell_6 ( .A1 (IN_reset), .A2 (signal_271), .ZN (signal_265) ) ;
    NAND2_X1 cell_7 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_272) ) ;
    XNOR2_X1 cell_8 ( .A (signal_304), .B (signal_275), .ZN (signal_274) ) ;
    XOR2_X1 cell_9 ( .A (signal_309), .B (signal_307), .Z (signal_275) ) ;
    NAND2_X1 cell_10 ( .A1 (signal_276), .A2 (signal_277), .ZN (signal_273) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_278), .A2 (signal_279), .ZN (signal_277) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_302), .A2 (signal_289), .ZN (signal_279) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_278) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_289), .A2 (signal_280), .ZN (signal_276) ) ;
    AND2_X1 cell_15 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_280) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_298), .A2 (signal_283), .ZN (signal_282) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_300), .A2 (signal_284), .ZN (signal_283) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_296), .A2 (signal_876), .ZN (signal_284) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_292), .A2 (signal_290), .ZN (signal_281) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_292), .A2 (IN_reset), .ZN (signal_291) ) ;
    NOR2_X1 cell_21 ( .A1 (IN_reset), .A2 (signal_294), .ZN (signal_293) ) ;
    NOR2_X1 cell_22 ( .A1 (IN_reset), .A2 (signal_296), .ZN (signal_295) ) ;
    NOR2_X1 cell_23 ( .A1 (IN_reset), .A2 (signal_298), .ZN (signal_297) ) ;
    NOR2_X1 cell_24 ( .A1 (IN_reset), .A2 (signal_300), .ZN (signal_299) ) ;
    NOR2_X1 cell_25 ( .A1 (signal_289), .A2 (IN_reset), .ZN (signal_303) ) ;
    NOR2_X1 cell_26 ( .A1 (signal_306), .A2 (IN_reset), .ZN (signal_305) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_309), .A2 (IN_reset), .ZN (signal_308) ) ;
    NOR2_X1 cell_28 ( .A1 (signal_288), .A2 (IN_reset), .ZN (signal_310) ) ;
    OR2_X1 cell_29 ( .A1 (signal_288), .A2 (signal_276), .ZN (signal_286) ) ;
    NAND2_X1 cell_30 ( .A1 (signal_272), .A2 (signal_286), .ZN (signal_311) ) ;
    NOR2_X1 cell_31 ( .A1 (signal_281), .A2 (signal_282), .ZN (signal_340) ) ;
    INV_X1 cell_32 ( .A (signal_286), .ZN (signal_285) ) ;
    OR2_X1 cell_33 ( .A1 (IN_reset), .A2 (signal_287), .ZN (signal_301) ) ;
    XNOR2_X1 cell_34 ( .A (signal_292), .B (signal_290), .ZN (signal_287) ) ;
    INV_X1 cell_35 ( .A (signal_340), .ZN (signal_341) ) ;
    INV_X1 cell_36 ( .A (signal_341), .ZN (signal_344) ) ;
    INV_X1 cell_37 ( .A (signal_341), .ZN (signal_342) ) ;
    INV_X1 cell_38 ( .A (signal_341), .ZN (signal_343) ) ;
    INV_X1 cell_167 ( .A (signal_345), .ZN (signal_346) ) ;
    INV_X1 cell_168 ( .A (signal_285), .ZN (signal_345) ) ;
    INV_X1 cell_169 ( .A (signal_345), .ZN (signal_348) ) ;
    INV_X1 cell_170 ( .A (signal_345), .ZN (signal_347) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_171 ( .s (signal_285), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({signal_1856, signal_1135}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_172 ( .s (signal_346), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({signal_1921, signal_1134}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_173 ( .s (signal_346), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({signal_1924, signal_1133}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_174 ( .s (signal_285), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({signal_1859, signal_1132}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_175 ( .s (signal_346), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({signal_1927, signal_1131}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_176 ( .s (signal_346), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({signal_1930, signal_1130}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_177 ( .s (signal_346), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({signal_1933, signal_1129}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_178 ( .s (signal_346), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({signal_1936, signal_1128}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_179 ( .s (signal_346), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({signal_1939, signal_1127}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_180 ( .s (signal_346), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({signal_1942, signal_1126}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_181 ( .s (signal_346), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({signal_1945, signal_1125}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_182 ( .s (signal_346), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({signal_1948, signal_1124}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_183 ( .s (signal_346), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({signal_1951, signal_1123}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_184 ( .s (signal_346), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({signal_1954, signal_1122}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_185 ( .s (signal_346), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({signal_1957, signal_1121}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_186 ( .s (signal_346), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({signal_1960, signal_1120}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_187 ( .s (signal_285), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({signal_1862, signal_1119}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_188 ( .s (signal_347), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({signal_1963, signal_1118}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_189 ( .s (signal_348), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({signal_1966, signal_1117}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_190 ( .s (signal_285), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({signal_1865, signal_1116}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_191 ( .s (signal_346), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({signal_1969, signal_1115}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_192 ( .s (signal_348), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({signal_1972, signal_1114}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_193 ( .s (signal_285), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({signal_1868, signal_1113}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_194 ( .s (signal_348), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({signal_1975, signal_1112}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_195 ( .s (signal_285), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({signal_1871, signal_1111}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_196 ( .s (signal_348), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({signal_1978, signal_1110}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_197 ( .s (signal_285), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({signal_1874, signal_1109}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_198 ( .s (signal_348), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({signal_1981, signal_1108}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_199 ( .s (signal_285), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({signal_1877, signal_1107}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_200 ( .s (signal_347), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({signal_1984, signal_1106}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_201 ( .s (signal_347), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({signal_1987, signal_1105}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_202 ( .s (signal_347), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({signal_1990, signal_1104}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_203 ( .s (signal_285), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({signal_1880, signal_1103}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_204 ( .s (signal_348), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({signal_1993, signal_1102}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_205 ( .s (signal_285), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({signal_1883, signal_1101}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_206 ( .s (signal_285), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({signal_1886, signal_1100}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_207 ( .s (signal_285), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({signal_1889, signal_1099}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_208 ( .s (signal_347), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({signal_1996, signal_1098}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_209 ( .s (signal_347), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({signal_1999, signal_1097}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_210 ( .s (signal_285), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({signal_1892, signal_1096}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_211 ( .s (signal_347), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({signal_2002, signal_1095}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_212 ( .s (signal_347), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({signal_2005, signal_1094}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_213 ( .s (signal_347), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({signal_2008, signal_1093}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_214 ( .s (signal_347), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({signal_2011, signal_1092}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_215 ( .s (signal_347), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({signal_2014, signal_1091}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_216 ( .s (signal_347), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({signal_2017, signal_1090}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_217 ( .s (signal_347), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({signal_2020, signal_1089}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_218 ( .s (signal_347), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({signal_2023, signal_1088}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_219 ( .s (signal_347), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({signal_2026, signal_1087}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_220 ( .s (signal_347), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({signal_2029, signal_1086}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_221 ( .s (signal_347), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({signal_2032, signal_1085}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_222 ( .s (signal_347), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({signal_2035, signal_1084}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_223 ( .s (signal_348), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({signal_2038, signal_1083}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_224 ( .s (signal_348), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({signal_2041, signal_1082}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_225 ( .s (signal_348), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({signal_2044, signal_1081}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_226 ( .s (signal_348), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({signal_2047, signal_1080}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_227 ( .s (signal_348), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({signal_2050, signal_1079}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_228 ( .s (signal_348), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({signal_2053, signal_1078}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_229 ( .s (signal_348), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({signal_2056, signal_1077}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_230 ( .s (signal_348), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({signal_2059, signal_1076}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_231 ( .s (signal_348), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({signal_2062, signal_1075}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_232 ( .s (signal_348), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({signal_2065, signal_1074}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_233 ( .s (signal_348), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({signal_2068, signal_1073}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_234 ( .s (signal_348), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({signal_2071, signal_1072}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({signal_1942, signal_1126}), .c ({signal_2080, signal_1062}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({signal_1939, signal_1127}), .c ({signal_2082, signal_1063}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({signal_1936, signal_1128}), .c ({signal_2084, signal_1064}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({signal_1933, signal_1129}), .c ({signal_2086, signal_1065}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({signal_2071, signal_1072}), .c ({signal_2088, signal_1008}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({signal_2068, signal_1073}), .c ({signal_2090, signal_1009}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({signal_2065, signal_1074}), .c ({signal_2092, signal_1010}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({signal_2062, signal_1075}), .c ({signal_2094, signal_1011}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({signal_1930, signal_1130}), .c ({signal_2096, signal_1066}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({signal_2059, signal_1076}), .c ({signal_2098, signal_1012}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({signal_2056, signal_1077}), .c ({signal_2100, signal_1013}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({signal_2053, signal_1078}), .c ({signal_2102, signal_1014}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({signal_2050, signal_1079}), .c ({signal_2104, signal_1015}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({signal_2047, signal_1080}), .c ({signal_2106, signal_1016}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({signal_2044, signal_1081}), .c ({signal_2108, signal_1017}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({signal_2041, signal_1082}), .c ({signal_2110, signal_1018}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({signal_2038, signal_1083}), .c ({signal_2112, signal_1019}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({signal_2035, signal_1084}), .c ({signal_2114, signal_1020}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({signal_2032, signal_1085}), .c ({signal_2116, signal_1021}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({signal_1927, signal_1131}), .c ({signal_2118, signal_1067}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({signal_2029, signal_1086}), .c ({signal_2120, signal_1022}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({signal_2026, signal_1087}), .c ({signal_2122, signal_1023}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_257 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({signal_2023, signal_1088}), .c ({signal_2124, signal_1024}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({signal_2020, signal_1089}), .c ({signal_2126, signal_1025}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({signal_2017, signal_1090}), .c ({signal_2128, signal_1026}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({signal_2014, signal_1091}), .c ({signal_2130, signal_1027}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({signal_2011, signal_1092}), .c ({signal_2132, signal_1028}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({signal_2008, signal_1093}), .c ({signal_2134, signal_1029}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({signal_2005, signal_1094}), .c ({signal_2136, signal_1030}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({signal_2002, signal_1095}), .c ({signal_2138, signal_1031}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({signal_1859, signal_1132}), .c ({signal_1894, signal_1068}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({signal_1892, signal_1096}), .c ({signal_1896, signal_1032}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_267 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({signal_1999, signal_1097}), .c ({signal_2140, signal_1033}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_268 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({signal_1996, signal_1098}), .c ({signal_2142, signal_1034}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({signal_1889, signal_1099}), .c ({signal_1898, signal_1035}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({signal_1886, signal_1100}), .c ({signal_1900, signal_1036}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({signal_1883, signal_1101}), .c ({signal_1902, signal_1037}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({signal_1993, signal_1102}), .c ({signal_2144, signal_1038}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({signal_1880, signal_1103}), .c ({signal_1904, signal_1039}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({signal_1990, signal_1104}), .c ({signal_2146, signal_1040}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({signal_1987, signal_1105}), .c ({signal_2148, signal_1041}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({signal_1924, signal_1133}), .c ({signal_2150, signal_1069}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({signal_1984, signal_1106}), .c ({signal_2152, signal_1042}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({signal_1877, signal_1107}), .c ({signal_1906, signal_1043}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({signal_1981, signal_1108}), .c ({signal_2154, signal_1044}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_280 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({signal_1874, signal_1109}), .c ({signal_1908, signal_1045}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_281 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({signal_1978, signal_1110}), .c ({signal_2156, signal_1046}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_282 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({signal_1871, signal_1111}), .c ({signal_1910, signal_1047}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_283 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({signal_1975, signal_1112}), .c ({signal_2158, signal_1048}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_284 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({signal_1868, signal_1113}), .c ({signal_1912, signal_1049}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_285 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({signal_1972, signal_1114}), .c ({signal_2160, signal_1050}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_286 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({signal_1969, signal_1115}), .c ({signal_2162, signal_1051}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_287 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({signal_1921, signal_1134}), .c ({signal_2164, signal_1070}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_288 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({signal_1865, signal_1116}), .c ({signal_1914, signal_1052}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_289 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({signal_1966, signal_1117}), .c ({signal_2166, signal_1053}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_290 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({signal_1963, signal_1118}), .c ({signal_2168, signal_1054}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_291 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({signal_1862, signal_1119}), .c ({signal_1916, signal_1055}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_292 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({signal_1960, signal_1120}), .c ({signal_2170, signal_1056}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_293 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({signal_1957, signal_1121}), .c ({signal_2172, signal_1057}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_294 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({signal_1954, signal_1122}), .c ({signal_2174, signal_1058}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_295 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({signal_1951, signal_1123}), .c ({signal_2176, signal_1059}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_296 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({signal_1948, signal_1124}), .c ({signal_2178, signal_1060}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_297 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({signal_1945, signal_1125}), .c ({signal_2180, signal_1061}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_298 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({signal_1856, signal_1135}), .c ({signal_1918, signal_1071}) ) ;
    INV_X1 cell_299 ( .A (signal_349), .ZN (signal_351) ) ;
    INV_X1 cell_300 ( .A (signal_311), .ZN (signal_349) ) ;
    INV_X1 cell_301 ( .A (signal_349), .ZN (signal_350) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_302 ( .s (signal_311), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({signal_1918, signal_1071}), .c ({signal_2072, signal_312}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_303 ( .s (signal_311), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({signal_2164, signal_1070}), .c ({signal_2192, signal_313}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_304 ( .s (signal_311), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({signal_2150, signal_1069}), .c ({signal_2193, signal_314}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_305 ( .s (signal_311), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({signal_1894, signal_1068}), .c ({signal_2073, signal_315}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_306 ( .s (signal_350), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({signal_2118, signal_1067}), .c ({signal_2194, signal_316}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_307 ( .s (signal_350), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({signal_2096, signal_1066}), .c ({signal_2195, signal_317}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_308 ( .s (signal_350), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({signal_2086, signal_1065}), .c ({signal_2196, signal_318}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_309 ( .s (signal_350), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({signal_2084, signal_1064}), .c ({signal_2197, signal_1000}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_310 ( .s (signal_350), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({signal_2082, signal_1063}), .c ({signal_2198, signal_999}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_311 ( .s (signal_350), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({signal_2080, signal_1062}), .c ({signal_2199, signal_998}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_312 ( .s (signal_350), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({signal_2180, signal_1061}), .c ({signal_2200, signal_997}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_313 ( .s (signal_350), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({signal_2178, signal_1060}), .c ({signal_2201, signal_996}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_314 ( .s (signal_350), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({signal_2176, signal_1059}), .c ({signal_2202, signal_995}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_315 ( .s (signal_350), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({signal_2174, signal_1058}), .c ({signal_2203, signal_994}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_316 ( .s (signal_350), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({signal_2172, signal_1057}), .c ({signal_2204, signal_993}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_317 ( .s (signal_350), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({signal_2170, signal_1056}), .c ({signal_2205, signal_992}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_318 ( .s (signal_311), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({signal_1916, signal_1055}), .c ({signal_2074, signal_319}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_319 ( .s (signal_311), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({signal_2168, signal_1054}), .c ({signal_2206, signal_320}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_320 ( .s (signal_311), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({signal_2166, signal_1053}), .c ({signal_2207, signal_321}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_321 ( .s (signal_311), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({signal_1914, signal_1052}), .c ({signal_2075, signal_322}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_322 ( .s (signal_350), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({signal_2162, signal_1051}), .c ({signal_2208, signal_323}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_323 ( .s (signal_311), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({signal_2160, signal_1050}), .c ({signal_2209, signal_324}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_324 ( .s (signal_311), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({signal_1912, signal_1049}), .c ({signal_2076, signal_325}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_325 ( .s (signal_311), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({signal_2158, signal_1048}), .c ({signal_2210, signal_984}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_326 ( .s (signal_311), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({signal_1910, signal_1047}), .c ({signal_2077, signal_983}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_327 ( .s (signal_311), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({signal_2156, signal_1046}), .c ({signal_2211, signal_982}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_328 ( .s (signal_311), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({signal_1908, signal_1045}), .c ({signal_2078, signal_981}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_329 ( .s (signal_311), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({signal_2154, signal_1044}), .c ({signal_2212, signal_980}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_330 ( .s (signal_351), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({signal_1906, signal_1043}), .c ({signal_2181, signal_979}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_331 ( .s (signal_351), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({signal_2152, signal_1042}), .c ({signal_2213, signal_978}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_332 ( .s (signal_351), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({signal_2148, signal_1041}), .c ({signal_2214, signal_977}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_333 ( .s (signal_351), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({signal_2146, signal_1040}), .c ({signal_2215, signal_976}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_334 ( .s (signal_351), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({signal_1904, signal_1039}), .c ({signal_2182, signal_326}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_335 ( .s (signal_351), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({signal_2144, signal_1038}), .c ({signal_2216, signal_327}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_336 ( .s (signal_351), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({signal_1902, signal_1037}), .c ({signal_2183, signal_328}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_337 ( .s (signal_351), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({signal_1900, signal_1036}), .c ({signal_2184, signal_329}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_338 ( .s (signal_351), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({signal_1898, signal_1035}), .c ({signal_2185, signal_330}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_339 ( .s (signal_311), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({signal_2142, signal_1034}), .c ({signal_2217, signal_331}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_340 ( .s (signal_351), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({signal_2140, signal_1033}), .c ({signal_2218, signal_332}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_341 ( .s (signal_351), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({signal_1896, signal_1032}), .c ({signal_2186, signal_968}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_342 ( .s (signal_351), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({signal_2138, signal_1031}), .c ({signal_2219, signal_967}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_343 ( .s (signal_351), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({signal_2136, signal_1030}), .c ({signal_2220, signal_966}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_344 ( .s (signal_351), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({signal_2134, signal_1029}), .c ({signal_2221, signal_965}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_345 ( .s (signal_351), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({signal_2132, signal_1028}), .c ({signal_2222, signal_964}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_346 ( .s (signal_351), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({signal_2130, signal_1027}), .c ({signal_2223, signal_963}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_347 ( .s (signal_351), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({signal_2128, signal_1026}), .c ({signal_2224, signal_962}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_348 ( .s (signal_351), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({signal_2126, signal_1025}), .c ({signal_2225, signal_961}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_349 ( .s (signal_351), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({signal_2124, signal_1024}), .c ({signal_2226, signal_960}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_350 ( .s (signal_351), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({signal_2122, signal_1023}), .c ({signal_2227, signal_333}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_351 ( .s (signal_351), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({signal_2120, signal_1022}), .c ({signal_2228, signal_334}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_352 ( .s (signal_311), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({signal_2116, signal_1021}), .c ({signal_2229, signal_335}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_353 ( .s (signal_351), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({signal_2114, signal_1020}), .c ({signal_2230, signal_336}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_354 ( .s (signal_351), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({signal_2112, signal_1019}), .c ({signal_2231, signal_337}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_355 ( .s (signal_351), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({signal_2110, signal_1018}), .c ({signal_2232, signal_338}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_356 ( .s (signal_351), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({signal_2108, signal_1017}), .c ({signal_2233, signal_339}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_357 ( .s (signal_351), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({signal_2106, signal_1016}), .c ({signal_2234, signal_952}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_358 ( .s (signal_351), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({signal_2104, signal_1015}), .c ({signal_2235, signal_951}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_359 ( .s (signal_351), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({signal_2102, signal_1014}), .c ({signal_2236, signal_950}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_360 ( .s (signal_351), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({signal_2100, signal_1013}), .c ({signal_2237, signal_949}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_361 ( .s (signal_351), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({signal_2098, signal_1012}), .c ({signal_2238, signal_948}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_362 ( .s (signal_351), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({signal_2094, signal_1011}), .c ({signal_2239, signal_947}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_363 ( .s (signal_351), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({signal_2092, signal_1010}), .c ({signal_2240, signal_946}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_364 ( .s (signal_351), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({signal_2090, signal_1009}), .c ({signal_2241, signal_945}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_365 ( .s (signal_351), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({signal_2088, signal_1008}), .c ({signal_2242, signal_944}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_366 ( .a ({1'b0, signal_874}), .b ({signal_2196, signal_318}), .c ({signal_2247, signal_1001}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_367 ( .a ({1'b0, signal_875}), .b ({signal_2195, signal_317}), .c ({signal_2248, signal_1002}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_368 ( .a ({1'b0, signal_877}), .b ({signal_2233, signal_339}), .c ({signal_2249, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_369 ( .a ({1'b0, signal_878}), .b ({signal_2232, signal_338}), .c ({signal_2250, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_370 ( .a ({1'b0, signal_879}), .b ({signal_2231, signal_337}), .c ({signal_2251, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_371 ( .a ({1'b0, 1'b0}), .b ({signal_2230, signal_336}), .c ({signal_2252, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_372 ( .a ({1'b0, 1'b0}), .b ({signal_2229, signal_335}), .c ({signal_2253, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_373 ( .a ({1'b0, signal_876}), .b ({signal_2194, signal_316}), .c ({signal_2254, signal_1003}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_374 ( .a ({1'b0, 1'b0}), .b ({signal_2228, signal_334}), .c ({signal_2255, signal_958}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_375 ( .a ({1'b0, 1'b0}), .b ({signal_2227, signal_333}), .c ({signal_2256, signal_959}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_2073, signal_315}), .c ({signal_2187, signal_1004}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_377 ( .a ({1'b0, signal_874}), .b ({signal_2218, signal_332}), .c ({signal_2257, signal_969}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_378 ( .a ({1'b0, signal_875}), .b ({signal_2217, signal_331}), .c ({signal_2258, signal_970}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_379 ( .a ({1'b0, signal_876}), .b ({signal_2185, signal_330}), .c ({signal_2243, signal_971}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_380 ( .a ({1'b0, 1'b0}), .b ({signal_2184, signal_329}), .c ({signal_2244, signal_972}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_381 ( .a ({1'b0, 1'b0}), .b ({signal_2183, signal_328}), .c ({signal_2245, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_382 ( .a ({1'b0, 1'b0}), .b ({signal_2216, signal_327}), .c ({signal_2259, signal_974}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_383 ( .a ({1'b0, 1'b0}), .b ({signal_2182, signal_326}), .c ({signal_2246, signal_975}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_384 ( .a ({1'b0, 1'b0}), .b ({signal_2193, signal_314}), .c ({signal_2260, signal_1005}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_385 ( .a ({1'b0, signal_877}), .b ({signal_2076, signal_325}), .c ({signal_2188, signal_985}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_386 ( .a ({1'b0, signal_878}), .b ({signal_2209, signal_324}), .c ({signal_2261, signal_986}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_387 ( .a ({1'b0, signal_879}), .b ({signal_2208, signal_323}), .c ({signal_2262, signal_987}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_388 ( .a ({1'b0, 1'b0}), .b ({signal_2192, signal_313}), .c ({signal_2263, signal_1006}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_389 ( .a ({1'b0, 1'b1}), .b ({signal_2075, signal_322}), .c ({signal_2189, signal_988}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_390 ( .a ({1'b0, 1'b0}), .b ({signal_2207, signal_321}), .c ({signal_2264, signal_989}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_391 ( .a ({1'b0, 1'b0}), .b ({signal_2206, signal_320}), .c ({signal_2265, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_392 ( .a ({1'b0, 1'b0}), .b ({signal_2074, signal_319}), .c ({signal_2190, signal_991}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_393 ( .a ({1'b0, 1'b0}), .b ({signal_2072, signal_312}), .c ({signal_2191, signal_1007}) ) ;
    INV_X1 cell_978 ( .A (signal_808), .ZN (signal_309) ) ;
    INV_X1 cell_980 ( .A (signal_307), .ZN (signal_306) ) ;
    INV_X1 cell_982 ( .A (signal_304), .ZN (signal_289) ) ;
    INV_X1 cell_984 ( .A (signal_288), .ZN (signal_302) ) ;
    INV_X1 cell_986 ( .A (signal_879), .ZN (signal_300) ) ;
    INV_X1 cell_988 ( .A (signal_878), .ZN (signal_298) ) ;
    INV_X1 cell_990 ( .A (signal_877), .ZN (signal_296) ) ;
    INV_X1 cell_992 ( .A (signal_876), .ZN (signal_294) ) ;
    INV_X1 cell_994 ( .A (signal_875), .ZN (signal_292) ) ;
    INV_X1 cell_996 ( .A (signal_874), .ZN (signal_290) ) ;

    /* cells in depth 1 */
    buf_clk cell_1726 ( .C (CLK), .D (signal_997), .Q (signal_3870) ) ;
    buf_clk cell_1728 ( .C (CLK), .D (signal_2200), .Q (signal_3872) ) ;
    buf_clk cell_1730 ( .C (CLK), .D (signal_993), .Q (signal_3874) ) ;
    buf_clk cell_1732 ( .C (CLK), .D (signal_2204), .Q (signal_3876) ) ;
    buf_clk cell_1734 ( .C (CLK), .D (signal_982), .Q (signal_3878) ) ;
    buf_clk cell_1736 ( .C (CLK), .D (signal_2211), .Q (signal_3880) ) ;
    buf_clk cell_1738 ( .C (CLK), .D (signal_977), .Q (signal_3882) ) ;
    buf_clk cell_1740 ( .C (CLK), .D (signal_2214), .Q (signal_3884) ) ;
    buf_clk cell_1742 ( .C (CLK), .D (signal_965), .Q (signal_3886) ) ;
    buf_clk cell_1744 ( .C (CLK), .D (signal_2221), .Q (signal_3888) ) ;
    buf_clk cell_1746 ( .C (CLK), .D (signal_961), .Q (signal_3890) ) ;
    buf_clk cell_1748 ( .C (CLK), .D (signal_2225), .Q (signal_3892) ) ;
    buf_clk cell_1750 ( .C (CLK), .D (signal_949), .Q (signal_3894) ) ;
    buf_clk cell_1752 ( .C (CLK), .D (signal_2237), .Q (signal_3896) ) ;
    buf_clk cell_1754 ( .C (CLK), .D (signal_945), .Q (signal_3898) ) ;
    buf_clk cell_1756 ( .C (CLK), .D (signal_2241), .Q (signal_3900) ) ;
    buf_clk cell_1758 ( .C (CLK), .D (signal_1005), .Q (signal_3902) ) ;
    buf_clk cell_1760 ( .C (CLK), .D (signal_2260), .Q (signal_3904) ) ;
    buf_clk cell_1762 ( .C (CLK), .D (signal_1002), .Q (signal_3906) ) ;
    buf_clk cell_1764 ( .C (CLK), .D (signal_2248), .Q (signal_3908) ) ;
    buf_clk cell_1766 ( .C (CLK), .D (signal_989), .Q (signal_3910) ) ;
    buf_clk cell_1768 ( .C (CLK), .D (signal_2264), .Q (signal_3912) ) ;
    buf_clk cell_1770 ( .C (CLK), .D (signal_986), .Q (signal_3914) ) ;
    buf_clk cell_1772 ( .C (CLK), .D (signal_2261), .Q (signal_3916) ) ;
    buf_clk cell_1774 ( .C (CLK), .D (signal_975), .Q (signal_3918) ) ;
    buf_clk cell_1776 ( .C (CLK), .D (signal_2246), .Q (signal_3920) ) ;
    buf_clk cell_1778 ( .C (CLK), .D (signal_969), .Q (signal_3922) ) ;
    buf_clk cell_1780 ( .C (CLK), .D (signal_2257), .Q (signal_3924) ) ;
    buf_clk cell_1782 ( .C (CLK), .D (signal_958), .Q (signal_3926) ) ;
    buf_clk cell_1784 ( .C (CLK), .D (signal_2255), .Q (signal_3928) ) ;
    buf_clk cell_1786 ( .C (CLK), .D (signal_954), .Q (signal_3930) ) ;
    buf_clk cell_1788 ( .C (CLK), .D (signal_2250), .Q (signal_3932) ) ;
    buf_clk cell_1790 ( .C (CLK), .D (signal_964), .Q (signal_3934) ) ;
    buf_clk cell_1792 ( .C (CLK), .D (signal_2222), .Q (signal_3936) ) ;
    buf_clk cell_1794 ( .C (CLK), .D (signal_987), .Q (signal_3938) ) ;
    buf_clk cell_1796 ( .C (CLK), .D (signal_2262), .Q (signal_3940) ) ;
    buf_clk cell_1798 ( .C (CLK), .D (signal_970), .Q (signal_3942) ) ;
    buf_clk cell_1800 ( .C (CLK), .D (signal_2258), .Q (signal_3944) ) ;
    buf_clk cell_1802 ( .C (CLK), .D (signal_1003), .Q (signal_3946) ) ;
    buf_clk cell_1804 ( .C (CLK), .D (signal_2254), .Q (signal_3948) ) ;
    buf_clk cell_1806 ( .C (CLK), .D (signal_984), .Q (signal_3950) ) ;
    buf_clk cell_1808 ( .C (CLK), .D (signal_2210), .Q (signal_3952) ) ;
    buf_clk cell_1810 ( .C (CLK), .D (signal_998), .Q (signal_3954) ) ;
    buf_clk cell_1814 ( .C (CLK), .D (signal_2199), .Q (signal_3958) ) ;
    buf_clk cell_1822 ( .C (CLK), .D (signal_994), .Q (signal_3966) ) ;
    buf_clk cell_1826 ( .C (CLK), .D (signal_2203), .Q (signal_3970) ) ;
    buf_clk cell_1834 ( .C (CLK), .D (signal_981), .Q (signal_3978) ) ;
    buf_clk cell_1838 ( .C (CLK), .D (signal_2078), .Q (signal_3982) ) ;
    buf_clk cell_1846 ( .C (CLK), .D (signal_978), .Q (signal_3990) ) ;
    buf_clk cell_1850 ( .C (CLK), .D (signal_2213), .Q (signal_3994) ) ;
    buf_clk cell_1858 ( .C (CLK), .D (signal_966), .Q (signal_4002) ) ;
    buf_clk cell_1862 ( .C (CLK), .D (signal_2220), .Q (signal_4006) ) ;
    buf_clk cell_1870 ( .C (CLK), .D (signal_962), .Q (signal_4014) ) ;
    buf_clk cell_1874 ( .C (CLK), .D (signal_2224), .Q (signal_4018) ) ;
    buf_clk cell_1882 ( .C (CLK), .D (signal_950), .Q (signal_4026) ) ;
    buf_clk cell_1886 ( .C (CLK), .D (signal_2236), .Q (signal_4030) ) ;
    buf_clk cell_1894 ( .C (CLK), .D (signal_946), .Q (signal_4038) ) ;
    buf_clk cell_1898 ( .C (CLK), .D (signal_2240), .Q (signal_4042) ) ;
    buf_clk cell_1906 ( .C (CLK), .D (signal_1007), .Q (signal_4050) ) ;
    buf_clk cell_1910 ( .C (CLK), .D (signal_2191), .Q (signal_4054) ) ;
    buf_clk cell_1922 ( .C (CLK), .D (signal_1001), .Q (signal_4066) ) ;
    buf_clk cell_1926 ( .C (CLK), .D (signal_2247), .Q (signal_4070) ) ;
    buf_clk cell_1938 ( .C (CLK), .D (signal_991), .Q (signal_4082) ) ;
    buf_clk cell_1942 ( .C (CLK), .D (signal_2190), .Q (signal_4086) ) ;
    buf_clk cell_1966 ( .C (CLK), .D (signal_973), .Q (signal_4110) ) ;
    buf_clk cell_1970 ( .C (CLK), .D (signal_2245), .Q (signal_4114) ) ;
    buf_clk cell_1982 ( .C (CLK), .D (signal_971), .Q (signal_4126) ) ;
    buf_clk cell_1986 ( .C (CLK), .D (signal_2243), .Q (signal_4130) ) ;
    buf_clk cell_1998 ( .C (CLK), .D (signal_957), .Q (signal_4142) ) ;
    buf_clk cell_2002 ( .C (CLK), .D (signal_2253), .Q (signal_4146) ) ;
    buf_clk cell_2014 ( .C (CLK), .D (signal_953), .Q (signal_4158) ) ;
    buf_clk cell_2018 ( .C (CLK), .D (signal_2249), .Q (signal_4162) ) ;
    buf_clk cell_2158 ( .C (CLK), .D (signal_944), .Q (signal_4302) ) ;
    buf_clk cell_2162 ( .C (CLK), .D (signal_2242), .Q (signal_4306) ) ;
    buf_clk cell_2174 ( .C (CLK), .D (signal_992), .Q (signal_4318) ) ;
    buf_clk cell_2178 ( .C (CLK), .D (signal_2205), .Q (signal_4322) ) ;
    buf_clk cell_2190 ( .C (CLK), .D (signal_343), .Q (signal_4334) ) ;
    buf_clk cell_2198 ( .C (CLK), .D (signal_313), .Q (signal_4342) ) ;
    buf_clk cell_2206 ( .C (CLK), .D (signal_2192), .Q (signal_4350) ) ;
    buf_clk cell_2214 ( .C (CLK), .D (signal_342), .Q (signal_4358) ) ;
    buf_clk cell_2222 ( .C (CLK), .D (signal_315), .Q (signal_4366) ) ;
    buf_clk cell_2230 ( .C (CLK), .D (signal_2073), .Q (signal_4374) ) ;
    buf_clk cell_2238 ( .C (CLK), .D (signal_317), .Q (signal_4382) ) ;
    buf_clk cell_2246 ( .C (CLK), .D (signal_2195), .Q (signal_4390) ) ;
    buf_clk cell_2254 ( .C (CLK), .D (signal_1000), .Q (signal_4398) ) ;
    buf_clk cell_2262 ( .C (CLK), .D (signal_2197), .Q (signal_4406) ) ;
    buf_clk cell_2278 ( .C (CLK), .D (signal_996), .Q (signal_4422) ) ;
    buf_clk cell_2286 ( .C (CLK), .D (signal_2201), .Q (signal_4430) ) ;
    buf_clk cell_2310 ( .C (CLK), .D (signal_321), .Q (signal_4454) ) ;
    buf_clk cell_2318 ( .C (CLK), .D (signal_2207), .Q (signal_4462) ) ;
    buf_clk cell_2326 ( .C (CLK), .D (signal_325), .Q (signal_4470) ) ;
    buf_clk cell_2334 ( .C (CLK), .D (signal_2076), .Q (signal_4478) ) ;
    buf_clk cell_2350 ( .C (CLK), .D (signal_344), .Q (signal_4494) ) ;
    buf_clk cell_2370 ( .C (CLK), .D (IN_reset), .Q (signal_4514) ) ;
    buf_clk cell_2378 ( .C (CLK), .D (IN_plaintext_s0[1]), .Q (signal_4522) ) ;
    buf_clk cell_2386 ( .C (CLK), .D (IN_plaintext_s1[1]), .Q (signal_4530) ) ;
    buf_clk cell_2394 ( .C (CLK), .D (IN_plaintext_s0[3]), .Q (signal_4538) ) ;
    buf_clk cell_2402 ( .C (CLK), .D (IN_plaintext_s1[3]), .Q (signal_4546) ) ;
    buf_clk cell_2410 ( .C (CLK), .D (IN_plaintext_s0[5]), .Q (signal_4554) ) ;
    buf_clk cell_2418 ( .C (CLK), .D (IN_plaintext_s1[5]), .Q (signal_4562) ) ;
    buf_clk cell_2426 ( .C (CLK), .D (IN_plaintext_s0[7]), .Q (signal_4570) ) ;
    buf_clk cell_2434 ( .C (CLK), .D (IN_plaintext_s1[7]), .Q (signal_4578) ) ;
    buf_clk cell_2442 ( .C (CLK), .D (IN_plaintext_s0[9]), .Q (signal_4586) ) ;
    buf_clk cell_2450 ( .C (CLK), .D (IN_plaintext_s1[9]), .Q (signal_4594) ) ;
    buf_clk cell_2458 ( .C (CLK), .D (IN_plaintext_s0[11]), .Q (signal_4602) ) ;
    buf_clk cell_2466 ( .C (CLK), .D (IN_plaintext_s1[11]), .Q (signal_4610) ) ;
    buf_clk cell_2474 ( .C (CLK), .D (IN_plaintext_s0[13]), .Q (signal_4618) ) ;
    buf_clk cell_2482 ( .C (CLK), .D (IN_plaintext_s1[13]), .Q (signal_4626) ) ;
    buf_clk cell_2490 ( .C (CLK), .D (IN_plaintext_s0[15]), .Q (signal_4634) ) ;
    buf_clk cell_2498 ( .C (CLK), .D (IN_plaintext_s1[15]), .Q (signal_4642) ) ;
    buf_clk cell_2506 ( .C (CLK), .D (IN_plaintext_s0[18]), .Q (signal_4650) ) ;
    buf_clk cell_2514 ( .C (CLK), .D (IN_plaintext_s1[18]), .Q (signal_4658) ) ;
    buf_clk cell_2522 ( .C (CLK), .D (IN_plaintext_s0[22]), .Q (signal_4666) ) ;
    buf_clk cell_2530 ( .C (CLK), .D (IN_plaintext_s1[22]), .Q (signal_4674) ) ;
    buf_clk cell_2538 ( .C (CLK), .D (IN_plaintext_s0[26]), .Q (signal_4682) ) ;
    buf_clk cell_2546 ( .C (CLK), .D (IN_plaintext_s1[26]), .Q (signal_4690) ) ;
    buf_clk cell_2554 ( .C (CLK), .D (IN_plaintext_s0[30]), .Q (signal_4698) ) ;
    buf_clk cell_2562 ( .C (CLK), .D (IN_plaintext_s1[30]), .Q (signal_4706) ) ;
    buf_clk cell_2586 ( .C (CLK), .D (signal_999), .Q (signal_4730) ) ;
    buf_clk cell_2594 ( .C (CLK), .D (signal_2198), .Q (signal_4738) ) ;
    buf_clk cell_2602 ( .C (CLK), .D (signal_995), .Q (signal_4746) ) ;
    buf_clk cell_2610 ( .C (CLK), .D (signal_2202), .Q (signal_4754) ) ;
    buf_clk cell_2638 ( .C (CLK), .D (signal_983), .Q (signal_4782) ) ;
    buf_clk cell_2646 ( .C (CLK), .D (signal_2077), .Q (signal_4790) ) ;
    buf_clk cell_2654 ( .C (CLK), .D (signal_979), .Q (signal_4798) ) ;
    buf_clk cell_2662 ( .C (CLK), .D (signal_2181), .Q (signal_4806) ) ;
    buf_clk cell_2690 ( .C (CLK), .D (signal_967), .Q (signal_4834) ) ;
    buf_clk cell_2698 ( .C (CLK), .D (signal_2219), .Q (signal_4842) ) ;
    buf_clk cell_2706 ( .C (CLK), .D (signal_963), .Q (signal_4850) ) ;
    buf_clk cell_2714 ( .C (CLK), .D (signal_2223), .Q (signal_4858) ) ;
    buf_clk cell_2722 ( .C (CLK), .D (signal_959), .Q (signal_4866) ) ;
    buf_clk cell_2730 ( .C (CLK), .D (signal_2256), .Q (signal_4874) ) ;
    buf_clk cell_2738 ( .C (CLK), .D (signal_955), .Q (signal_4882) ) ;
    buf_clk cell_2746 ( .C (CLK), .D (signal_2251), .Q (signal_4890) ) ;
    buf_clk cell_2754 ( .C (CLK), .D (signal_951), .Q (signal_4898) ) ;
    buf_clk cell_2762 ( .C (CLK), .D (signal_2235), .Q (signal_4906) ) ;
    buf_clk cell_2770 ( .C (CLK), .D (signal_947), .Q (signal_4914) ) ;
    buf_clk cell_2778 ( .C (CLK), .D (signal_2239), .Q (signal_4922) ) ;
    buf_clk cell_2786 ( .C (CLK), .D (signal_1004), .Q (signal_4930) ) ;
    buf_clk cell_2792 ( .C (CLK), .D (signal_2187), .Q (signal_4936) ) ;
    buf_clk cell_2798 ( .C (CLK), .D (signal_988), .Q (signal_4942) ) ;
    buf_clk cell_2804 ( .C (CLK), .D (signal_2189), .Q (signal_4948) ) ;
    buf_clk cell_2810 ( .C (CLK), .D (signal_985), .Q (signal_4954) ) ;
    buf_clk cell_2816 ( .C (CLK), .D (signal_2188), .Q (signal_4960) ) ;
    buf_clk cell_2822 ( .C (CLK), .D (signal_972), .Q (signal_4966) ) ;
    buf_clk cell_2828 ( .C (CLK), .D (signal_2244), .Q (signal_4972) ) ;
    buf_clk cell_2834 ( .C (CLK), .D (signal_968), .Q (signal_4978) ) ;
    buf_clk cell_2840 ( .C (CLK), .D (signal_2186), .Q (signal_4984) ) ;
    buf_clk cell_2846 ( .C (CLK), .D (signal_956), .Q (signal_4990) ) ;
    buf_clk cell_2852 ( .C (CLK), .D (signal_2252), .Q (signal_4996) ) ;
    buf_clk cell_2858 ( .C (CLK), .D (signal_952), .Q (signal_5002) ) ;
    buf_clk cell_2864 ( .C (CLK), .D (signal_2234), .Q (signal_5008) ) ;
    buf_clk cell_2970 ( .C (CLK), .D (signal_980), .Q (signal_5114) ) ;
    buf_clk cell_2976 ( .C (CLK), .D (signal_2212), .Q (signal_5120) ) ;
    buf_clk cell_3054 ( .C (CLK), .D (signal_976), .Q (signal_5198) ) ;
    buf_clk cell_3062 ( .C (CLK), .D (signal_2215), .Q (signal_5206) ) ;
    buf_clk cell_3446 ( .C (CLK), .D (signal_312), .Q (signal_5590) ) ;
    buf_clk cell_3462 ( .C (CLK), .D (signal_2072), .Q (signal_5606) ) ;
    buf_clk cell_3486 ( .C (CLK), .D (signal_314), .Q (signal_5630) ) ;
    buf_clk cell_3502 ( .C (CLK), .D (signal_2193), .Q (signal_5646) ) ;
    buf_clk cell_3526 ( .C (CLK), .D (signal_316), .Q (signal_5670) ) ;
    buf_clk cell_3542 ( .C (CLK), .D (signal_2194), .Q (signal_5686) ) ;
    buf_clk cell_3558 ( .C (CLK), .D (signal_318), .Q (signal_5702) ) ;
    buf_clk cell_3574 ( .C (CLK), .D (signal_2196), .Q (signal_5718) ) ;
    buf_clk cell_3634 ( .C (CLK), .D (signal_319), .Q (signal_5778) ) ;
    buf_clk cell_3650 ( .C (CLK), .D (signal_2074), .Q (signal_5794) ) ;
    buf_clk cell_3666 ( .C (CLK), .D (signal_320), .Q (signal_5810) ) ;
    buf_clk cell_3682 ( .C (CLK), .D (signal_2206), .Q (signal_5826) ) ;
    buf_clk cell_3698 ( .C (CLK), .D (signal_322), .Q (signal_5842) ) ;
    buf_clk cell_3714 ( .C (CLK), .D (signal_2075), .Q (signal_5858) ) ;
    buf_clk cell_3730 ( .C (CLK), .D (signal_323), .Q (signal_5874) ) ;
    buf_clk cell_3746 ( .C (CLK), .D (signal_2208), .Q (signal_5890) ) ;
    buf_clk cell_3762 ( .C (CLK), .D (signal_324), .Q (signal_5906) ) ;
    buf_clk cell_3778 ( .C (CLK), .D (signal_2209), .Q (signal_5922) ) ;
    buf_clk cell_3886 ( .C (CLK), .D (signal_326), .Q (signal_6030) ) ;
    buf_clk cell_3902 ( .C (CLK), .D (signal_2182), .Q (signal_6046) ) ;
    buf_clk cell_3918 ( .C (CLK), .D (signal_327), .Q (signal_6062) ) ;
    buf_clk cell_3934 ( .C (CLK), .D (signal_2216), .Q (signal_6078) ) ;
    buf_clk cell_3950 ( .C (CLK), .D (signal_328), .Q (signal_6094) ) ;
    buf_clk cell_3966 ( .C (CLK), .D (signal_2183), .Q (signal_6110) ) ;
    buf_clk cell_3982 ( .C (CLK), .D (signal_329), .Q (signal_6126) ) ;
    buf_clk cell_3998 ( .C (CLK), .D (signal_2184), .Q (signal_6142) ) ;
    buf_clk cell_4014 ( .C (CLK), .D (signal_330), .Q (signal_6158) ) ;
    buf_clk cell_4030 ( .C (CLK), .D (signal_2185), .Q (signal_6174) ) ;
    buf_clk cell_4046 ( .C (CLK), .D (signal_331), .Q (signal_6190) ) ;
    buf_clk cell_4062 ( .C (CLK), .D (signal_2217), .Q (signal_6206) ) ;
    buf_clk cell_4078 ( .C (CLK), .D (signal_332), .Q (signal_6222) ) ;
    buf_clk cell_4094 ( .C (CLK), .D (signal_2218), .Q (signal_6238) ) ;
    buf_clk cell_4178 ( .C (CLK), .D (signal_340), .Q (signal_6322) ) ;
    buf_clk cell_4286 ( .C (CLK), .D (signal_960), .Q (signal_6430) ) ;
    buf_clk cell_4302 ( .C (CLK), .D (signal_2226), .Q (signal_6446) ) ;
    buf_clk cell_4318 ( .C (CLK), .D (signal_333), .Q (signal_6462) ) ;
    buf_clk cell_4334 ( .C (CLK), .D (signal_2227), .Q (signal_6478) ) ;
    buf_clk cell_4350 ( .C (CLK), .D (signal_334), .Q (signal_6494) ) ;
    buf_clk cell_4366 ( .C (CLK), .D (signal_2228), .Q (signal_6510) ) ;
    buf_clk cell_4382 ( .C (CLK), .D (signal_335), .Q (signal_6526) ) ;
    buf_clk cell_4398 ( .C (CLK), .D (signal_2229), .Q (signal_6542) ) ;
    buf_clk cell_4414 ( .C (CLK), .D (signal_336), .Q (signal_6558) ) ;
    buf_clk cell_4430 ( .C (CLK), .D (signal_2230), .Q (signal_6574) ) ;
    buf_clk cell_4446 ( .C (CLK), .D (signal_337), .Q (signal_6590) ) ;
    buf_clk cell_4462 ( .C (CLK), .D (signal_2231), .Q (signal_6606) ) ;
    buf_clk cell_4478 ( .C (CLK), .D (signal_338), .Q (signal_6622) ) ;
    buf_clk cell_4494 ( .C (CLK), .D (signal_2232), .Q (signal_6638) ) ;
    buf_clk cell_4510 ( .C (CLK), .D (signal_339), .Q (signal_6654) ) ;
    buf_clk cell_4526 ( .C (CLK), .D (signal_2233), .Q (signal_6670) ) ;
    buf_clk cell_4630 ( .C (CLK), .D (signal_948), .Q (signal_6774) ) ;
    buf_clk cell_4646 ( .C (CLK), .D (signal_2238), .Q (signal_6790) ) ;
    buf_clk cell_4742 ( .C (CLK), .D (IN_plaintext_s0[0]), .Q (signal_6886) ) ;
    buf_clk cell_4758 ( .C (CLK), .D (IN_plaintext_s1[0]), .Q (signal_6902) ) ;
    buf_clk cell_4774 ( .C (CLK), .D (IN_plaintext_s0[2]), .Q (signal_6918) ) ;
    buf_clk cell_4790 ( .C (CLK), .D (IN_plaintext_s1[2]), .Q (signal_6934) ) ;
    buf_clk cell_4806 ( .C (CLK), .D (IN_plaintext_s0[4]), .Q (signal_6950) ) ;
    buf_clk cell_4822 ( .C (CLK), .D (IN_plaintext_s1[4]), .Q (signal_6966) ) ;
    buf_clk cell_4838 ( .C (CLK), .D (IN_plaintext_s0[6]), .Q (signal_6982) ) ;
    buf_clk cell_4854 ( .C (CLK), .D (IN_plaintext_s1[6]), .Q (signal_6998) ) ;
    buf_clk cell_4870 ( .C (CLK), .D (IN_plaintext_s0[8]), .Q (signal_7014) ) ;
    buf_clk cell_4886 ( .C (CLK), .D (IN_plaintext_s1[8]), .Q (signal_7030) ) ;
    buf_clk cell_4902 ( .C (CLK), .D (IN_plaintext_s0[10]), .Q (signal_7046) ) ;
    buf_clk cell_4918 ( .C (CLK), .D (IN_plaintext_s1[10]), .Q (signal_7062) ) ;
    buf_clk cell_4934 ( .C (CLK), .D (IN_plaintext_s0[12]), .Q (signal_7078) ) ;
    buf_clk cell_4950 ( .C (CLK), .D (IN_plaintext_s1[12]), .Q (signal_7094) ) ;
    buf_clk cell_4966 ( .C (CLK), .D (IN_plaintext_s0[14]), .Q (signal_7110) ) ;
    buf_clk cell_4982 ( .C (CLK), .D (IN_plaintext_s1[14]), .Q (signal_7126) ) ;
    buf_clk cell_4998 ( .C (CLK), .D (IN_plaintext_s0[16]), .Q (signal_7142) ) ;
    buf_clk cell_5014 ( .C (CLK), .D (IN_plaintext_s1[16]), .Q (signal_7158) ) ;
    buf_clk cell_5030 ( .C (CLK), .D (IN_plaintext_s0[17]), .Q (signal_7174) ) ;
    buf_clk cell_5046 ( .C (CLK), .D (IN_plaintext_s1[17]), .Q (signal_7190) ) ;
    buf_clk cell_5062 ( .C (CLK), .D (IN_plaintext_s0[19]), .Q (signal_7206) ) ;
    buf_clk cell_5078 ( .C (CLK), .D (IN_plaintext_s1[19]), .Q (signal_7222) ) ;
    buf_clk cell_5094 ( .C (CLK), .D (IN_plaintext_s0[20]), .Q (signal_7238) ) ;
    buf_clk cell_5110 ( .C (CLK), .D (IN_plaintext_s1[20]), .Q (signal_7254) ) ;
    buf_clk cell_5126 ( .C (CLK), .D (IN_plaintext_s0[21]), .Q (signal_7270) ) ;
    buf_clk cell_5142 ( .C (CLK), .D (IN_plaintext_s1[21]), .Q (signal_7286) ) ;
    buf_clk cell_5158 ( .C (CLK), .D (IN_plaintext_s0[23]), .Q (signal_7302) ) ;
    buf_clk cell_5174 ( .C (CLK), .D (IN_plaintext_s1[23]), .Q (signal_7318) ) ;
    buf_clk cell_5190 ( .C (CLK), .D (IN_plaintext_s0[24]), .Q (signal_7334) ) ;
    buf_clk cell_5206 ( .C (CLK), .D (IN_plaintext_s1[24]), .Q (signal_7350) ) ;
    buf_clk cell_5222 ( .C (CLK), .D (IN_plaintext_s0[25]), .Q (signal_7366) ) ;
    buf_clk cell_5238 ( .C (CLK), .D (IN_plaintext_s1[25]), .Q (signal_7382) ) ;
    buf_clk cell_5254 ( .C (CLK), .D (IN_plaintext_s0[27]), .Q (signal_7398) ) ;
    buf_clk cell_5270 ( .C (CLK), .D (IN_plaintext_s1[27]), .Q (signal_7414) ) ;
    buf_clk cell_5286 ( .C (CLK), .D (IN_plaintext_s0[28]), .Q (signal_7430) ) ;
    buf_clk cell_5302 ( .C (CLK), .D (IN_plaintext_s1[28]), .Q (signal_7446) ) ;
    buf_clk cell_5318 ( .C (CLK), .D (IN_plaintext_s0[29]), .Q (signal_7462) ) ;
    buf_clk cell_5334 ( .C (CLK), .D (IN_plaintext_s1[29]), .Q (signal_7478) ) ;
    buf_clk cell_5350 ( .C (CLK), .D (IN_plaintext_s0[31]), .Q (signal_7494) ) ;
    buf_clk cell_5366 ( .C (CLK), .D (IN_plaintext_s1[31]), .Q (signal_7510) ) ;
    buf_clk cell_5382 ( .C (CLK), .D (IN_plaintext_s0[32]), .Q (signal_7526) ) ;
    buf_clk cell_5398 ( .C (CLK), .D (IN_plaintext_s1[32]), .Q (signal_7542) ) ;
    buf_clk cell_5414 ( .C (CLK), .D (IN_plaintext_s0[33]), .Q (signal_7558) ) ;
    buf_clk cell_5430 ( .C (CLK), .D (IN_plaintext_s1[33]), .Q (signal_7574) ) ;
    buf_clk cell_5446 ( .C (CLK), .D (IN_plaintext_s0[34]), .Q (signal_7590) ) ;
    buf_clk cell_5462 ( .C (CLK), .D (IN_plaintext_s1[34]), .Q (signal_7606) ) ;
    buf_clk cell_5478 ( .C (CLK), .D (IN_plaintext_s0[35]), .Q (signal_7622) ) ;
    buf_clk cell_5494 ( .C (CLK), .D (IN_plaintext_s1[35]), .Q (signal_7638) ) ;
    buf_clk cell_5510 ( .C (CLK), .D (IN_plaintext_s0[36]), .Q (signal_7654) ) ;
    buf_clk cell_5526 ( .C (CLK), .D (IN_plaintext_s1[36]), .Q (signal_7670) ) ;
    buf_clk cell_5542 ( .C (CLK), .D (IN_plaintext_s0[37]), .Q (signal_7686) ) ;
    buf_clk cell_5558 ( .C (CLK), .D (IN_plaintext_s1[37]), .Q (signal_7702) ) ;
    buf_clk cell_5574 ( .C (CLK), .D (IN_plaintext_s0[38]), .Q (signal_7718) ) ;
    buf_clk cell_5590 ( .C (CLK), .D (IN_plaintext_s1[38]), .Q (signal_7734) ) ;
    buf_clk cell_5606 ( .C (CLK), .D (IN_plaintext_s0[39]), .Q (signal_7750) ) ;
    buf_clk cell_5622 ( .C (CLK), .D (IN_plaintext_s1[39]), .Q (signal_7766) ) ;
    buf_clk cell_5638 ( .C (CLK), .D (IN_plaintext_s0[40]), .Q (signal_7782) ) ;
    buf_clk cell_5654 ( .C (CLK), .D (IN_plaintext_s1[40]), .Q (signal_7798) ) ;
    buf_clk cell_5670 ( .C (CLK), .D (IN_plaintext_s0[41]), .Q (signal_7814) ) ;
    buf_clk cell_5686 ( .C (CLK), .D (IN_plaintext_s1[41]), .Q (signal_7830) ) ;
    buf_clk cell_5702 ( .C (CLK), .D (IN_plaintext_s0[42]), .Q (signal_7846) ) ;
    buf_clk cell_5718 ( .C (CLK), .D (IN_plaintext_s1[42]), .Q (signal_7862) ) ;
    buf_clk cell_5734 ( .C (CLK), .D (IN_plaintext_s0[43]), .Q (signal_7878) ) ;
    buf_clk cell_5750 ( .C (CLK), .D (IN_plaintext_s1[43]), .Q (signal_7894) ) ;
    buf_clk cell_5766 ( .C (CLK), .D (IN_plaintext_s0[44]), .Q (signal_7910) ) ;
    buf_clk cell_5782 ( .C (CLK), .D (IN_plaintext_s1[44]), .Q (signal_7926) ) ;
    buf_clk cell_5798 ( .C (CLK), .D (IN_plaintext_s0[45]), .Q (signal_7942) ) ;
    buf_clk cell_5814 ( .C (CLK), .D (IN_plaintext_s1[45]), .Q (signal_7958) ) ;
    buf_clk cell_5830 ( .C (CLK), .D (IN_plaintext_s0[46]), .Q (signal_7974) ) ;
    buf_clk cell_5846 ( .C (CLK), .D (IN_plaintext_s1[46]), .Q (signal_7990) ) ;
    buf_clk cell_5862 ( .C (CLK), .D (IN_plaintext_s0[47]), .Q (signal_8006) ) ;
    buf_clk cell_5878 ( .C (CLK), .D (IN_plaintext_s1[47]), .Q (signal_8022) ) ;
    buf_clk cell_5894 ( .C (CLK), .D (IN_plaintext_s0[48]), .Q (signal_8038) ) ;
    buf_clk cell_5910 ( .C (CLK), .D (IN_plaintext_s1[48]), .Q (signal_8054) ) ;
    buf_clk cell_5926 ( .C (CLK), .D (IN_plaintext_s0[49]), .Q (signal_8070) ) ;
    buf_clk cell_5942 ( .C (CLK), .D (IN_plaintext_s1[49]), .Q (signal_8086) ) ;
    buf_clk cell_5958 ( .C (CLK), .D (IN_plaintext_s0[50]), .Q (signal_8102) ) ;
    buf_clk cell_5974 ( .C (CLK), .D (IN_plaintext_s1[50]), .Q (signal_8118) ) ;
    buf_clk cell_5990 ( .C (CLK), .D (IN_plaintext_s0[51]), .Q (signal_8134) ) ;
    buf_clk cell_6006 ( .C (CLK), .D (IN_plaintext_s1[51]), .Q (signal_8150) ) ;
    buf_clk cell_6022 ( .C (CLK), .D (IN_plaintext_s0[52]), .Q (signal_8166) ) ;
    buf_clk cell_6038 ( .C (CLK), .D (IN_plaintext_s1[52]), .Q (signal_8182) ) ;
    buf_clk cell_6054 ( .C (CLK), .D (IN_plaintext_s0[53]), .Q (signal_8198) ) ;
    buf_clk cell_6070 ( .C (CLK), .D (IN_plaintext_s1[53]), .Q (signal_8214) ) ;
    buf_clk cell_6086 ( .C (CLK), .D (IN_plaintext_s0[54]), .Q (signal_8230) ) ;
    buf_clk cell_6102 ( .C (CLK), .D (IN_plaintext_s1[54]), .Q (signal_8246) ) ;
    buf_clk cell_6118 ( .C (CLK), .D (IN_plaintext_s0[55]), .Q (signal_8262) ) ;
    buf_clk cell_6134 ( .C (CLK), .D (IN_plaintext_s1[55]), .Q (signal_8278) ) ;
    buf_clk cell_6150 ( .C (CLK), .D (IN_plaintext_s0[56]), .Q (signal_8294) ) ;
    buf_clk cell_6166 ( .C (CLK), .D (IN_plaintext_s1[56]), .Q (signal_8310) ) ;
    buf_clk cell_6182 ( .C (CLK), .D (IN_plaintext_s0[57]), .Q (signal_8326) ) ;
    buf_clk cell_6198 ( .C (CLK), .D (IN_plaintext_s1[57]), .Q (signal_8342) ) ;
    buf_clk cell_6214 ( .C (CLK), .D (IN_plaintext_s0[58]), .Q (signal_8358) ) ;
    buf_clk cell_6230 ( .C (CLK), .D (IN_plaintext_s1[58]), .Q (signal_8374) ) ;
    buf_clk cell_6246 ( .C (CLK), .D (IN_plaintext_s0[59]), .Q (signal_8390) ) ;
    buf_clk cell_6262 ( .C (CLK), .D (IN_plaintext_s1[59]), .Q (signal_8406) ) ;
    buf_clk cell_6278 ( .C (CLK), .D (IN_plaintext_s0[60]), .Q (signal_8422) ) ;
    buf_clk cell_6294 ( .C (CLK), .D (IN_plaintext_s1[60]), .Q (signal_8438) ) ;
    buf_clk cell_6310 ( .C (CLK), .D (IN_plaintext_s0[61]), .Q (signal_8454) ) ;
    buf_clk cell_6326 ( .C (CLK), .D (IN_plaintext_s1[61]), .Q (signal_8470) ) ;
    buf_clk cell_6342 ( .C (CLK), .D (IN_plaintext_s0[62]), .Q (signal_8486) ) ;
    buf_clk cell_6358 ( .C (CLK), .D (IN_plaintext_s1[62]), .Q (signal_8502) ) ;
    buf_clk cell_6374 ( .C (CLK), .D (IN_plaintext_s0[63]), .Q (signal_8518) ) ;
    buf_clk cell_6390 ( .C (CLK), .D (IN_plaintext_s1[63]), .Q (signal_8534) ) ;
    buf_clk cell_7590 ( .C (CLK), .D (signal_310), .Q (signal_9734) ) ;
    buf_clk cell_7606 ( .C (CLK), .D (signal_308), .Q (signal_9750) ) ;
    buf_clk cell_7622 ( .C (CLK), .D (signal_305), .Q (signal_9766) ) ;
    buf_clk cell_7638 ( .C (CLK), .D (signal_303), .Q (signal_9782) ) ;
    buf_clk cell_7654 ( .C (CLK), .D (signal_301), .Q (signal_9798) ) ;
    buf_clk cell_7670 ( .C (CLK), .D (signal_299), .Q (signal_9814) ) ;
    buf_clk cell_7686 ( .C (CLK), .D (signal_297), .Q (signal_9830) ) ;
    buf_clk cell_7702 ( .C (CLK), .D (signal_295), .Q (signal_9846) ) ;
    buf_clk cell_7718 ( .C (CLK), .D (signal_293), .Q (signal_9862) ) ;
    buf_clk cell_7734 ( .C (CLK), .D (signal_291), .Q (signal_9878) ) ;
    buf_clk cell_7942 ( .C (CLK), .D (signal_265), .Q (signal_10086) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1128 ( .s ({signal_2201, signal_996}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[0]), .c ({signal_2266, signal_1328}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1129 ( .s ({signal_2201, signal_996}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[1]), .c ({signal_2267, signal_1329}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1130 ( .s ({signal_2205, signal_992}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[2]), .c ({signal_2268, signal_1330}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1131 ( .s ({signal_2205, signal_992}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[3]), .c ({signal_2269, signal_1331}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1132 ( .s ({signal_2212, signal_980}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[4]), .c ({signal_2270, signal_1332}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1133 ( .s ({signal_2212, signal_980}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[5]), .c ({signal_2271, signal_1333}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1134 ( .s ({signal_2215, signal_976}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[6]), .c ({signal_2272, signal_1334}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1135 ( .s ({signal_2215, signal_976}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[7]), .c ({signal_2273, signal_1335}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1136 ( .s ({signal_2222, signal_964}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[8]), .c ({signal_2274, signal_1336}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1137 ( .s ({signal_2222, signal_964}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[9]), .c ({signal_2275, signal_1337}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1138 ( .s ({signal_2226, signal_960}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[10]), .c ({signal_2276, signal_1338}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1139 ( .s ({signal_2226, signal_960}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[11]), .c ({signal_2277, signal_1339}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1140 ( .s ({signal_2238, signal_948}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[12]), .c ({signal_2278, signal_1340}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1141 ( .s ({signal_2238, signal_948}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[13]), .c ({signal_2279, signal_1341}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1142 ( .s ({signal_2242, signal_944}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[14]), .c ({signal_2280, signal_1342}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1143 ( .s ({signal_2242, signal_944}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[15]), .c ({signal_2281, signal_1343}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1144 ( .s ({signal_2260, signal_1005}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[16]), .c ({signal_2290, signal_1344}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1145 ( .s ({signal_2263, signal_1006}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[17]), .c ({signal_2291, signal_1345}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1146 ( .s ({signal_2263, signal_1006}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[18]), .c ({signal_2292, signal_1346}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1147 ( .s ({signal_2254, signal_1003}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[19]), .c ({signal_2293, signal_1347}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1148 ( .s ({signal_2254, signal_1003}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[20]), .c ({signal_2294, signal_1348}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1149 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[21]), .c ({signal_2295, signal_1349}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1150 ( .s ({signal_2264, signal_989}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[22]), .c ({signal_2296, signal_1350}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1151 ( .s ({signal_2265, signal_990}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[23]), .c ({signal_2297, signal_1351}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1152 ( .s ({signal_2265, signal_990}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[24]), .c ({signal_2298, signal_1352}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1153 ( .s ({signal_2262, signal_987}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[25]), .c ({signal_2299, signal_1353}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1154 ( .s ({signal_2262, signal_987}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[26]), .c ({signal_2300, signal_1354}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1155 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[27]), .c ({signal_2301, signal_1355}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1156 ( .s ({signal_2246, signal_975}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[28]), .c ({signal_2282, signal_1356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1157 ( .s ({signal_2259, signal_974}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[29]), .c ({signal_2302, signal_1357}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1158 ( .s ({signal_2259, signal_974}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[30]), .c ({signal_2303, signal_1358}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1159 ( .s ({signal_2257, signal_969}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[31]), .c ({signal_2304, signal_1359}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1160 ( .s ({signal_2258, signal_970}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[32]), .c ({signal_2305, signal_1360}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1161 ( .s ({signal_2258, signal_970}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[33]), .c ({signal_2306, signal_1361}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1162 ( .s ({signal_2256, signal_959}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[34]), .c ({signal_2307, signal_1362}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1163 ( .s ({signal_2256, signal_959}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[35]), .c ({signal_2308, signal_1363}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1164 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[36]), .c ({signal_2309, signal_1364}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1165 ( .s ({signal_2251, signal_955}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[37]), .c ({signal_2310, signal_1365}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1166 ( .s ({signal_2251, signal_955}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[38]), .c ({signal_2311, signal_1366}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1167 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[39]), .c ({signal_2312, signal_1367}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1168 ( .s ({signal_2221, signal_965}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[40]), .c ({signal_2283, signal_1368}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1169 ( .s ({signal_2241, signal_945}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[41]), .c ({signal_2284, signal_1369}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1170 ( .s ({signal_2225, signal_961}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[42]), .c ({signal_2285, signal_1370}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1171 ( .s ({signal_2257, signal_969}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[43]), .c ({signal_2313, signal_1371}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1172 ( .s ({signal_2264, signal_989}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[44]), .c ({signal_2314, signal_1372}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1173 ( .s ({signal_2261, signal_986}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[45]), .c ({signal_2315, signal_1373}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1174 ( .s ({signal_2255, signal_958}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[46]), .c ({signal_2316, signal_1374}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1175 ( .s ({signal_2248, signal_1002}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[47]), .c ({signal_2317, signal_1375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1176 ( .s ({signal_2250, signal_954}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[48]), .c ({signal_2318, signal_1376}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1177 ( .s ({signal_2246, signal_975}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[49]), .c ({signal_2286, signal_1377}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1178 ( .s ({signal_2200, signal_997}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[50]), .c ({signal_2287, signal_1378}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1179 ( .s ({signal_2204, signal_993}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[51]), .c ({signal_2288, signal_1379}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1180 ( .s ({signal_2237, signal_949}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[52]), .c ({signal_2289, signal_1380}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1181 ( .s ({signal_2260, signal_1005}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[53]), .c ({signal_2319, signal_1381}) ) ;
    buf_clk cell_1727 ( .C (CLK), .D (signal_3870), .Q (signal_3871) ) ;
    buf_clk cell_1729 ( .C (CLK), .D (signal_3872), .Q (signal_3873) ) ;
    buf_clk cell_1731 ( .C (CLK), .D (signal_3874), .Q (signal_3875) ) ;
    buf_clk cell_1733 ( .C (CLK), .D (signal_3876), .Q (signal_3877) ) ;
    buf_clk cell_1735 ( .C (CLK), .D (signal_3878), .Q (signal_3879) ) ;
    buf_clk cell_1737 ( .C (CLK), .D (signal_3880), .Q (signal_3881) ) ;
    buf_clk cell_1739 ( .C (CLK), .D (signal_3882), .Q (signal_3883) ) ;
    buf_clk cell_1741 ( .C (CLK), .D (signal_3884), .Q (signal_3885) ) ;
    buf_clk cell_1743 ( .C (CLK), .D (signal_3886), .Q (signal_3887) ) ;
    buf_clk cell_1745 ( .C (CLK), .D (signal_3888), .Q (signal_3889) ) ;
    buf_clk cell_1747 ( .C (CLK), .D (signal_3890), .Q (signal_3891) ) ;
    buf_clk cell_1749 ( .C (CLK), .D (signal_3892), .Q (signal_3893) ) ;
    buf_clk cell_1751 ( .C (CLK), .D (signal_3894), .Q (signal_3895) ) ;
    buf_clk cell_1753 ( .C (CLK), .D (signal_3896), .Q (signal_3897) ) ;
    buf_clk cell_1755 ( .C (CLK), .D (signal_3898), .Q (signal_3899) ) ;
    buf_clk cell_1757 ( .C (CLK), .D (signal_3900), .Q (signal_3901) ) ;
    buf_clk cell_1759 ( .C (CLK), .D (signal_3902), .Q (signal_3903) ) ;
    buf_clk cell_1761 ( .C (CLK), .D (signal_3904), .Q (signal_3905) ) ;
    buf_clk cell_1763 ( .C (CLK), .D (signal_3906), .Q (signal_3907) ) ;
    buf_clk cell_1765 ( .C (CLK), .D (signal_3908), .Q (signal_3909) ) ;
    buf_clk cell_1767 ( .C (CLK), .D (signal_3910), .Q (signal_3911) ) ;
    buf_clk cell_1769 ( .C (CLK), .D (signal_3912), .Q (signal_3913) ) ;
    buf_clk cell_1771 ( .C (CLK), .D (signal_3914), .Q (signal_3915) ) ;
    buf_clk cell_1773 ( .C (CLK), .D (signal_3916), .Q (signal_3917) ) ;
    buf_clk cell_1775 ( .C (CLK), .D (signal_3918), .Q (signal_3919) ) ;
    buf_clk cell_1777 ( .C (CLK), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_1779 ( .C (CLK), .D (signal_3922), .Q (signal_3923) ) ;
    buf_clk cell_1781 ( .C (CLK), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_1783 ( .C (CLK), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_1785 ( .C (CLK), .D (signal_3928), .Q (signal_3929) ) ;
    buf_clk cell_1787 ( .C (CLK), .D (signal_3930), .Q (signal_3931) ) ;
    buf_clk cell_1789 ( .C (CLK), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_1791 ( .C (CLK), .D (signal_3934), .Q (signal_3935) ) ;
    buf_clk cell_1793 ( .C (CLK), .D (signal_3936), .Q (signal_3937) ) ;
    buf_clk cell_1795 ( .C (CLK), .D (signal_3938), .Q (signal_3939) ) ;
    buf_clk cell_1797 ( .C (CLK), .D (signal_3940), .Q (signal_3941) ) ;
    buf_clk cell_1799 ( .C (CLK), .D (signal_3942), .Q (signal_3943) ) ;
    buf_clk cell_1801 ( .C (CLK), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_1803 ( .C (CLK), .D (signal_3946), .Q (signal_3947) ) ;
    buf_clk cell_1805 ( .C (CLK), .D (signal_3948), .Q (signal_3949) ) ;
    buf_clk cell_1807 ( .C (CLK), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_1809 ( .C (CLK), .D (signal_3952), .Q (signal_3953) ) ;
    buf_clk cell_1811 ( .C (CLK), .D (signal_3954), .Q (signal_3955) ) ;
    buf_clk cell_1815 ( .C (CLK), .D (signal_3958), .Q (signal_3959) ) ;
    buf_clk cell_1823 ( .C (CLK), .D (signal_3966), .Q (signal_3967) ) ;
    buf_clk cell_1827 ( .C (CLK), .D (signal_3970), .Q (signal_3971) ) ;
    buf_clk cell_1835 ( .C (CLK), .D (signal_3978), .Q (signal_3979) ) ;
    buf_clk cell_1839 ( .C (CLK), .D (signal_3982), .Q (signal_3983) ) ;
    buf_clk cell_1847 ( .C (CLK), .D (signal_3990), .Q (signal_3991) ) ;
    buf_clk cell_1851 ( .C (CLK), .D (signal_3994), .Q (signal_3995) ) ;
    buf_clk cell_1859 ( .C (CLK), .D (signal_4002), .Q (signal_4003) ) ;
    buf_clk cell_1863 ( .C (CLK), .D (signal_4006), .Q (signal_4007) ) ;
    buf_clk cell_1871 ( .C (CLK), .D (signal_4014), .Q (signal_4015) ) ;
    buf_clk cell_1875 ( .C (CLK), .D (signal_4018), .Q (signal_4019) ) ;
    buf_clk cell_1883 ( .C (CLK), .D (signal_4026), .Q (signal_4027) ) ;
    buf_clk cell_1887 ( .C (CLK), .D (signal_4030), .Q (signal_4031) ) ;
    buf_clk cell_1895 ( .C (CLK), .D (signal_4038), .Q (signal_4039) ) ;
    buf_clk cell_1899 ( .C (CLK), .D (signal_4042), .Q (signal_4043) ) ;
    buf_clk cell_1907 ( .C (CLK), .D (signal_4050), .Q (signal_4051) ) ;
    buf_clk cell_1911 ( .C (CLK), .D (signal_4054), .Q (signal_4055) ) ;
    buf_clk cell_1923 ( .C (CLK), .D (signal_4066), .Q (signal_4067) ) ;
    buf_clk cell_1927 ( .C (CLK), .D (signal_4070), .Q (signal_4071) ) ;
    buf_clk cell_1939 ( .C (CLK), .D (signal_4082), .Q (signal_4083) ) ;
    buf_clk cell_1943 ( .C (CLK), .D (signal_4086), .Q (signal_4087) ) ;
    buf_clk cell_1967 ( .C (CLK), .D (signal_4110), .Q (signal_4111) ) ;
    buf_clk cell_1971 ( .C (CLK), .D (signal_4114), .Q (signal_4115) ) ;
    buf_clk cell_1983 ( .C (CLK), .D (signal_4126), .Q (signal_4127) ) ;
    buf_clk cell_1987 ( .C (CLK), .D (signal_4130), .Q (signal_4131) ) ;
    buf_clk cell_1999 ( .C (CLK), .D (signal_4142), .Q (signal_4143) ) ;
    buf_clk cell_2003 ( .C (CLK), .D (signal_4146), .Q (signal_4147) ) ;
    buf_clk cell_2015 ( .C (CLK), .D (signal_4158), .Q (signal_4159) ) ;
    buf_clk cell_2019 ( .C (CLK), .D (signal_4162), .Q (signal_4163) ) ;
    buf_clk cell_2159 ( .C (CLK), .D (signal_4302), .Q (signal_4303) ) ;
    buf_clk cell_2163 ( .C (CLK), .D (signal_4306), .Q (signal_4307) ) ;
    buf_clk cell_2175 ( .C (CLK), .D (signal_4318), .Q (signal_4319) ) ;
    buf_clk cell_2179 ( .C (CLK), .D (signal_4322), .Q (signal_4323) ) ;
    buf_clk cell_2191 ( .C (CLK), .D (signal_4334), .Q (signal_4335) ) ;
    buf_clk cell_2199 ( .C (CLK), .D (signal_4342), .Q (signal_4343) ) ;
    buf_clk cell_2207 ( .C (CLK), .D (signal_4350), .Q (signal_4351) ) ;
    buf_clk cell_2215 ( .C (CLK), .D (signal_4358), .Q (signal_4359) ) ;
    buf_clk cell_2223 ( .C (CLK), .D (signal_4366), .Q (signal_4367) ) ;
    buf_clk cell_2231 ( .C (CLK), .D (signal_4374), .Q (signal_4375) ) ;
    buf_clk cell_2239 ( .C (CLK), .D (signal_4382), .Q (signal_4383) ) ;
    buf_clk cell_2247 ( .C (CLK), .D (signal_4390), .Q (signal_4391) ) ;
    buf_clk cell_2255 ( .C (CLK), .D (signal_4398), .Q (signal_4399) ) ;
    buf_clk cell_2263 ( .C (CLK), .D (signal_4406), .Q (signal_4407) ) ;
    buf_clk cell_2279 ( .C (CLK), .D (signal_4422), .Q (signal_4423) ) ;
    buf_clk cell_2287 ( .C (CLK), .D (signal_4430), .Q (signal_4431) ) ;
    buf_clk cell_2311 ( .C (CLK), .D (signal_4454), .Q (signal_4455) ) ;
    buf_clk cell_2319 ( .C (CLK), .D (signal_4462), .Q (signal_4463) ) ;
    buf_clk cell_2327 ( .C (CLK), .D (signal_4470), .Q (signal_4471) ) ;
    buf_clk cell_2335 ( .C (CLK), .D (signal_4478), .Q (signal_4479) ) ;
    buf_clk cell_2351 ( .C (CLK), .D (signal_4494), .Q (signal_4495) ) ;
    buf_clk cell_2371 ( .C (CLK), .D (signal_4514), .Q (signal_4515) ) ;
    buf_clk cell_2379 ( .C (CLK), .D (signal_4522), .Q (signal_4523) ) ;
    buf_clk cell_2387 ( .C (CLK), .D (signal_4530), .Q (signal_4531) ) ;
    buf_clk cell_2395 ( .C (CLK), .D (signal_4538), .Q (signal_4539) ) ;
    buf_clk cell_2403 ( .C (CLK), .D (signal_4546), .Q (signal_4547) ) ;
    buf_clk cell_2411 ( .C (CLK), .D (signal_4554), .Q (signal_4555) ) ;
    buf_clk cell_2419 ( .C (CLK), .D (signal_4562), .Q (signal_4563) ) ;
    buf_clk cell_2427 ( .C (CLK), .D (signal_4570), .Q (signal_4571) ) ;
    buf_clk cell_2435 ( .C (CLK), .D (signal_4578), .Q (signal_4579) ) ;
    buf_clk cell_2443 ( .C (CLK), .D (signal_4586), .Q (signal_4587) ) ;
    buf_clk cell_2451 ( .C (CLK), .D (signal_4594), .Q (signal_4595) ) ;
    buf_clk cell_2459 ( .C (CLK), .D (signal_4602), .Q (signal_4603) ) ;
    buf_clk cell_2467 ( .C (CLK), .D (signal_4610), .Q (signal_4611) ) ;
    buf_clk cell_2475 ( .C (CLK), .D (signal_4618), .Q (signal_4619) ) ;
    buf_clk cell_2483 ( .C (CLK), .D (signal_4626), .Q (signal_4627) ) ;
    buf_clk cell_2491 ( .C (CLK), .D (signal_4634), .Q (signal_4635) ) ;
    buf_clk cell_2499 ( .C (CLK), .D (signal_4642), .Q (signal_4643) ) ;
    buf_clk cell_2507 ( .C (CLK), .D (signal_4650), .Q (signal_4651) ) ;
    buf_clk cell_2515 ( .C (CLK), .D (signal_4658), .Q (signal_4659) ) ;
    buf_clk cell_2523 ( .C (CLK), .D (signal_4666), .Q (signal_4667) ) ;
    buf_clk cell_2531 ( .C (CLK), .D (signal_4674), .Q (signal_4675) ) ;
    buf_clk cell_2539 ( .C (CLK), .D (signal_4682), .Q (signal_4683) ) ;
    buf_clk cell_2547 ( .C (CLK), .D (signal_4690), .Q (signal_4691) ) ;
    buf_clk cell_2555 ( .C (CLK), .D (signal_4698), .Q (signal_4699) ) ;
    buf_clk cell_2563 ( .C (CLK), .D (signal_4706), .Q (signal_4707) ) ;
    buf_clk cell_2587 ( .C (CLK), .D (signal_4730), .Q (signal_4731) ) ;
    buf_clk cell_2595 ( .C (CLK), .D (signal_4738), .Q (signal_4739) ) ;
    buf_clk cell_2603 ( .C (CLK), .D (signal_4746), .Q (signal_4747) ) ;
    buf_clk cell_2611 ( .C (CLK), .D (signal_4754), .Q (signal_4755) ) ;
    buf_clk cell_2639 ( .C (CLK), .D (signal_4782), .Q (signal_4783) ) ;
    buf_clk cell_2647 ( .C (CLK), .D (signal_4790), .Q (signal_4791) ) ;
    buf_clk cell_2655 ( .C (CLK), .D (signal_4798), .Q (signal_4799) ) ;
    buf_clk cell_2663 ( .C (CLK), .D (signal_4806), .Q (signal_4807) ) ;
    buf_clk cell_2691 ( .C (CLK), .D (signal_4834), .Q (signal_4835) ) ;
    buf_clk cell_2699 ( .C (CLK), .D (signal_4842), .Q (signal_4843) ) ;
    buf_clk cell_2707 ( .C (CLK), .D (signal_4850), .Q (signal_4851) ) ;
    buf_clk cell_2715 ( .C (CLK), .D (signal_4858), .Q (signal_4859) ) ;
    buf_clk cell_2723 ( .C (CLK), .D (signal_4866), .Q (signal_4867) ) ;
    buf_clk cell_2731 ( .C (CLK), .D (signal_4874), .Q (signal_4875) ) ;
    buf_clk cell_2739 ( .C (CLK), .D (signal_4882), .Q (signal_4883) ) ;
    buf_clk cell_2747 ( .C (CLK), .D (signal_4890), .Q (signal_4891) ) ;
    buf_clk cell_2755 ( .C (CLK), .D (signal_4898), .Q (signal_4899) ) ;
    buf_clk cell_2763 ( .C (CLK), .D (signal_4906), .Q (signal_4907) ) ;
    buf_clk cell_2771 ( .C (CLK), .D (signal_4914), .Q (signal_4915) ) ;
    buf_clk cell_2779 ( .C (CLK), .D (signal_4922), .Q (signal_4923) ) ;
    buf_clk cell_2787 ( .C (CLK), .D (signal_4930), .Q (signal_4931) ) ;
    buf_clk cell_2793 ( .C (CLK), .D (signal_4936), .Q (signal_4937) ) ;
    buf_clk cell_2799 ( .C (CLK), .D (signal_4942), .Q (signal_4943) ) ;
    buf_clk cell_2805 ( .C (CLK), .D (signal_4948), .Q (signal_4949) ) ;
    buf_clk cell_2811 ( .C (CLK), .D (signal_4954), .Q (signal_4955) ) ;
    buf_clk cell_2817 ( .C (CLK), .D (signal_4960), .Q (signal_4961) ) ;
    buf_clk cell_2823 ( .C (CLK), .D (signal_4966), .Q (signal_4967) ) ;
    buf_clk cell_2829 ( .C (CLK), .D (signal_4972), .Q (signal_4973) ) ;
    buf_clk cell_2835 ( .C (CLK), .D (signal_4978), .Q (signal_4979) ) ;
    buf_clk cell_2841 ( .C (CLK), .D (signal_4984), .Q (signal_4985) ) ;
    buf_clk cell_2847 ( .C (CLK), .D (signal_4990), .Q (signal_4991) ) ;
    buf_clk cell_2853 ( .C (CLK), .D (signal_4996), .Q (signal_4997) ) ;
    buf_clk cell_2859 ( .C (CLK), .D (signal_5002), .Q (signal_5003) ) ;
    buf_clk cell_2865 ( .C (CLK), .D (signal_5008), .Q (signal_5009) ) ;
    buf_clk cell_2971 ( .C (CLK), .D (signal_5114), .Q (signal_5115) ) ;
    buf_clk cell_2977 ( .C (CLK), .D (signal_5120), .Q (signal_5121) ) ;
    buf_clk cell_3055 ( .C (CLK), .D (signal_5198), .Q (signal_5199) ) ;
    buf_clk cell_3063 ( .C (CLK), .D (signal_5206), .Q (signal_5207) ) ;
    buf_clk cell_3447 ( .C (CLK), .D (signal_5590), .Q (signal_5591) ) ;
    buf_clk cell_3463 ( .C (CLK), .D (signal_5606), .Q (signal_5607) ) ;
    buf_clk cell_3487 ( .C (CLK), .D (signal_5630), .Q (signal_5631) ) ;
    buf_clk cell_3503 ( .C (CLK), .D (signal_5646), .Q (signal_5647) ) ;
    buf_clk cell_3527 ( .C (CLK), .D (signal_5670), .Q (signal_5671) ) ;
    buf_clk cell_3543 ( .C (CLK), .D (signal_5686), .Q (signal_5687) ) ;
    buf_clk cell_3559 ( .C (CLK), .D (signal_5702), .Q (signal_5703) ) ;
    buf_clk cell_3575 ( .C (CLK), .D (signal_5718), .Q (signal_5719) ) ;
    buf_clk cell_3635 ( .C (CLK), .D (signal_5778), .Q (signal_5779) ) ;
    buf_clk cell_3651 ( .C (CLK), .D (signal_5794), .Q (signal_5795) ) ;
    buf_clk cell_3667 ( .C (CLK), .D (signal_5810), .Q (signal_5811) ) ;
    buf_clk cell_3683 ( .C (CLK), .D (signal_5826), .Q (signal_5827) ) ;
    buf_clk cell_3699 ( .C (CLK), .D (signal_5842), .Q (signal_5843) ) ;
    buf_clk cell_3715 ( .C (CLK), .D (signal_5858), .Q (signal_5859) ) ;
    buf_clk cell_3731 ( .C (CLK), .D (signal_5874), .Q (signal_5875) ) ;
    buf_clk cell_3747 ( .C (CLK), .D (signal_5890), .Q (signal_5891) ) ;
    buf_clk cell_3763 ( .C (CLK), .D (signal_5906), .Q (signal_5907) ) ;
    buf_clk cell_3779 ( .C (CLK), .D (signal_5922), .Q (signal_5923) ) ;
    buf_clk cell_3887 ( .C (CLK), .D (signal_6030), .Q (signal_6031) ) ;
    buf_clk cell_3903 ( .C (CLK), .D (signal_6046), .Q (signal_6047) ) ;
    buf_clk cell_3919 ( .C (CLK), .D (signal_6062), .Q (signal_6063) ) ;
    buf_clk cell_3935 ( .C (CLK), .D (signal_6078), .Q (signal_6079) ) ;
    buf_clk cell_3951 ( .C (CLK), .D (signal_6094), .Q (signal_6095) ) ;
    buf_clk cell_3967 ( .C (CLK), .D (signal_6110), .Q (signal_6111) ) ;
    buf_clk cell_3983 ( .C (CLK), .D (signal_6126), .Q (signal_6127) ) ;
    buf_clk cell_3999 ( .C (CLK), .D (signal_6142), .Q (signal_6143) ) ;
    buf_clk cell_4015 ( .C (CLK), .D (signal_6158), .Q (signal_6159) ) ;
    buf_clk cell_4031 ( .C (CLK), .D (signal_6174), .Q (signal_6175) ) ;
    buf_clk cell_4047 ( .C (CLK), .D (signal_6190), .Q (signal_6191) ) ;
    buf_clk cell_4063 ( .C (CLK), .D (signal_6206), .Q (signal_6207) ) ;
    buf_clk cell_4079 ( .C (CLK), .D (signal_6222), .Q (signal_6223) ) ;
    buf_clk cell_4095 ( .C (CLK), .D (signal_6238), .Q (signal_6239) ) ;
    buf_clk cell_4179 ( .C (CLK), .D (signal_6322), .Q (signal_6323) ) ;
    buf_clk cell_4287 ( .C (CLK), .D (signal_6430), .Q (signal_6431) ) ;
    buf_clk cell_4303 ( .C (CLK), .D (signal_6446), .Q (signal_6447) ) ;
    buf_clk cell_4319 ( .C (CLK), .D (signal_6462), .Q (signal_6463) ) ;
    buf_clk cell_4335 ( .C (CLK), .D (signal_6478), .Q (signal_6479) ) ;
    buf_clk cell_4351 ( .C (CLK), .D (signal_6494), .Q (signal_6495) ) ;
    buf_clk cell_4367 ( .C (CLK), .D (signal_6510), .Q (signal_6511) ) ;
    buf_clk cell_4383 ( .C (CLK), .D (signal_6526), .Q (signal_6527) ) ;
    buf_clk cell_4399 ( .C (CLK), .D (signal_6542), .Q (signal_6543) ) ;
    buf_clk cell_4415 ( .C (CLK), .D (signal_6558), .Q (signal_6559) ) ;
    buf_clk cell_4431 ( .C (CLK), .D (signal_6574), .Q (signal_6575) ) ;
    buf_clk cell_4447 ( .C (CLK), .D (signal_6590), .Q (signal_6591) ) ;
    buf_clk cell_4463 ( .C (CLK), .D (signal_6606), .Q (signal_6607) ) ;
    buf_clk cell_4479 ( .C (CLK), .D (signal_6622), .Q (signal_6623) ) ;
    buf_clk cell_4495 ( .C (CLK), .D (signal_6638), .Q (signal_6639) ) ;
    buf_clk cell_4511 ( .C (CLK), .D (signal_6654), .Q (signal_6655) ) ;
    buf_clk cell_4527 ( .C (CLK), .D (signal_6670), .Q (signal_6671) ) ;
    buf_clk cell_4631 ( .C (CLK), .D (signal_6774), .Q (signal_6775) ) ;
    buf_clk cell_4647 ( .C (CLK), .D (signal_6790), .Q (signal_6791) ) ;
    buf_clk cell_4743 ( .C (CLK), .D (signal_6886), .Q (signal_6887) ) ;
    buf_clk cell_4759 ( .C (CLK), .D (signal_6902), .Q (signal_6903) ) ;
    buf_clk cell_4775 ( .C (CLK), .D (signal_6918), .Q (signal_6919) ) ;
    buf_clk cell_4791 ( .C (CLK), .D (signal_6934), .Q (signal_6935) ) ;
    buf_clk cell_4807 ( .C (CLK), .D (signal_6950), .Q (signal_6951) ) ;
    buf_clk cell_4823 ( .C (CLK), .D (signal_6966), .Q (signal_6967) ) ;
    buf_clk cell_4839 ( .C (CLK), .D (signal_6982), .Q (signal_6983) ) ;
    buf_clk cell_4855 ( .C (CLK), .D (signal_6998), .Q (signal_6999) ) ;
    buf_clk cell_4871 ( .C (CLK), .D (signal_7014), .Q (signal_7015) ) ;
    buf_clk cell_4887 ( .C (CLK), .D (signal_7030), .Q (signal_7031) ) ;
    buf_clk cell_4903 ( .C (CLK), .D (signal_7046), .Q (signal_7047) ) ;
    buf_clk cell_4919 ( .C (CLK), .D (signal_7062), .Q (signal_7063) ) ;
    buf_clk cell_4935 ( .C (CLK), .D (signal_7078), .Q (signal_7079) ) ;
    buf_clk cell_4951 ( .C (CLK), .D (signal_7094), .Q (signal_7095) ) ;
    buf_clk cell_4967 ( .C (CLK), .D (signal_7110), .Q (signal_7111) ) ;
    buf_clk cell_4983 ( .C (CLK), .D (signal_7126), .Q (signal_7127) ) ;
    buf_clk cell_4999 ( .C (CLK), .D (signal_7142), .Q (signal_7143) ) ;
    buf_clk cell_5015 ( .C (CLK), .D (signal_7158), .Q (signal_7159) ) ;
    buf_clk cell_5031 ( .C (CLK), .D (signal_7174), .Q (signal_7175) ) ;
    buf_clk cell_5047 ( .C (CLK), .D (signal_7190), .Q (signal_7191) ) ;
    buf_clk cell_5063 ( .C (CLK), .D (signal_7206), .Q (signal_7207) ) ;
    buf_clk cell_5079 ( .C (CLK), .D (signal_7222), .Q (signal_7223) ) ;
    buf_clk cell_5095 ( .C (CLK), .D (signal_7238), .Q (signal_7239) ) ;
    buf_clk cell_5111 ( .C (CLK), .D (signal_7254), .Q (signal_7255) ) ;
    buf_clk cell_5127 ( .C (CLK), .D (signal_7270), .Q (signal_7271) ) ;
    buf_clk cell_5143 ( .C (CLK), .D (signal_7286), .Q (signal_7287) ) ;
    buf_clk cell_5159 ( .C (CLK), .D (signal_7302), .Q (signal_7303) ) ;
    buf_clk cell_5175 ( .C (CLK), .D (signal_7318), .Q (signal_7319) ) ;
    buf_clk cell_5191 ( .C (CLK), .D (signal_7334), .Q (signal_7335) ) ;
    buf_clk cell_5207 ( .C (CLK), .D (signal_7350), .Q (signal_7351) ) ;
    buf_clk cell_5223 ( .C (CLK), .D (signal_7366), .Q (signal_7367) ) ;
    buf_clk cell_5239 ( .C (CLK), .D (signal_7382), .Q (signal_7383) ) ;
    buf_clk cell_5255 ( .C (CLK), .D (signal_7398), .Q (signal_7399) ) ;
    buf_clk cell_5271 ( .C (CLK), .D (signal_7414), .Q (signal_7415) ) ;
    buf_clk cell_5287 ( .C (CLK), .D (signal_7430), .Q (signal_7431) ) ;
    buf_clk cell_5303 ( .C (CLK), .D (signal_7446), .Q (signal_7447) ) ;
    buf_clk cell_5319 ( .C (CLK), .D (signal_7462), .Q (signal_7463) ) ;
    buf_clk cell_5335 ( .C (CLK), .D (signal_7478), .Q (signal_7479) ) ;
    buf_clk cell_5351 ( .C (CLK), .D (signal_7494), .Q (signal_7495) ) ;
    buf_clk cell_5367 ( .C (CLK), .D (signal_7510), .Q (signal_7511) ) ;
    buf_clk cell_5383 ( .C (CLK), .D (signal_7526), .Q (signal_7527) ) ;
    buf_clk cell_5399 ( .C (CLK), .D (signal_7542), .Q (signal_7543) ) ;
    buf_clk cell_5415 ( .C (CLK), .D (signal_7558), .Q (signal_7559) ) ;
    buf_clk cell_5431 ( .C (CLK), .D (signal_7574), .Q (signal_7575) ) ;
    buf_clk cell_5447 ( .C (CLK), .D (signal_7590), .Q (signal_7591) ) ;
    buf_clk cell_5463 ( .C (CLK), .D (signal_7606), .Q (signal_7607) ) ;
    buf_clk cell_5479 ( .C (CLK), .D (signal_7622), .Q (signal_7623) ) ;
    buf_clk cell_5495 ( .C (CLK), .D (signal_7638), .Q (signal_7639) ) ;
    buf_clk cell_5511 ( .C (CLK), .D (signal_7654), .Q (signal_7655) ) ;
    buf_clk cell_5527 ( .C (CLK), .D (signal_7670), .Q (signal_7671) ) ;
    buf_clk cell_5543 ( .C (CLK), .D (signal_7686), .Q (signal_7687) ) ;
    buf_clk cell_5559 ( .C (CLK), .D (signal_7702), .Q (signal_7703) ) ;
    buf_clk cell_5575 ( .C (CLK), .D (signal_7718), .Q (signal_7719) ) ;
    buf_clk cell_5591 ( .C (CLK), .D (signal_7734), .Q (signal_7735) ) ;
    buf_clk cell_5607 ( .C (CLK), .D (signal_7750), .Q (signal_7751) ) ;
    buf_clk cell_5623 ( .C (CLK), .D (signal_7766), .Q (signal_7767) ) ;
    buf_clk cell_5639 ( .C (CLK), .D (signal_7782), .Q (signal_7783) ) ;
    buf_clk cell_5655 ( .C (CLK), .D (signal_7798), .Q (signal_7799) ) ;
    buf_clk cell_5671 ( .C (CLK), .D (signal_7814), .Q (signal_7815) ) ;
    buf_clk cell_5687 ( .C (CLK), .D (signal_7830), .Q (signal_7831) ) ;
    buf_clk cell_5703 ( .C (CLK), .D (signal_7846), .Q (signal_7847) ) ;
    buf_clk cell_5719 ( .C (CLK), .D (signal_7862), .Q (signal_7863) ) ;
    buf_clk cell_5735 ( .C (CLK), .D (signal_7878), .Q (signal_7879) ) ;
    buf_clk cell_5751 ( .C (CLK), .D (signal_7894), .Q (signal_7895) ) ;
    buf_clk cell_5767 ( .C (CLK), .D (signal_7910), .Q (signal_7911) ) ;
    buf_clk cell_5783 ( .C (CLK), .D (signal_7926), .Q (signal_7927) ) ;
    buf_clk cell_5799 ( .C (CLK), .D (signal_7942), .Q (signal_7943) ) ;
    buf_clk cell_5815 ( .C (CLK), .D (signal_7958), .Q (signal_7959) ) ;
    buf_clk cell_5831 ( .C (CLK), .D (signal_7974), .Q (signal_7975) ) ;
    buf_clk cell_5847 ( .C (CLK), .D (signal_7990), .Q (signal_7991) ) ;
    buf_clk cell_5863 ( .C (CLK), .D (signal_8006), .Q (signal_8007) ) ;
    buf_clk cell_5879 ( .C (CLK), .D (signal_8022), .Q (signal_8023) ) ;
    buf_clk cell_5895 ( .C (CLK), .D (signal_8038), .Q (signal_8039) ) ;
    buf_clk cell_5911 ( .C (CLK), .D (signal_8054), .Q (signal_8055) ) ;
    buf_clk cell_5927 ( .C (CLK), .D (signal_8070), .Q (signal_8071) ) ;
    buf_clk cell_5943 ( .C (CLK), .D (signal_8086), .Q (signal_8087) ) ;
    buf_clk cell_5959 ( .C (CLK), .D (signal_8102), .Q (signal_8103) ) ;
    buf_clk cell_5975 ( .C (CLK), .D (signal_8118), .Q (signal_8119) ) ;
    buf_clk cell_5991 ( .C (CLK), .D (signal_8134), .Q (signal_8135) ) ;
    buf_clk cell_6007 ( .C (CLK), .D (signal_8150), .Q (signal_8151) ) ;
    buf_clk cell_6023 ( .C (CLK), .D (signal_8166), .Q (signal_8167) ) ;
    buf_clk cell_6039 ( .C (CLK), .D (signal_8182), .Q (signal_8183) ) ;
    buf_clk cell_6055 ( .C (CLK), .D (signal_8198), .Q (signal_8199) ) ;
    buf_clk cell_6071 ( .C (CLK), .D (signal_8214), .Q (signal_8215) ) ;
    buf_clk cell_6087 ( .C (CLK), .D (signal_8230), .Q (signal_8231) ) ;
    buf_clk cell_6103 ( .C (CLK), .D (signal_8246), .Q (signal_8247) ) ;
    buf_clk cell_6119 ( .C (CLK), .D (signal_8262), .Q (signal_8263) ) ;
    buf_clk cell_6135 ( .C (CLK), .D (signal_8278), .Q (signal_8279) ) ;
    buf_clk cell_6151 ( .C (CLK), .D (signal_8294), .Q (signal_8295) ) ;
    buf_clk cell_6167 ( .C (CLK), .D (signal_8310), .Q (signal_8311) ) ;
    buf_clk cell_6183 ( .C (CLK), .D (signal_8326), .Q (signal_8327) ) ;
    buf_clk cell_6199 ( .C (CLK), .D (signal_8342), .Q (signal_8343) ) ;
    buf_clk cell_6215 ( .C (CLK), .D (signal_8358), .Q (signal_8359) ) ;
    buf_clk cell_6231 ( .C (CLK), .D (signal_8374), .Q (signal_8375) ) ;
    buf_clk cell_6247 ( .C (CLK), .D (signal_8390), .Q (signal_8391) ) ;
    buf_clk cell_6263 ( .C (CLK), .D (signal_8406), .Q (signal_8407) ) ;
    buf_clk cell_6279 ( .C (CLK), .D (signal_8422), .Q (signal_8423) ) ;
    buf_clk cell_6295 ( .C (CLK), .D (signal_8438), .Q (signal_8439) ) ;
    buf_clk cell_6311 ( .C (CLK), .D (signal_8454), .Q (signal_8455) ) ;
    buf_clk cell_6327 ( .C (CLK), .D (signal_8470), .Q (signal_8471) ) ;
    buf_clk cell_6343 ( .C (CLK), .D (signal_8486), .Q (signal_8487) ) ;
    buf_clk cell_6359 ( .C (CLK), .D (signal_8502), .Q (signal_8503) ) ;
    buf_clk cell_6375 ( .C (CLK), .D (signal_8518), .Q (signal_8519) ) ;
    buf_clk cell_6391 ( .C (CLK), .D (signal_8534), .Q (signal_8535) ) ;
    buf_clk cell_7591 ( .C (CLK), .D (signal_9734), .Q (signal_9735) ) ;
    buf_clk cell_7607 ( .C (CLK), .D (signal_9750), .Q (signal_9751) ) ;
    buf_clk cell_7623 ( .C (CLK), .D (signal_9766), .Q (signal_9767) ) ;
    buf_clk cell_7639 ( .C (CLK), .D (signal_9782), .Q (signal_9783) ) ;
    buf_clk cell_7655 ( .C (CLK), .D (signal_9798), .Q (signal_9799) ) ;
    buf_clk cell_7671 ( .C (CLK), .D (signal_9814), .Q (signal_9815) ) ;
    buf_clk cell_7687 ( .C (CLK), .D (signal_9830), .Q (signal_9831) ) ;
    buf_clk cell_7703 ( .C (CLK), .D (signal_9846), .Q (signal_9847) ) ;
    buf_clk cell_7719 ( .C (CLK), .D (signal_9862), .Q (signal_9863) ) ;
    buf_clk cell_7735 ( .C (CLK), .D (signal_9878), .Q (signal_9879) ) ;
    buf_clk cell_7943 ( .C (CLK), .D (signal_10086), .Q (signal_10087) ) ;

    /* cells in depth 3 */
    buf_clk cell_1812 ( .C (CLK), .D (signal_3955), .Q (signal_3956) ) ;
    buf_clk cell_1816 ( .C (CLK), .D (signal_3959), .Q (signal_3960) ) ;
    buf_clk cell_1818 ( .C (CLK), .D (signal_1329), .Q (signal_3962) ) ;
    buf_clk cell_1820 ( .C (CLK), .D (signal_2267), .Q (signal_3964) ) ;
    buf_clk cell_1824 ( .C (CLK), .D (signal_3967), .Q (signal_3968) ) ;
    buf_clk cell_1828 ( .C (CLK), .D (signal_3971), .Q (signal_3972) ) ;
    buf_clk cell_1830 ( .C (CLK), .D (signal_1331), .Q (signal_3974) ) ;
    buf_clk cell_1832 ( .C (CLK), .D (signal_2269), .Q (signal_3976) ) ;
    buf_clk cell_1836 ( .C (CLK), .D (signal_3979), .Q (signal_3980) ) ;
    buf_clk cell_1840 ( .C (CLK), .D (signal_3983), .Q (signal_3984) ) ;
    buf_clk cell_1842 ( .C (CLK), .D (signal_1333), .Q (signal_3986) ) ;
    buf_clk cell_1844 ( .C (CLK), .D (signal_2271), .Q (signal_3988) ) ;
    buf_clk cell_1848 ( .C (CLK), .D (signal_3991), .Q (signal_3992) ) ;
    buf_clk cell_1852 ( .C (CLK), .D (signal_3995), .Q (signal_3996) ) ;
    buf_clk cell_1854 ( .C (CLK), .D (signal_1335), .Q (signal_3998) ) ;
    buf_clk cell_1856 ( .C (CLK), .D (signal_2273), .Q (signal_4000) ) ;
    buf_clk cell_1860 ( .C (CLK), .D (signal_4003), .Q (signal_4004) ) ;
    buf_clk cell_1864 ( .C (CLK), .D (signal_4007), .Q (signal_4008) ) ;
    buf_clk cell_1866 ( .C (CLK), .D (signal_1337), .Q (signal_4010) ) ;
    buf_clk cell_1868 ( .C (CLK), .D (signal_2275), .Q (signal_4012) ) ;
    buf_clk cell_1872 ( .C (CLK), .D (signal_4015), .Q (signal_4016) ) ;
    buf_clk cell_1876 ( .C (CLK), .D (signal_4019), .Q (signal_4020) ) ;
    buf_clk cell_1878 ( .C (CLK), .D (signal_1339), .Q (signal_4022) ) ;
    buf_clk cell_1880 ( .C (CLK), .D (signal_2277), .Q (signal_4024) ) ;
    buf_clk cell_1884 ( .C (CLK), .D (signal_4027), .Q (signal_4028) ) ;
    buf_clk cell_1888 ( .C (CLK), .D (signal_4031), .Q (signal_4032) ) ;
    buf_clk cell_1890 ( .C (CLK), .D (signal_1341), .Q (signal_4034) ) ;
    buf_clk cell_1892 ( .C (CLK), .D (signal_2279), .Q (signal_4036) ) ;
    buf_clk cell_1896 ( .C (CLK), .D (signal_4039), .Q (signal_4040) ) ;
    buf_clk cell_1900 ( .C (CLK), .D (signal_4043), .Q (signal_4044) ) ;
    buf_clk cell_1902 ( .C (CLK), .D (signal_1343), .Q (signal_4046) ) ;
    buf_clk cell_1904 ( .C (CLK), .D (signal_2281), .Q (signal_4048) ) ;
    buf_clk cell_1908 ( .C (CLK), .D (signal_4051), .Q (signal_4052) ) ;
    buf_clk cell_1912 ( .C (CLK), .D (signal_4055), .Q (signal_4056) ) ;
    buf_clk cell_1914 ( .C (CLK), .D (signal_1344), .Q (signal_4058) ) ;
    buf_clk cell_1916 ( .C (CLK), .D (signal_2290), .Q (signal_4060) ) ;
    buf_clk cell_1918 ( .C (CLK), .D (signal_1346), .Q (signal_4062) ) ;
    buf_clk cell_1920 ( .C (CLK), .D (signal_2292), .Q (signal_4064) ) ;
    buf_clk cell_1924 ( .C (CLK), .D (signal_4067), .Q (signal_4068) ) ;
    buf_clk cell_1928 ( .C (CLK), .D (signal_4071), .Q (signal_4072) ) ;
    buf_clk cell_1930 ( .C (CLK), .D (signal_1347), .Q (signal_4074) ) ;
    buf_clk cell_1932 ( .C (CLK), .D (signal_2293), .Q (signal_4076) ) ;
    buf_clk cell_1934 ( .C (CLK), .D (signal_1349), .Q (signal_4078) ) ;
    buf_clk cell_1936 ( .C (CLK), .D (signal_2295), .Q (signal_4080) ) ;
    buf_clk cell_1940 ( .C (CLK), .D (signal_4083), .Q (signal_4084) ) ;
    buf_clk cell_1944 ( .C (CLK), .D (signal_4087), .Q (signal_4088) ) ;
    buf_clk cell_1946 ( .C (CLK), .D (signal_1350), .Q (signal_4090) ) ;
    buf_clk cell_1948 ( .C (CLK), .D (signal_2296), .Q (signal_4092) ) ;
    buf_clk cell_1950 ( .C (CLK), .D (signal_1352), .Q (signal_4094) ) ;
    buf_clk cell_1952 ( .C (CLK), .D (signal_2298), .Q (signal_4096) ) ;
    buf_clk cell_1954 ( .C (CLK), .D (signal_3951), .Q (signal_4098) ) ;
    buf_clk cell_1956 ( .C (CLK), .D (signal_3953), .Q (signal_4100) ) ;
    buf_clk cell_1958 ( .C (CLK), .D (signal_1353), .Q (signal_4102) ) ;
    buf_clk cell_1960 ( .C (CLK), .D (signal_2299), .Q (signal_4104) ) ;
    buf_clk cell_1962 ( .C (CLK), .D (signal_1355), .Q (signal_4106) ) ;
    buf_clk cell_1964 ( .C (CLK), .D (signal_2301), .Q (signal_4108) ) ;
    buf_clk cell_1968 ( .C (CLK), .D (signal_4111), .Q (signal_4112) ) ;
    buf_clk cell_1972 ( .C (CLK), .D (signal_4115), .Q (signal_4116) ) ;
    buf_clk cell_1974 ( .C (CLK), .D (signal_1356), .Q (signal_4118) ) ;
    buf_clk cell_1976 ( .C (CLK), .D (signal_2282), .Q (signal_4120) ) ;
    buf_clk cell_1978 ( .C (CLK), .D (signal_1358), .Q (signal_4122) ) ;
    buf_clk cell_1980 ( .C (CLK), .D (signal_2303), .Q (signal_4124) ) ;
    buf_clk cell_1984 ( .C (CLK), .D (signal_4127), .Q (signal_4128) ) ;
    buf_clk cell_1988 ( .C (CLK), .D (signal_4131), .Q (signal_4132) ) ;
    buf_clk cell_1990 ( .C (CLK), .D (signal_1359), .Q (signal_4134) ) ;
    buf_clk cell_1992 ( .C (CLK), .D (signal_2304), .Q (signal_4136) ) ;
    buf_clk cell_1994 ( .C (CLK), .D (signal_1361), .Q (signal_4138) ) ;
    buf_clk cell_1996 ( .C (CLK), .D (signal_2306), .Q (signal_4140) ) ;
    buf_clk cell_2000 ( .C (CLK), .D (signal_4143), .Q (signal_4144) ) ;
    buf_clk cell_2004 ( .C (CLK), .D (signal_4147), .Q (signal_4148) ) ;
    buf_clk cell_2006 ( .C (CLK), .D (signal_1362), .Q (signal_4150) ) ;
    buf_clk cell_2008 ( .C (CLK), .D (signal_2307), .Q (signal_4152) ) ;
    buf_clk cell_2010 ( .C (CLK), .D (signal_1364), .Q (signal_4154) ) ;
    buf_clk cell_2012 ( .C (CLK), .D (signal_2309), .Q (signal_4156) ) ;
    buf_clk cell_2016 ( .C (CLK), .D (signal_4159), .Q (signal_4160) ) ;
    buf_clk cell_2020 ( .C (CLK), .D (signal_4163), .Q (signal_4164) ) ;
    buf_clk cell_2022 ( .C (CLK), .D (signal_1365), .Q (signal_4166) ) ;
    buf_clk cell_2024 ( .C (CLK), .D (signal_2310), .Q (signal_4168) ) ;
    buf_clk cell_2026 ( .C (CLK), .D (signal_1367), .Q (signal_4170) ) ;
    buf_clk cell_2028 ( .C (CLK), .D (signal_2312), .Q (signal_4172) ) ;
    buf_clk cell_2030 ( .C (CLK), .D (signal_1336), .Q (signal_4174) ) ;
    buf_clk cell_2032 ( .C (CLK), .D (signal_2274), .Q (signal_4176) ) ;
    buf_clk cell_2034 ( .C (CLK), .D (signal_1368), .Q (signal_4178) ) ;
    buf_clk cell_2036 ( .C (CLK), .D (signal_2283), .Q (signal_4180) ) ;
    buf_clk cell_2038 ( .C (CLK), .D (signal_1369), .Q (signal_4182) ) ;
    buf_clk cell_2040 ( .C (CLK), .D (signal_2284), .Q (signal_4184) ) ;
    buf_clk cell_2042 ( .C (CLK), .D (signal_1342), .Q (signal_4186) ) ;
    buf_clk cell_2044 ( .C (CLK), .D (signal_2280), .Q (signal_4188) ) ;
    buf_clk cell_2046 ( .C (CLK), .D (signal_1338), .Q (signal_4190) ) ;
    buf_clk cell_2048 ( .C (CLK), .D (signal_2276), .Q (signal_4192) ) ;
    buf_clk cell_2050 ( .C (CLK), .D (signal_1370), .Q (signal_4194) ) ;
    buf_clk cell_2052 ( .C (CLK), .D (signal_2285), .Q (signal_4196) ) ;
    buf_clk cell_2054 ( .C (CLK), .D (signal_1334), .Q (signal_4198) ) ;
    buf_clk cell_2056 ( .C (CLK), .D (signal_2272), .Q (signal_4200) ) ;
    buf_clk cell_2058 ( .C (CLK), .D (signal_1371), .Q (signal_4202) ) ;
    buf_clk cell_2060 ( .C (CLK), .D (signal_2313), .Q (signal_4204) ) ;
    buf_clk cell_2062 ( .C (CLK), .D (signal_1360), .Q (signal_4206) ) ;
    buf_clk cell_2064 ( .C (CLK), .D (signal_2305), .Q (signal_4208) ) ;
    buf_clk cell_2066 ( .C (CLK), .D (signal_1372), .Q (signal_4210) ) ;
    buf_clk cell_2068 ( .C (CLK), .D (signal_2314), .Q (signal_4212) ) ;
    buf_clk cell_2070 ( .C (CLK), .D (signal_1351), .Q (signal_4214) ) ;
    buf_clk cell_2072 ( .C (CLK), .D (signal_2297), .Q (signal_4216) ) ;
    buf_clk cell_2074 ( .C (CLK), .D (signal_1340), .Q (signal_4218) ) ;
    buf_clk cell_2076 ( .C (CLK), .D (signal_2278), .Q (signal_4220) ) ;
    buf_clk cell_2078 ( .C (CLK), .D (signal_1373), .Q (signal_4222) ) ;
    buf_clk cell_2080 ( .C (CLK), .D (signal_2315), .Q (signal_4224) ) ;
    buf_clk cell_2082 ( .C (CLK), .D (signal_3887), .Q (signal_4226) ) ;
    buf_clk cell_2084 ( .C (CLK), .D (signal_3889), .Q (signal_4228) ) ;
    buf_clk cell_2086 ( .C (CLK), .D (signal_3935), .Q (signal_4230) ) ;
    buf_clk cell_2088 ( .C (CLK), .D (signal_3937), .Q (signal_4232) ) ;
    buf_clk cell_2090 ( .C (CLK), .D (signal_3915), .Q (signal_4234) ) ;
    buf_clk cell_2092 ( .C (CLK), .D (signal_3917), .Q (signal_4236) ) ;
    buf_clk cell_2094 ( .C (CLK), .D (signal_3903), .Q (signal_4238) ) ;
    buf_clk cell_2096 ( .C (CLK), .D (signal_3905), .Q (signal_4240) ) ;
    buf_clk cell_2098 ( .C (CLK), .D (signal_1374), .Q (signal_4242) ) ;
    buf_clk cell_2100 ( .C (CLK), .D (signal_2316), .Q (signal_4244) ) ;
    buf_clk cell_2102 ( .C (CLK), .D (signal_1332), .Q (signal_4246) ) ;
    buf_clk cell_2104 ( .C (CLK), .D (signal_2270), .Q (signal_4248) ) ;
    buf_clk cell_2106 ( .C (CLK), .D (signal_1363), .Q (signal_4250) ) ;
    buf_clk cell_2108 ( .C (CLK), .D (signal_2308), .Q (signal_4252) ) ;
    buf_clk cell_2110 ( .C (CLK), .D (signal_1375), .Q (signal_4254) ) ;
    buf_clk cell_2112 ( .C (CLK), .D (signal_2317), .Q (signal_4256) ) ;
    buf_clk cell_2114 ( .C (CLK), .D (signal_1357), .Q (signal_4258) ) ;
    buf_clk cell_2116 ( .C (CLK), .D (signal_2302), .Q (signal_4260) ) ;
    buf_clk cell_2118 ( .C (CLK), .D (signal_1376), .Q (signal_4262) ) ;
    buf_clk cell_2120 ( .C (CLK), .D (signal_2318), .Q (signal_4264) ) ;
    buf_clk cell_2122 ( .C (CLK), .D (signal_1377), .Q (signal_4266) ) ;
    buf_clk cell_2124 ( .C (CLK), .D (signal_2286), .Q (signal_4268) ) ;
    buf_clk cell_2126 ( .C (CLK), .D (signal_1378), .Q (signal_4270) ) ;
    buf_clk cell_2128 ( .C (CLK), .D (signal_2287), .Q (signal_4272) ) ;
    buf_clk cell_2130 ( .C (CLK), .D (signal_1366), .Q (signal_4274) ) ;
    buf_clk cell_2132 ( .C (CLK), .D (signal_2311), .Q (signal_4276) ) ;
    buf_clk cell_2134 ( .C (CLK), .D (signal_1328), .Q (signal_4278) ) ;
    buf_clk cell_2136 ( .C (CLK), .D (signal_2266), .Q (signal_4280) ) ;
    buf_clk cell_2138 ( .C (CLK), .D (signal_1379), .Q (signal_4282) ) ;
    buf_clk cell_2140 ( .C (CLK), .D (signal_2288), .Q (signal_4284) ) ;
    buf_clk cell_2142 ( .C (CLK), .D (signal_1380), .Q (signal_4286) ) ;
    buf_clk cell_2144 ( .C (CLK), .D (signal_2289), .Q (signal_4288) ) ;
    buf_clk cell_2146 ( .C (CLK), .D (signal_3923), .Q (signal_4290) ) ;
    buf_clk cell_2148 ( .C (CLK), .D (signal_3925), .Q (signal_4292) ) ;
    buf_clk cell_2150 ( .C (CLK), .D (signal_3943), .Q (signal_4294) ) ;
    buf_clk cell_2152 ( .C (CLK), .D (signal_3945), .Q (signal_4296) ) ;
    buf_clk cell_2154 ( .C (CLK), .D (signal_1381), .Q (signal_4298) ) ;
    buf_clk cell_2156 ( .C (CLK), .D (signal_2319), .Q (signal_4300) ) ;
    buf_clk cell_2160 ( .C (CLK), .D (signal_4303), .Q (signal_4304) ) ;
    buf_clk cell_2164 ( .C (CLK), .D (signal_4307), .Q (signal_4308) ) ;
    buf_clk cell_2166 ( .C (CLK), .D (signal_1345), .Q (signal_4310) ) ;
    buf_clk cell_2168 ( .C (CLK), .D (signal_2291), .Q (signal_4312) ) ;
    buf_clk cell_2170 ( .C (CLK), .D (signal_3947), .Q (signal_4314) ) ;
    buf_clk cell_2172 ( .C (CLK), .D (signal_3949), .Q (signal_4316) ) ;
    buf_clk cell_2176 ( .C (CLK), .D (signal_4319), .Q (signal_4320) ) ;
    buf_clk cell_2180 ( .C (CLK), .D (signal_4323), .Q (signal_4324) ) ;
    buf_clk cell_2182 ( .C (CLK), .D (signal_3875), .Q (signal_4326) ) ;
    buf_clk cell_2184 ( .C (CLK), .D (signal_3877), .Q (signal_4328) ) ;
    buf_clk cell_2186 ( .C (CLK), .D (signal_1330), .Q (signal_4330) ) ;
    buf_clk cell_2188 ( .C (CLK), .D (signal_2268), .Q (signal_4332) ) ;
    buf_clk cell_2192 ( .C (CLK), .D (signal_4335), .Q (signal_4336) ) ;
    buf_clk cell_2200 ( .C (CLK), .D (signal_4343), .Q (signal_4344) ) ;
    buf_clk cell_2208 ( .C (CLK), .D (signal_4351), .Q (signal_4352) ) ;
    buf_clk cell_2216 ( .C (CLK), .D (signal_4359), .Q (signal_4360) ) ;
    buf_clk cell_2224 ( .C (CLK), .D (signal_4367), .Q (signal_4368) ) ;
    buf_clk cell_2232 ( .C (CLK), .D (signal_4375), .Q (signal_4376) ) ;
    buf_clk cell_2240 ( .C (CLK), .D (signal_4383), .Q (signal_4384) ) ;
    buf_clk cell_2248 ( .C (CLK), .D (signal_4391), .Q (signal_4392) ) ;
    buf_clk cell_2256 ( .C (CLK), .D (signal_4399), .Q (signal_4400) ) ;
    buf_clk cell_2264 ( .C (CLK), .D (signal_4407), .Q (signal_4408) ) ;
    buf_clk cell_2280 ( .C (CLK), .D (signal_4423), .Q (signal_4424) ) ;
    buf_clk cell_2288 ( .C (CLK), .D (signal_4431), .Q (signal_4432) ) ;
    buf_clk cell_2312 ( .C (CLK), .D (signal_4455), .Q (signal_4456) ) ;
    buf_clk cell_2320 ( .C (CLK), .D (signal_4463), .Q (signal_4464) ) ;
    buf_clk cell_2328 ( .C (CLK), .D (signal_4471), .Q (signal_4472) ) ;
    buf_clk cell_2336 ( .C (CLK), .D (signal_4479), .Q (signal_4480) ) ;
    buf_clk cell_2352 ( .C (CLK), .D (signal_4495), .Q (signal_4496) ) ;
    buf_clk cell_2358 ( .C (CLK), .D (signal_3883), .Q (signal_4502) ) ;
    buf_clk cell_2364 ( .C (CLK), .D (signal_3885), .Q (signal_4508) ) ;
    buf_clk cell_2372 ( .C (CLK), .D (signal_4515), .Q (signal_4516) ) ;
    buf_clk cell_2380 ( .C (CLK), .D (signal_4523), .Q (signal_4524) ) ;
    buf_clk cell_2388 ( .C (CLK), .D (signal_4531), .Q (signal_4532) ) ;
    buf_clk cell_2396 ( .C (CLK), .D (signal_4539), .Q (signal_4540) ) ;
    buf_clk cell_2404 ( .C (CLK), .D (signal_4547), .Q (signal_4548) ) ;
    buf_clk cell_2412 ( .C (CLK), .D (signal_4555), .Q (signal_4556) ) ;
    buf_clk cell_2420 ( .C (CLK), .D (signal_4563), .Q (signal_4564) ) ;
    buf_clk cell_2428 ( .C (CLK), .D (signal_4571), .Q (signal_4572) ) ;
    buf_clk cell_2436 ( .C (CLK), .D (signal_4579), .Q (signal_4580) ) ;
    buf_clk cell_2444 ( .C (CLK), .D (signal_4587), .Q (signal_4588) ) ;
    buf_clk cell_2452 ( .C (CLK), .D (signal_4595), .Q (signal_4596) ) ;
    buf_clk cell_2460 ( .C (CLK), .D (signal_4603), .Q (signal_4604) ) ;
    buf_clk cell_2468 ( .C (CLK), .D (signal_4611), .Q (signal_4612) ) ;
    buf_clk cell_2476 ( .C (CLK), .D (signal_4619), .Q (signal_4620) ) ;
    buf_clk cell_2484 ( .C (CLK), .D (signal_4627), .Q (signal_4628) ) ;
    buf_clk cell_2492 ( .C (CLK), .D (signal_4635), .Q (signal_4636) ) ;
    buf_clk cell_2500 ( .C (CLK), .D (signal_4643), .Q (signal_4644) ) ;
    buf_clk cell_2508 ( .C (CLK), .D (signal_4651), .Q (signal_4652) ) ;
    buf_clk cell_2516 ( .C (CLK), .D (signal_4659), .Q (signal_4660) ) ;
    buf_clk cell_2524 ( .C (CLK), .D (signal_4667), .Q (signal_4668) ) ;
    buf_clk cell_2532 ( .C (CLK), .D (signal_4675), .Q (signal_4676) ) ;
    buf_clk cell_2540 ( .C (CLK), .D (signal_4683), .Q (signal_4684) ) ;
    buf_clk cell_2548 ( .C (CLK), .D (signal_4691), .Q (signal_4692) ) ;
    buf_clk cell_2556 ( .C (CLK), .D (signal_4699), .Q (signal_4700) ) ;
    buf_clk cell_2564 ( .C (CLK), .D (signal_4707), .Q (signal_4708) ) ;
    buf_clk cell_2588 ( .C (CLK), .D (signal_4731), .Q (signal_4732) ) ;
    buf_clk cell_2596 ( .C (CLK), .D (signal_4739), .Q (signal_4740) ) ;
    buf_clk cell_2604 ( .C (CLK), .D (signal_4747), .Q (signal_4748) ) ;
    buf_clk cell_2612 ( .C (CLK), .D (signal_4755), .Q (signal_4756) ) ;
    buf_clk cell_2626 ( .C (CLK), .D (signal_3939), .Q (signal_4770) ) ;
    buf_clk cell_2632 ( .C (CLK), .D (signal_3941), .Q (signal_4776) ) ;
    buf_clk cell_2640 ( .C (CLK), .D (signal_4783), .Q (signal_4784) ) ;
    buf_clk cell_2648 ( .C (CLK), .D (signal_4791), .Q (signal_4792) ) ;
    buf_clk cell_2656 ( .C (CLK), .D (signal_4799), .Q (signal_4800) ) ;
    buf_clk cell_2664 ( .C (CLK), .D (signal_4807), .Q (signal_4808) ) ;
    buf_clk cell_2670 ( .C (CLK), .D (signal_3919), .Q (signal_4814) ) ;
    buf_clk cell_2676 ( .C (CLK), .D (signal_3921), .Q (signal_4820) ) ;
    buf_clk cell_2692 ( .C (CLK), .D (signal_4835), .Q (signal_4836) ) ;
    buf_clk cell_2700 ( .C (CLK), .D (signal_4843), .Q (signal_4844) ) ;
    buf_clk cell_2708 ( .C (CLK), .D (signal_4851), .Q (signal_4852) ) ;
    buf_clk cell_2716 ( .C (CLK), .D (signal_4859), .Q (signal_4860) ) ;
    buf_clk cell_2724 ( .C (CLK), .D (signal_4867), .Q (signal_4868) ) ;
    buf_clk cell_2732 ( .C (CLK), .D (signal_4875), .Q (signal_4876) ) ;
    buf_clk cell_2740 ( .C (CLK), .D (signal_4883), .Q (signal_4884) ) ;
    buf_clk cell_2748 ( .C (CLK), .D (signal_4891), .Q (signal_4892) ) ;
    buf_clk cell_2756 ( .C (CLK), .D (signal_4899), .Q (signal_4900) ) ;
    buf_clk cell_2764 ( .C (CLK), .D (signal_4907), .Q (signal_4908) ) ;
    buf_clk cell_2772 ( .C (CLK), .D (signal_4915), .Q (signal_4916) ) ;
    buf_clk cell_2780 ( .C (CLK), .D (signal_4923), .Q (signal_4924) ) ;
    buf_clk cell_2788 ( .C (CLK), .D (signal_4931), .Q (signal_4932) ) ;
    buf_clk cell_2794 ( .C (CLK), .D (signal_4937), .Q (signal_4938) ) ;
    buf_clk cell_2800 ( .C (CLK), .D (signal_4943), .Q (signal_4944) ) ;
    buf_clk cell_2806 ( .C (CLK), .D (signal_4949), .Q (signal_4950) ) ;
    buf_clk cell_2812 ( .C (CLK), .D (signal_4955), .Q (signal_4956) ) ;
    buf_clk cell_2818 ( .C (CLK), .D (signal_4961), .Q (signal_4962) ) ;
    buf_clk cell_2824 ( .C (CLK), .D (signal_4967), .Q (signal_4968) ) ;
    buf_clk cell_2830 ( .C (CLK), .D (signal_4973), .Q (signal_4974) ) ;
    buf_clk cell_2836 ( .C (CLK), .D (signal_4979), .Q (signal_4980) ) ;
    buf_clk cell_2842 ( .C (CLK), .D (signal_4985), .Q (signal_4986) ) ;
    buf_clk cell_2848 ( .C (CLK), .D (signal_4991), .Q (signal_4992) ) ;
    buf_clk cell_2854 ( .C (CLK), .D (signal_4997), .Q (signal_4998) ) ;
    buf_clk cell_2860 ( .C (CLK), .D (signal_5003), .Q (signal_5004) ) ;
    buf_clk cell_2866 ( .C (CLK), .D (signal_5009), .Q (signal_5010) ) ;
    buf_clk cell_2934 ( .C (CLK), .D (signal_3899), .Q (signal_5078) ) ;
    buf_clk cell_2938 ( .C (CLK), .D (signal_3901), .Q (signal_5082) ) ;
    buf_clk cell_2972 ( .C (CLK), .D (signal_5115), .Q (signal_5116) ) ;
    buf_clk cell_2978 ( .C (CLK), .D (signal_5121), .Q (signal_5122) ) ;
    buf_clk cell_2982 ( .C (CLK), .D (signal_3871), .Q (signal_5126) ) ;
    buf_clk cell_2986 ( .C (CLK), .D (signal_3873), .Q (signal_5130) ) ;
    buf_clk cell_3014 ( .C (CLK), .D (signal_3879), .Q (signal_5158) ) ;
    buf_clk cell_3020 ( .C (CLK), .D (signal_3881), .Q (signal_5164) ) ;
    buf_clk cell_3056 ( .C (CLK), .D (signal_5199), .Q (signal_5200) ) ;
    buf_clk cell_3064 ( .C (CLK), .D (signal_5207), .Q (signal_5208) ) ;
    buf_clk cell_3194 ( .C (CLK), .D (signal_3907), .Q (signal_5338) ) ;
    buf_clk cell_3202 ( .C (CLK), .D (signal_3909), .Q (signal_5346) ) ;
    buf_clk cell_3448 ( .C (CLK), .D (signal_5591), .Q (signal_5592) ) ;
    buf_clk cell_3464 ( .C (CLK), .D (signal_5607), .Q (signal_5608) ) ;
    buf_clk cell_3488 ( .C (CLK), .D (signal_5631), .Q (signal_5632) ) ;
    buf_clk cell_3504 ( .C (CLK), .D (signal_5647), .Q (signal_5648) ) ;
    buf_clk cell_3528 ( .C (CLK), .D (signal_5671), .Q (signal_5672) ) ;
    buf_clk cell_3544 ( .C (CLK), .D (signal_5687), .Q (signal_5688) ) ;
    buf_clk cell_3560 ( .C (CLK), .D (signal_5703), .Q (signal_5704) ) ;
    buf_clk cell_3576 ( .C (CLK), .D (signal_5719), .Q (signal_5720) ) ;
    buf_clk cell_3636 ( .C (CLK), .D (signal_5779), .Q (signal_5780) ) ;
    buf_clk cell_3652 ( .C (CLK), .D (signal_5795), .Q (signal_5796) ) ;
    buf_clk cell_3668 ( .C (CLK), .D (signal_5811), .Q (signal_5812) ) ;
    buf_clk cell_3684 ( .C (CLK), .D (signal_5827), .Q (signal_5828) ) ;
    buf_clk cell_3700 ( .C (CLK), .D (signal_5843), .Q (signal_5844) ) ;
    buf_clk cell_3716 ( .C (CLK), .D (signal_5859), .Q (signal_5860) ) ;
    buf_clk cell_3732 ( .C (CLK), .D (signal_5875), .Q (signal_5876) ) ;
    buf_clk cell_3748 ( .C (CLK), .D (signal_5891), .Q (signal_5892) ) ;
    buf_clk cell_3764 ( .C (CLK), .D (signal_5907), .Q (signal_5908) ) ;
    buf_clk cell_3780 ( .C (CLK), .D (signal_5923), .Q (signal_5924) ) ;
    buf_clk cell_3888 ( .C (CLK), .D (signal_6031), .Q (signal_6032) ) ;
    buf_clk cell_3904 ( .C (CLK), .D (signal_6047), .Q (signal_6048) ) ;
    buf_clk cell_3920 ( .C (CLK), .D (signal_6063), .Q (signal_6064) ) ;
    buf_clk cell_3936 ( .C (CLK), .D (signal_6079), .Q (signal_6080) ) ;
    buf_clk cell_3952 ( .C (CLK), .D (signal_6095), .Q (signal_6096) ) ;
    buf_clk cell_3968 ( .C (CLK), .D (signal_6111), .Q (signal_6112) ) ;
    buf_clk cell_3984 ( .C (CLK), .D (signal_6127), .Q (signal_6128) ) ;
    buf_clk cell_4000 ( .C (CLK), .D (signal_6143), .Q (signal_6144) ) ;
    buf_clk cell_4016 ( .C (CLK), .D (signal_6159), .Q (signal_6160) ) ;
    buf_clk cell_4032 ( .C (CLK), .D (signal_6175), .Q (signal_6176) ) ;
    buf_clk cell_4048 ( .C (CLK), .D (signal_6191), .Q (signal_6192) ) ;
    buf_clk cell_4064 ( .C (CLK), .D (signal_6207), .Q (signal_6208) ) ;
    buf_clk cell_4080 ( .C (CLK), .D (signal_6223), .Q (signal_6224) ) ;
    buf_clk cell_4096 ( .C (CLK), .D (signal_6239), .Q (signal_6240) ) ;
    buf_clk cell_4180 ( .C (CLK), .D (signal_6323), .Q (signal_6324) ) ;
    buf_clk cell_4258 ( .C (CLK), .D (signal_3891), .Q (signal_6402) ) ;
    buf_clk cell_4272 ( .C (CLK), .D (signal_3893), .Q (signal_6416) ) ;
    buf_clk cell_4288 ( .C (CLK), .D (signal_6431), .Q (signal_6432) ) ;
    buf_clk cell_4304 ( .C (CLK), .D (signal_6447), .Q (signal_6448) ) ;
    buf_clk cell_4320 ( .C (CLK), .D (signal_6463), .Q (signal_6464) ) ;
    buf_clk cell_4336 ( .C (CLK), .D (signal_6479), .Q (signal_6480) ) ;
    buf_clk cell_4352 ( .C (CLK), .D (signal_6495), .Q (signal_6496) ) ;
    buf_clk cell_4368 ( .C (CLK), .D (signal_6511), .Q (signal_6512) ) ;
    buf_clk cell_4384 ( .C (CLK), .D (signal_6527), .Q (signal_6528) ) ;
    buf_clk cell_4400 ( .C (CLK), .D (signal_6543), .Q (signal_6544) ) ;
    buf_clk cell_4416 ( .C (CLK), .D (signal_6559), .Q (signal_6560) ) ;
    buf_clk cell_4432 ( .C (CLK), .D (signal_6575), .Q (signal_6576) ) ;
    buf_clk cell_4448 ( .C (CLK), .D (signal_6591), .Q (signal_6592) ) ;
    buf_clk cell_4464 ( .C (CLK), .D (signal_6607), .Q (signal_6608) ) ;
    buf_clk cell_4480 ( .C (CLK), .D (signal_6623), .Q (signal_6624) ) ;
    buf_clk cell_4496 ( .C (CLK), .D (signal_6639), .Q (signal_6640) ) ;
    buf_clk cell_4512 ( .C (CLK), .D (signal_6655), .Q (signal_6656) ) ;
    buf_clk cell_4528 ( .C (CLK), .D (signal_6671), .Q (signal_6672) ) ;
    buf_clk cell_4602 ( .C (CLK), .D (signal_3895), .Q (signal_6746) ) ;
    buf_clk cell_4616 ( .C (CLK), .D (signal_3897), .Q (signal_6760) ) ;
    buf_clk cell_4632 ( .C (CLK), .D (signal_6775), .Q (signal_6776) ) ;
    buf_clk cell_4648 ( .C (CLK), .D (signal_6791), .Q (signal_6792) ) ;
    buf_clk cell_4744 ( .C (CLK), .D (signal_6887), .Q (signal_6888) ) ;
    buf_clk cell_4760 ( .C (CLK), .D (signal_6903), .Q (signal_6904) ) ;
    buf_clk cell_4776 ( .C (CLK), .D (signal_6919), .Q (signal_6920) ) ;
    buf_clk cell_4792 ( .C (CLK), .D (signal_6935), .Q (signal_6936) ) ;
    buf_clk cell_4808 ( .C (CLK), .D (signal_6951), .Q (signal_6952) ) ;
    buf_clk cell_4824 ( .C (CLK), .D (signal_6967), .Q (signal_6968) ) ;
    buf_clk cell_4840 ( .C (CLK), .D (signal_6983), .Q (signal_6984) ) ;
    buf_clk cell_4856 ( .C (CLK), .D (signal_6999), .Q (signal_7000) ) ;
    buf_clk cell_4872 ( .C (CLK), .D (signal_7015), .Q (signal_7016) ) ;
    buf_clk cell_4888 ( .C (CLK), .D (signal_7031), .Q (signal_7032) ) ;
    buf_clk cell_4904 ( .C (CLK), .D (signal_7047), .Q (signal_7048) ) ;
    buf_clk cell_4920 ( .C (CLK), .D (signal_7063), .Q (signal_7064) ) ;
    buf_clk cell_4936 ( .C (CLK), .D (signal_7079), .Q (signal_7080) ) ;
    buf_clk cell_4952 ( .C (CLK), .D (signal_7095), .Q (signal_7096) ) ;
    buf_clk cell_4968 ( .C (CLK), .D (signal_7111), .Q (signal_7112) ) ;
    buf_clk cell_4984 ( .C (CLK), .D (signal_7127), .Q (signal_7128) ) ;
    buf_clk cell_5000 ( .C (CLK), .D (signal_7143), .Q (signal_7144) ) ;
    buf_clk cell_5016 ( .C (CLK), .D (signal_7159), .Q (signal_7160) ) ;
    buf_clk cell_5032 ( .C (CLK), .D (signal_7175), .Q (signal_7176) ) ;
    buf_clk cell_5048 ( .C (CLK), .D (signal_7191), .Q (signal_7192) ) ;
    buf_clk cell_5064 ( .C (CLK), .D (signal_7207), .Q (signal_7208) ) ;
    buf_clk cell_5080 ( .C (CLK), .D (signal_7223), .Q (signal_7224) ) ;
    buf_clk cell_5096 ( .C (CLK), .D (signal_7239), .Q (signal_7240) ) ;
    buf_clk cell_5112 ( .C (CLK), .D (signal_7255), .Q (signal_7256) ) ;
    buf_clk cell_5128 ( .C (CLK), .D (signal_7271), .Q (signal_7272) ) ;
    buf_clk cell_5144 ( .C (CLK), .D (signal_7287), .Q (signal_7288) ) ;
    buf_clk cell_5160 ( .C (CLK), .D (signal_7303), .Q (signal_7304) ) ;
    buf_clk cell_5176 ( .C (CLK), .D (signal_7319), .Q (signal_7320) ) ;
    buf_clk cell_5192 ( .C (CLK), .D (signal_7335), .Q (signal_7336) ) ;
    buf_clk cell_5208 ( .C (CLK), .D (signal_7351), .Q (signal_7352) ) ;
    buf_clk cell_5224 ( .C (CLK), .D (signal_7367), .Q (signal_7368) ) ;
    buf_clk cell_5240 ( .C (CLK), .D (signal_7383), .Q (signal_7384) ) ;
    buf_clk cell_5256 ( .C (CLK), .D (signal_7399), .Q (signal_7400) ) ;
    buf_clk cell_5272 ( .C (CLK), .D (signal_7415), .Q (signal_7416) ) ;
    buf_clk cell_5288 ( .C (CLK), .D (signal_7431), .Q (signal_7432) ) ;
    buf_clk cell_5304 ( .C (CLK), .D (signal_7447), .Q (signal_7448) ) ;
    buf_clk cell_5320 ( .C (CLK), .D (signal_7463), .Q (signal_7464) ) ;
    buf_clk cell_5336 ( .C (CLK), .D (signal_7479), .Q (signal_7480) ) ;
    buf_clk cell_5352 ( .C (CLK), .D (signal_7495), .Q (signal_7496) ) ;
    buf_clk cell_5368 ( .C (CLK), .D (signal_7511), .Q (signal_7512) ) ;
    buf_clk cell_5384 ( .C (CLK), .D (signal_7527), .Q (signal_7528) ) ;
    buf_clk cell_5400 ( .C (CLK), .D (signal_7543), .Q (signal_7544) ) ;
    buf_clk cell_5416 ( .C (CLK), .D (signal_7559), .Q (signal_7560) ) ;
    buf_clk cell_5432 ( .C (CLK), .D (signal_7575), .Q (signal_7576) ) ;
    buf_clk cell_5448 ( .C (CLK), .D (signal_7591), .Q (signal_7592) ) ;
    buf_clk cell_5464 ( .C (CLK), .D (signal_7607), .Q (signal_7608) ) ;
    buf_clk cell_5480 ( .C (CLK), .D (signal_7623), .Q (signal_7624) ) ;
    buf_clk cell_5496 ( .C (CLK), .D (signal_7639), .Q (signal_7640) ) ;
    buf_clk cell_5512 ( .C (CLK), .D (signal_7655), .Q (signal_7656) ) ;
    buf_clk cell_5528 ( .C (CLK), .D (signal_7671), .Q (signal_7672) ) ;
    buf_clk cell_5544 ( .C (CLK), .D (signal_7687), .Q (signal_7688) ) ;
    buf_clk cell_5560 ( .C (CLK), .D (signal_7703), .Q (signal_7704) ) ;
    buf_clk cell_5576 ( .C (CLK), .D (signal_7719), .Q (signal_7720) ) ;
    buf_clk cell_5592 ( .C (CLK), .D (signal_7735), .Q (signal_7736) ) ;
    buf_clk cell_5608 ( .C (CLK), .D (signal_7751), .Q (signal_7752) ) ;
    buf_clk cell_5624 ( .C (CLK), .D (signal_7767), .Q (signal_7768) ) ;
    buf_clk cell_5640 ( .C (CLK), .D (signal_7783), .Q (signal_7784) ) ;
    buf_clk cell_5656 ( .C (CLK), .D (signal_7799), .Q (signal_7800) ) ;
    buf_clk cell_5672 ( .C (CLK), .D (signal_7815), .Q (signal_7816) ) ;
    buf_clk cell_5688 ( .C (CLK), .D (signal_7831), .Q (signal_7832) ) ;
    buf_clk cell_5704 ( .C (CLK), .D (signal_7847), .Q (signal_7848) ) ;
    buf_clk cell_5720 ( .C (CLK), .D (signal_7863), .Q (signal_7864) ) ;
    buf_clk cell_5736 ( .C (CLK), .D (signal_7879), .Q (signal_7880) ) ;
    buf_clk cell_5752 ( .C (CLK), .D (signal_7895), .Q (signal_7896) ) ;
    buf_clk cell_5768 ( .C (CLK), .D (signal_7911), .Q (signal_7912) ) ;
    buf_clk cell_5784 ( .C (CLK), .D (signal_7927), .Q (signal_7928) ) ;
    buf_clk cell_5800 ( .C (CLK), .D (signal_7943), .Q (signal_7944) ) ;
    buf_clk cell_5816 ( .C (CLK), .D (signal_7959), .Q (signal_7960) ) ;
    buf_clk cell_5832 ( .C (CLK), .D (signal_7975), .Q (signal_7976) ) ;
    buf_clk cell_5848 ( .C (CLK), .D (signal_7991), .Q (signal_7992) ) ;
    buf_clk cell_5864 ( .C (CLK), .D (signal_8007), .Q (signal_8008) ) ;
    buf_clk cell_5880 ( .C (CLK), .D (signal_8023), .Q (signal_8024) ) ;
    buf_clk cell_5896 ( .C (CLK), .D (signal_8039), .Q (signal_8040) ) ;
    buf_clk cell_5912 ( .C (CLK), .D (signal_8055), .Q (signal_8056) ) ;
    buf_clk cell_5928 ( .C (CLK), .D (signal_8071), .Q (signal_8072) ) ;
    buf_clk cell_5944 ( .C (CLK), .D (signal_8087), .Q (signal_8088) ) ;
    buf_clk cell_5960 ( .C (CLK), .D (signal_8103), .Q (signal_8104) ) ;
    buf_clk cell_5976 ( .C (CLK), .D (signal_8119), .Q (signal_8120) ) ;
    buf_clk cell_5992 ( .C (CLK), .D (signal_8135), .Q (signal_8136) ) ;
    buf_clk cell_6008 ( .C (CLK), .D (signal_8151), .Q (signal_8152) ) ;
    buf_clk cell_6024 ( .C (CLK), .D (signal_8167), .Q (signal_8168) ) ;
    buf_clk cell_6040 ( .C (CLK), .D (signal_8183), .Q (signal_8184) ) ;
    buf_clk cell_6056 ( .C (CLK), .D (signal_8199), .Q (signal_8200) ) ;
    buf_clk cell_6072 ( .C (CLK), .D (signal_8215), .Q (signal_8216) ) ;
    buf_clk cell_6088 ( .C (CLK), .D (signal_8231), .Q (signal_8232) ) ;
    buf_clk cell_6104 ( .C (CLK), .D (signal_8247), .Q (signal_8248) ) ;
    buf_clk cell_6120 ( .C (CLK), .D (signal_8263), .Q (signal_8264) ) ;
    buf_clk cell_6136 ( .C (CLK), .D (signal_8279), .Q (signal_8280) ) ;
    buf_clk cell_6152 ( .C (CLK), .D (signal_8295), .Q (signal_8296) ) ;
    buf_clk cell_6168 ( .C (CLK), .D (signal_8311), .Q (signal_8312) ) ;
    buf_clk cell_6184 ( .C (CLK), .D (signal_8327), .Q (signal_8328) ) ;
    buf_clk cell_6200 ( .C (CLK), .D (signal_8343), .Q (signal_8344) ) ;
    buf_clk cell_6216 ( .C (CLK), .D (signal_8359), .Q (signal_8360) ) ;
    buf_clk cell_6232 ( .C (CLK), .D (signal_8375), .Q (signal_8376) ) ;
    buf_clk cell_6248 ( .C (CLK), .D (signal_8391), .Q (signal_8392) ) ;
    buf_clk cell_6264 ( .C (CLK), .D (signal_8407), .Q (signal_8408) ) ;
    buf_clk cell_6280 ( .C (CLK), .D (signal_8423), .Q (signal_8424) ) ;
    buf_clk cell_6296 ( .C (CLK), .D (signal_8439), .Q (signal_8440) ) ;
    buf_clk cell_6312 ( .C (CLK), .D (signal_8455), .Q (signal_8456) ) ;
    buf_clk cell_6328 ( .C (CLK), .D (signal_8471), .Q (signal_8472) ) ;
    buf_clk cell_6344 ( .C (CLK), .D (signal_8487), .Q (signal_8488) ) ;
    buf_clk cell_6360 ( .C (CLK), .D (signal_8503), .Q (signal_8504) ) ;
    buf_clk cell_6376 ( .C (CLK), .D (signal_8519), .Q (signal_8520) ) ;
    buf_clk cell_6392 ( .C (CLK), .D (signal_8535), .Q (signal_8536) ) ;
    buf_clk cell_7592 ( .C (CLK), .D (signal_9735), .Q (signal_9736) ) ;
    buf_clk cell_7608 ( .C (CLK), .D (signal_9751), .Q (signal_9752) ) ;
    buf_clk cell_7624 ( .C (CLK), .D (signal_9767), .Q (signal_9768) ) ;
    buf_clk cell_7640 ( .C (CLK), .D (signal_9783), .Q (signal_9784) ) ;
    buf_clk cell_7656 ( .C (CLK), .D (signal_9799), .Q (signal_9800) ) ;
    buf_clk cell_7672 ( .C (CLK), .D (signal_9815), .Q (signal_9816) ) ;
    buf_clk cell_7688 ( .C (CLK), .D (signal_9831), .Q (signal_9832) ) ;
    buf_clk cell_7704 ( .C (CLK), .D (signal_9847), .Q (signal_9848) ) ;
    buf_clk cell_7720 ( .C (CLK), .D (signal_9863), .Q (signal_9864) ) ;
    buf_clk cell_7736 ( .C (CLK), .D (signal_9879), .Q (signal_9880) ) ;
    buf_clk cell_7944 ( .C (CLK), .D (signal_10087), .Q (signal_10088) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1182 ( .s ({signal_3873, signal_3871}), .b ({1'b0, 1'b0}), .a ({signal_2266, signal_1328}), .clk (CLK), .r (Fresh[54]), .c ({signal_2320, signal_1382}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1183 ( .s ({signal_3873, signal_3871}), .b ({signal_2267, signal_1329}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[55]), .c ({signal_2321, signal_1383}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1184 ( .s ({signal_3873, signal_3871}), .b ({signal_2266, signal_1328}), .a ({signal_2267, signal_1329}), .clk (CLK), .r (Fresh[56]), .c ({signal_2322, signal_1384}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1185 ( .s ({signal_3877, signal_3875}), .b ({1'b0, 1'b0}), .a ({signal_2268, signal_1330}), .clk (CLK), .r (Fresh[57]), .c ({signal_2323, signal_1385}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1186 ( .s ({signal_3877, signal_3875}), .b ({signal_2269, signal_1331}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[58]), .c ({signal_2324, signal_1386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1187 ( .s ({signal_3877, signal_3875}), .b ({signal_2268, signal_1330}), .a ({signal_2269, signal_1331}), .clk (CLK), .r (Fresh[59]), .c ({signal_2325, signal_1387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1188 ( .s ({signal_3881, signal_3879}), .b ({1'b0, 1'b1}), .a ({signal_2270, signal_1332}), .clk (CLK), .r (Fresh[60]), .c ({signal_2326, signal_1388}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1189 ( .s ({signal_3881, signal_3879}), .b ({signal_2271, signal_1333}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[61]), .c ({signal_2327, signal_1389}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1190 ( .s ({signal_3881, signal_3879}), .b ({signal_2271, signal_1333}), .a ({signal_2270, signal_1332}), .clk (CLK), .r (Fresh[62]), .c ({signal_2328, signal_1390}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1191 ( .s ({signal_3885, signal_3883}), .b ({1'b0, 1'b0}), .a ({signal_2272, signal_1334}), .clk (CLK), .r (Fresh[63]), .c ({signal_2329, signal_1391}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1192 ( .s ({signal_3885, signal_3883}), .b ({signal_2273, signal_1335}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[64]), .c ({signal_2330, signal_1392}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1193 ( .s ({signal_3885, signal_3883}), .b ({signal_2272, signal_1334}), .a ({signal_2273, signal_1335}), .clk (CLK), .r (Fresh[65]), .c ({signal_2331, signal_1393}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1194 ( .s ({signal_3889, signal_3887}), .b ({1'b0, 1'b0}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[66]), .c ({signal_2332, signal_1394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1195 ( .s ({signal_3889, signal_3887}), .b ({signal_2275, signal_1337}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[67]), .c ({signal_2333, signal_1395}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1196 ( .s ({signal_3889, signal_3887}), .b ({signal_2274, signal_1336}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[68]), .c ({signal_2334, signal_1396}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1197 ( .s ({signal_3893, signal_3891}), .b ({1'b0, 1'b0}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[69]), .c ({signal_2335, signal_1397}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1198 ( .s ({signal_3893, signal_3891}), .b ({signal_2277, signal_1339}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[70]), .c ({signal_2336, signal_1398}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1199 ( .s ({signal_3893, signal_3891}), .b ({signal_2276, signal_1338}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[71]), .c ({signal_2337, signal_1399}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1200 ( .s ({signal_3897, signal_3895}), .b ({1'b0, 1'b0}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[72]), .c ({signal_2338, signal_1400}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1201 ( .s ({signal_3897, signal_3895}), .b ({signal_2279, signal_1341}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[73]), .c ({signal_2339, signal_1401}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1202 ( .s ({signal_3897, signal_3895}), .b ({signal_2278, signal_1340}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[74]), .c ({signal_2340, signal_1402}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1203 ( .s ({signal_3901, signal_3899}), .b ({1'b0, 1'b0}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[75]), .c ({signal_2341, signal_1403}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1204 ( .s ({signal_3901, signal_3899}), .b ({signal_2281, signal_1343}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[76]), .c ({signal_2342, signal_1404}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1205 ( .s ({signal_3901, signal_3899}), .b ({signal_2280, signal_1342}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[77]), .c ({signal_2343, signal_1405}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1206 ( .s ({signal_3905, signal_3903}), .b ({signal_2291, signal_1345}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[78]), .c ({signal_2380, signal_1406}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1207 ( .s ({signal_3905, signal_3903}), .b ({signal_2292, signal_1346}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[79]), .c ({signal_2381, signal_1407}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1208 ( .s ({signal_3909, signal_3907}), .b ({1'b0, 1'b0}), .a ({signal_2294, signal_1348}), .clk (CLK), .r (Fresh[80]), .c ({signal_2382, signal_1408}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1209 ( .s ({signal_3909, signal_3907}), .b ({1'b0, 1'b1}), .a ({signal_2294, signal_1348}), .clk (CLK), .r (Fresh[81]), .c ({signal_2383, signal_1409}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1210 ( .s ({signal_3913, signal_3911}), .b ({signal_2297, signal_1351}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[82]), .c ({signal_2384, signal_1410}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1211 ( .s ({signal_3913, signal_3911}), .b ({signal_2298, signal_1352}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[83]), .c ({signal_2385, signal_1411}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1212 ( .s ({signal_3917, signal_3915}), .b ({1'b0, 1'b1}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[84]), .c ({signal_2386, signal_1412}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1213 ( .s ({signal_3917, signal_3915}), .b ({1'b0, 1'b0}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[85]), .c ({signal_2387, signal_1413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1214 ( .s ({signal_3921, signal_3919}), .b ({signal_2302, signal_1357}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[86]), .c ({signal_2388, signal_1414}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1215 ( .s ({signal_3921, signal_3919}), .b ({1'b0, 1'b1}), .a ({signal_2303, signal_1358}), .clk (CLK), .r (Fresh[87]), .c ({signal_2389, signal_1415}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1216 ( .s ({signal_3925, signal_3923}), .b ({signal_2305, signal_1360}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[88]), .c ({signal_2390, signal_1416}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1217 ( .s ({signal_3925, signal_3923}), .b ({signal_2306, signal_1361}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[89]), .c ({signal_2391, signal_1417}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1218 ( .s ({signal_3929, signal_3927}), .b ({1'b0, 1'b0}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[90]), .c ({signal_2392, signal_1418}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1219 ( .s ({signal_3929, signal_3927}), .b ({1'b0, 1'b1}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[91]), .c ({signal_2393, signal_1419}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1220 ( .s ({signal_3933, signal_3931}), .b ({1'b0, 1'b0}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[92]), .c ({signal_2394, signal_1420}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1221 ( .s ({signal_3933, signal_3931}), .b ({1'b0, 1'b1}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[93]), .c ({signal_2395, signal_1421}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1222 ( .s ({signal_3889, signal_3887}), .b ({signal_2275, signal_1337}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[94]), .c ({signal_2344, signal_1422}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1223 ( .s ({signal_3889, signal_3887}), .b ({1'b0, 1'b1}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[95]), .c ({signal_2345, signal_1423}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1224 ( .s ({signal_3889, signal_3887}), .b ({signal_2274, signal_1336}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[96]), .c ({signal_2346, signal_1424}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1225 ( .s ({signal_3889, signal_3887}), .b ({1'b0, 1'b0}), .a ({signal_2275, signal_1337}), .clk (CLK), .r (Fresh[97]), .c ({signal_2347, signal_1425}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1226 ( .s ({signal_3889, signal_3887}), .b ({1'b0, 1'b1}), .a ({signal_2274, signal_1336}), .clk (CLK), .r (Fresh[98]), .c ({signal_2348, signal_1426}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1227 ( .s ({signal_3901, signal_3899}), .b ({1'b0, 1'b0}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[99]), .c ({signal_2349, signal_1427}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1228 ( .s ({signal_3901, signal_3899}), .b ({1'b0, 1'b1}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[100]), .c ({signal_2350, signal_1428}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1229 ( .s ({signal_3901, signal_3899}), .b ({signal_2281, signal_1343}), .a ({signal_2280, signal_1342}), .clk (CLK), .r (Fresh[101]), .c ({signal_2351, signal_1429}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1230 ( .s ({signal_3893, signal_3891}), .b ({signal_2277, signal_1339}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[102]), .c ({signal_2352, signal_1430}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1231 ( .s ({signal_3893, signal_3891}), .b ({1'b0, 1'b0}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[103]), .c ({signal_2353, signal_1431}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1232 ( .s ({signal_3893, signal_3891}), .b ({1'b0, 1'b1}), .a ({signal_2276, signal_1338}), .clk (CLK), .r (Fresh[104]), .c ({signal_2354, signal_1432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1233 ( .s ({signal_3929, signal_3927}), .b ({signal_2307, signal_1362}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[105]), .c ({signal_2396, signal_1433}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1234 ( .s ({signal_3929, signal_3927}), .b ({1'b0, 1'b0}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[106]), .c ({signal_2397, signal_1434}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1235 ( .s ({signal_3893, signal_3891}), .b ({1'b0, 1'b1}), .a ({signal_2277, signal_1339}), .clk (CLK), .r (Fresh[107]), .c ({signal_2355, signal_1435}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1236 ( .s ({signal_3893, signal_3891}), .b ({signal_2276, signal_1338}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[108]), .c ({signal_2356, signal_1436}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1237 ( .s ({signal_3885, signal_3883}), .b ({signal_2273, signal_1335}), .a ({signal_2272, signal_1334}), .clk (CLK), .r (Fresh[109]), .c ({signal_2357, signal_1437}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1238 ( .s ({signal_3885, signal_3883}), .b ({1'b0, 1'b1}), .a ({signal_2273, signal_1335}), .clk (CLK), .r (Fresh[110]), .c ({signal_2358, signal_1438}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1239 ( .s ({signal_3885, signal_3883}), .b ({signal_2272, signal_1334}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[111]), .c ({signal_2359, signal_1439}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1240 ( .s ({signal_3921, signal_3919}), .b ({signal_2302, signal_1357}), .a ({signal_2303, signal_1358}), .clk (CLK), .r (Fresh[112]), .c ({signal_2398, signal_1440}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1241 ( .s ({signal_3921, signal_3919}), .b ({1'b0, 1'b0}), .a ({signal_2302, signal_1357}), .clk (CLK), .r (Fresh[113]), .c ({signal_2399, signal_1441}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1242 ( .s ({signal_3897, signal_3895}), .b ({signal_2279, signal_1341}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[114]), .c ({signal_2360, signal_1442}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1243 ( .s ({signal_3937, signal_3935}), .b ({signal_2301, signal_1355}), .a ({signal_2315, signal_1373}), .clk (CLK), .r (Fresh[115]), .c ({signal_2400, signal_1443}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1244 ( .s ({signal_3937, signal_3935}), .b ({signal_2315, signal_1373}), .a ({signal_2301, signal_1355}), .clk (CLK), .r (Fresh[116]), .c ({signal_2401, signal_1444}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1245 ( .s ({signal_3917, signal_3915}), .b ({1'b0, 1'b0}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[117]), .c ({signal_2402, signal_1445}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1246 ( .s ({signal_3917, signal_3915}), .b ({signal_2300, signal_1354}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[118]), .c ({signal_2403, signal_1446}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1247 ( .s ({signal_3917, signal_3915}), .b ({signal_2299, signal_1353}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[119]), .c ({signal_2404, signal_1447}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1248 ( .s ({signal_3941, signal_3939}), .b ({signal_2291, signal_1345}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[120]), .c ({signal_2405, signal_1448}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1249 ( .s ({signal_3941, signal_3939}), .b ({signal_2292, signal_1346}), .a ({signal_2291, signal_1345}), .clk (CLK), .r (Fresh[121]), .c ({signal_2406, signal_1449}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1250 ( .s ({signal_3905, signal_3903}), .b ({signal_2299, signal_1353}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[122]), .c ({signal_2407, signal_1450}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1251 ( .s ({signal_3905, signal_3903}), .b ({signal_2300, signal_1354}), .a ({signal_2299, signal_1353}), .clk (CLK), .r (Fresh[123]), .c ({signal_2408, signal_1451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1252 ( .s ({signal_3881, signal_3879}), .b ({signal_2270, signal_1332}), .a ({signal_2271, signal_1333}), .clk (CLK), .r (Fresh[124]), .c ({signal_2361, signal_1452}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1253 ( .s ({signal_3881, signal_3879}), .b ({1'b0, 1'b0}), .a ({signal_2271, signal_1333}), .clk (CLK), .r (Fresh[125]), .c ({signal_2362, signal_1453}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1254 ( .s ({signal_3881, signal_3879}), .b ({signal_2270, signal_1332}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[126]), .c ({signal_2363, signal_1454}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1255 ( .s ({signal_3929, signal_3927}), .b ({signal_2308, signal_1363}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[127]), .c ({signal_2409, signal_1455}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1256 ( .s ({signal_3921, signal_3919}), .b ({signal_2303, signal_1358}), .a ({signal_2302, signal_1357}), .clk (CLK), .r (Fresh[128]), .c ({signal_2410, signal_1456}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1257 ( .s ({signal_3873, signal_3871}), .b ({1'b0, 1'b0}), .a ({signal_2267, signal_1329}), .clk (CLK), .r (Fresh[129]), .c ({signal_2364, signal_1457}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1258 ( .s ({signal_3873, signal_3871}), .b ({1'b0, 1'b1}), .a ({signal_2266, signal_1328}), .clk (CLK), .r (Fresh[130]), .c ({signal_2365, signal_1458}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1259 ( .s ({signal_3873, signal_3871}), .b ({signal_2267, signal_1329}), .a ({signal_2266, signal_1328}), .clk (CLK), .r (Fresh[131]), .c ({signal_2366, signal_1459}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1260 ( .s ({signal_3933, signal_3931}), .b ({signal_2310, signal_1365}), .a ({signal_2311, signal_1366}), .clk (CLK), .r (Fresh[132]), .c ({signal_2411, signal_1460}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1261 ( .s ({signal_3933, signal_3931}), .b ({1'b0, 1'b0}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[133]), .c ({signal_2412, signal_1461}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1262 ( .s ({signal_3921, signal_3919}), .b ({signal_2303, signal_1358}), .a ({1'b0, 1'b1}), .clk (CLK), .r (Fresh[134]), .c ({signal_2413, signal_1462}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1263 ( .s ({signal_3933, signal_3931}), .b ({signal_2311, signal_1366}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[135]), .c ({signal_2414, signal_1463}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1264 ( .s ({signal_3873, signal_3871}), .b ({1'b0, 1'b1}), .a ({signal_2267, signal_1329}), .clk (CLK), .r (Fresh[136]), .c ({signal_2367, signal_1464}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1265 ( .s ({signal_3873, signal_3871}), .b ({signal_2266, signal_1328}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[137]), .c ({signal_2368, signal_1465}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1266 ( .s ({signal_3925, signal_3923}), .b ({1'b0, 1'b0}), .a ({signal_2306, signal_1361}), .clk (CLK), .r (Fresh[138]), .c ({signal_2415, signal_1466}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1267 ( .s ({signal_3925, signal_3923}), .b ({1'b0, 1'b1}), .a ({signal_2305, signal_1360}), .clk (CLK), .r (Fresh[139]), .c ({signal_2416, signal_1467}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1268 ( .s ({signal_3877, signal_3875}), .b ({1'b0, 1'b0}), .a ({signal_2269, signal_1331}), .clk (CLK), .r (Fresh[140]), .c ({signal_2369, signal_1468}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1269 ( .s ({signal_3877, signal_3875}), .b ({1'b0, 1'b1}), .a ({signal_2268, signal_1330}), .clk (CLK), .r (Fresh[141]), .c ({signal_2370, signal_1469}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1270 ( .s ({signal_3877, signal_3875}), .b ({signal_2269, signal_1331}), .a ({signal_2268, signal_1330}), .clk (CLK), .r (Fresh[142]), .c ({signal_2371, signal_1470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1271 ( .s ({signal_3925, signal_3923}), .b ({signal_2305, signal_1360}), .a ({signal_2306, signal_1361}), .clk (CLK), .r (Fresh[143]), .c ({signal_2417, signal_1471}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1272 ( .s ({signal_3925, signal_3923}), .b ({signal_2306, signal_1361}), .a ({signal_2305, signal_1360}), .clk (CLK), .r (Fresh[144]), .c ({signal_2418, signal_1472}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1273 ( .s ({signal_3897, signal_3895}), .b ({1'b0, 1'b0}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[145]), .c ({signal_2372, signal_1473}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1274 ( .s ({signal_3897, signal_3895}), .b ({1'b0, 1'b1}), .a ({signal_2278, signal_1340}), .clk (CLK), .r (Fresh[146]), .c ({signal_2373, signal_1474}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1275 ( .s ({signal_3945, signal_3943}), .b ({signal_2297, signal_1351}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[147]), .c ({signal_2419, signal_1475}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1276 ( .s ({signal_3925, signal_3923}), .b ({signal_2297, signal_1351}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[148]), .c ({signal_2420, signal_1476}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1277 ( .s ({signal_3913, signal_3911}), .b ({signal_2298, signal_1352}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[149]), .c ({signal_2421, signal_1477}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1278 ( .s ({signal_3913, signal_3911}), .b ({signal_2297, signal_1351}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[150]), .c ({signal_2422, signal_1478}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1279 ( .s ({signal_3945, signal_3943}), .b ({signal_2296, signal_1350}), .a ({signal_2314, signal_1372}), .clk (CLK), .r (Fresh[151]), .c ({signal_2423, signal_1479}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1280 ( .s ({signal_3925, signal_3923}), .b ({signal_2296, signal_1350}), .a ({signal_2314, signal_1372}), .clk (CLK), .r (Fresh[152]), .c ({signal_2424, signal_1480}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1281 ( .s ({signal_3945, signal_3943}), .b ({signal_2298, signal_1352}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[153]), .c ({signal_2425, signal_1481}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1282 ( .s ({signal_3945, signal_3943}), .b ({signal_2314, signal_1372}), .a ({signal_2296, signal_1350}), .clk (CLK), .r (Fresh[154]), .c ({signal_2426, signal_1482}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1283 ( .s ({signal_3901, signal_3899}), .b ({1'b0, 1'b1}), .a ({signal_2281, signal_1343}), .clk (CLK), .r (Fresh[155]), .c ({signal_2374, signal_1483}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1284 ( .s ({signal_3901, signal_3899}), .b ({signal_2280, signal_1342}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[156]), .c ({signal_2375, signal_1484}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1285 ( .s ({signal_3905, signal_3903}), .b ({signal_2291, signal_1345}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[157]), .c ({signal_2427, signal_1485}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1286 ( .s ({signal_3905, signal_3903}), .b ({signal_2292, signal_1346}), .a ({signal_2291, signal_1345}), .clk (CLK), .r (Fresh[158]), .c ({signal_2428, signal_1486}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1287 ( .s ({signal_3905, signal_3903}), .b ({1'b0, 1'b1}), .a ({signal_2291, signal_1345}), .clk (CLK), .r (Fresh[159]), .c ({signal_2429, signal_1487}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1288 ( .s ({signal_3905, signal_3903}), .b ({1'b0, 1'b0}), .a ({signal_2292, signal_1346}), .clk (CLK), .r (Fresh[160]), .c ({signal_2430, signal_1488}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1289 ( .s ({signal_3909, signal_3907}), .b ({signal_2293, signal_1347}), .a ({signal_2294, signal_1348}), .clk (CLK), .r (Fresh[161]), .c ({signal_2431, signal_1489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1290 ( .s ({signal_3909, signal_3907}), .b ({1'b0, 1'b0}), .a ({signal_2293, signal_1347}), .clk (CLK), .r (Fresh[162]), .c ({signal_2432, signal_1490}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1291 ( .s ({signal_3949, signal_3947}), .b ({signal_2308, signal_1363}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[163]), .c ({signal_2433, signal_1491}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1292 ( .s ({signal_3929, signal_3927}), .b ({1'b0, 1'b1}), .a ({signal_2307, signal_1362}), .clk (CLK), .r (Fresh[164]), .c ({signal_2434, signal_1492}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1293 ( .s ({signal_3949, signal_3947}), .b ({signal_2309, signal_1364}), .a ({signal_2316, signal_1374}), .clk (CLK), .r (Fresh[165]), .c ({signal_2435, signal_1493}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1294 ( .s ({signal_3949, signal_3947}), .b ({signal_2307, signal_1362}), .a ({signal_2308, signal_1363}), .clk (CLK), .r (Fresh[166]), .c ({signal_2436, signal_1494}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1295 ( .s ({signal_3949, signal_3947}), .b ({signal_2316, signal_1374}), .a ({signal_2309, signal_1364}), .clk (CLK), .r (Fresh[167]), .c ({signal_2437, signal_1495}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1296 ( .s ({signal_3909, signal_3907}), .b ({signal_2294, signal_1348}), .a ({signal_2293, signal_1347}), .clk (CLK), .r (Fresh[168]), .c ({signal_2438, signal_1496}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1297 ( .s ({signal_3933, signal_3931}), .b ({1'b0, 1'b1}), .a ({signal_2310, signal_1365}), .clk (CLK), .r (Fresh[169]), .c ({signal_2439, signal_1497}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1298 ( .s ({signal_3897, signal_3895}), .b ({1'b0, 1'b1}), .a ({signal_2279, signal_1341}), .clk (CLK), .r (Fresh[170]), .c ({signal_2376, signal_1498}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1299 ( .s ({signal_3897, signal_3895}), .b ({signal_2278, signal_1340}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[171]), .c ({signal_2377, signal_1499}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1300 ( .s ({signal_3913, signal_3911}), .b ({1'b0, 1'b0}), .a ({signal_2298, signal_1352}), .clk (CLK), .r (Fresh[172]), .c ({signal_2440, signal_1500}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1301 ( .s ({signal_3913, signal_3911}), .b ({1'b0, 1'b1}), .a ({signal_2297, signal_1351}), .clk (CLK), .r (Fresh[173]), .c ({signal_2441, signal_1501}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1302 ( .s ({signal_3877, signal_3875}), .b ({1'b0, 1'b1}), .a ({signal_2269, signal_1331}), .clk (CLK), .r (Fresh[174]), .c ({signal_2378, signal_1502}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1303 ( .s ({signal_3877, signal_3875}), .b ({signal_2268, signal_1330}), .a ({1'b0, 1'b0}), .clk (CLK), .r (Fresh[175]), .c ({signal_2379, signal_1503}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1304 ( .s ({signal_3953, signal_3951}), .b ({signal_2299, signal_1353}), .a ({signal_2300, signal_1354}), .clk (CLK), .r (Fresh[176]), .c ({signal_2442, signal_1504}) ) ;
    buf_clk cell_1813 ( .C (CLK), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_1817 ( .C (CLK), .D (signal_3960), .Q (signal_3961) ) ;
    buf_clk cell_1819 ( .C (CLK), .D (signal_3962), .Q (signal_3963) ) ;
    buf_clk cell_1821 ( .C (CLK), .D (signal_3964), .Q (signal_3965) ) ;
    buf_clk cell_1825 ( .C (CLK), .D (signal_3968), .Q (signal_3969) ) ;
    buf_clk cell_1829 ( .C (CLK), .D (signal_3972), .Q (signal_3973) ) ;
    buf_clk cell_1831 ( .C (CLK), .D (signal_3974), .Q (signal_3975) ) ;
    buf_clk cell_1833 ( .C (CLK), .D (signal_3976), .Q (signal_3977) ) ;
    buf_clk cell_1837 ( .C (CLK), .D (signal_3980), .Q (signal_3981) ) ;
    buf_clk cell_1841 ( .C (CLK), .D (signal_3984), .Q (signal_3985) ) ;
    buf_clk cell_1843 ( .C (CLK), .D (signal_3986), .Q (signal_3987) ) ;
    buf_clk cell_1845 ( .C (CLK), .D (signal_3988), .Q (signal_3989) ) ;
    buf_clk cell_1849 ( .C (CLK), .D (signal_3992), .Q (signal_3993) ) ;
    buf_clk cell_1853 ( .C (CLK), .D (signal_3996), .Q (signal_3997) ) ;
    buf_clk cell_1855 ( .C (CLK), .D (signal_3998), .Q (signal_3999) ) ;
    buf_clk cell_1857 ( .C (CLK), .D (signal_4000), .Q (signal_4001) ) ;
    buf_clk cell_1861 ( .C (CLK), .D (signal_4004), .Q (signal_4005) ) ;
    buf_clk cell_1865 ( .C (CLK), .D (signal_4008), .Q (signal_4009) ) ;
    buf_clk cell_1867 ( .C (CLK), .D (signal_4010), .Q (signal_4011) ) ;
    buf_clk cell_1869 ( .C (CLK), .D (signal_4012), .Q (signal_4013) ) ;
    buf_clk cell_1873 ( .C (CLK), .D (signal_4016), .Q (signal_4017) ) ;
    buf_clk cell_1877 ( .C (CLK), .D (signal_4020), .Q (signal_4021) ) ;
    buf_clk cell_1879 ( .C (CLK), .D (signal_4022), .Q (signal_4023) ) ;
    buf_clk cell_1881 ( .C (CLK), .D (signal_4024), .Q (signal_4025) ) ;
    buf_clk cell_1885 ( .C (CLK), .D (signal_4028), .Q (signal_4029) ) ;
    buf_clk cell_1889 ( .C (CLK), .D (signal_4032), .Q (signal_4033) ) ;
    buf_clk cell_1891 ( .C (CLK), .D (signal_4034), .Q (signal_4035) ) ;
    buf_clk cell_1893 ( .C (CLK), .D (signal_4036), .Q (signal_4037) ) ;
    buf_clk cell_1897 ( .C (CLK), .D (signal_4040), .Q (signal_4041) ) ;
    buf_clk cell_1901 ( .C (CLK), .D (signal_4044), .Q (signal_4045) ) ;
    buf_clk cell_1903 ( .C (CLK), .D (signal_4046), .Q (signal_4047) ) ;
    buf_clk cell_1905 ( .C (CLK), .D (signal_4048), .Q (signal_4049) ) ;
    buf_clk cell_1909 ( .C (CLK), .D (signal_4052), .Q (signal_4053) ) ;
    buf_clk cell_1913 ( .C (CLK), .D (signal_4056), .Q (signal_4057) ) ;
    buf_clk cell_1915 ( .C (CLK), .D (signal_4058), .Q (signal_4059) ) ;
    buf_clk cell_1917 ( .C (CLK), .D (signal_4060), .Q (signal_4061) ) ;
    buf_clk cell_1919 ( .C (CLK), .D (signal_4062), .Q (signal_4063) ) ;
    buf_clk cell_1921 ( .C (CLK), .D (signal_4064), .Q (signal_4065) ) ;
    buf_clk cell_1925 ( .C (CLK), .D (signal_4068), .Q (signal_4069) ) ;
    buf_clk cell_1929 ( .C (CLK), .D (signal_4072), .Q (signal_4073) ) ;
    buf_clk cell_1931 ( .C (CLK), .D (signal_4074), .Q (signal_4075) ) ;
    buf_clk cell_1933 ( .C (CLK), .D (signal_4076), .Q (signal_4077) ) ;
    buf_clk cell_1935 ( .C (CLK), .D (signal_4078), .Q (signal_4079) ) ;
    buf_clk cell_1937 ( .C (CLK), .D (signal_4080), .Q (signal_4081) ) ;
    buf_clk cell_1941 ( .C (CLK), .D (signal_4084), .Q (signal_4085) ) ;
    buf_clk cell_1945 ( .C (CLK), .D (signal_4088), .Q (signal_4089) ) ;
    buf_clk cell_1947 ( .C (CLK), .D (signal_4090), .Q (signal_4091) ) ;
    buf_clk cell_1949 ( .C (CLK), .D (signal_4092), .Q (signal_4093) ) ;
    buf_clk cell_1951 ( .C (CLK), .D (signal_4094), .Q (signal_4095) ) ;
    buf_clk cell_1953 ( .C (CLK), .D (signal_4096), .Q (signal_4097) ) ;
    buf_clk cell_1955 ( .C (CLK), .D (signal_4098), .Q (signal_4099) ) ;
    buf_clk cell_1957 ( .C (CLK), .D (signal_4100), .Q (signal_4101) ) ;
    buf_clk cell_1959 ( .C (CLK), .D (signal_4102), .Q (signal_4103) ) ;
    buf_clk cell_1961 ( .C (CLK), .D (signal_4104), .Q (signal_4105) ) ;
    buf_clk cell_1963 ( .C (CLK), .D (signal_4106), .Q (signal_4107) ) ;
    buf_clk cell_1965 ( .C (CLK), .D (signal_4108), .Q (signal_4109) ) ;
    buf_clk cell_1969 ( .C (CLK), .D (signal_4112), .Q (signal_4113) ) ;
    buf_clk cell_1973 ( .C (CLK), .D (signal_4116), .Q (signal_4117) ) ;
    buf_clk cell_1975 ( .C (CLK), .D (signal_4118), .Q (signal_4119) ) ;
    buf_clk cell_1977 ( .C (CLK), .D (signal_4120), .Q (signal_4121) ) ;
    buf_clk cell_1979 ( .C (CLK), .D (signal_4122), .Q (signal_4123) ) ;
    buf_clk cell_1981 ( .C (CLK), .D (signal_4124), .Q (signal_4125) ) ;
    buf_clk cell_1985 ( .C (CLK), .D (signal_4128), .Q (signal_4129) ) ;
    buf_clk cell_1989 ( .C (CLK), .D (signal_4132), .Q (signal_4133) ) ;
    buf_clk cell_1991 ( .C (CLK), .D (signal_4134), .Q (signal_4135) ) ;
    buf_clk cell_1993 ( .C (CLK), .D (signal_4136), .Q (signal_4137) ) ;
    buf_clk cell_1995 ( .C (CLK), .D (signal_4138), .Q (signal_4139) ) ;
    buf_clk cell_1997 ( .C (CLK), .D (signal_4140), .Q (signal_4141) ) ;
    buf_clk cell_2001 ( .C (CLK), .D (signal_4144), .Q (signal_4145) ) ;
    buf_clk cell_2005 ( .C (CLK), .D (signal_4148), .Q (signal_4149) ) ;
    buf_clk cell_2007 ( .C (CLK), .D (signal_4150), .Q (signal_4151) ) ;
    buf_clk cell_2009 ( .C (CLK), .D (signal_4152), .Q (signal_4153) ) ;
    buf_clk cell_2011 ( .C (CLK), .D (signal_4154), .Q (signal_4155) ) ;
    buf_clk cell_2013 ( .C (CLK), .D (signal_4156), .Q (signal_4157) ) ;
    buf_clk cell_2017 ( .C (CLK), .D (signal_4160), .Q (signal_4161) ) ;
    buf_clk cell_2021 ( .C (CLK), .D (signal_4164), .Q (signal_4165) ) ;
    buf_clk cell_2023 ( .C (CLK), .D (signal_4166), .Q (signal_4167) ) ;
    buf_clk cell_2025 ( .C (CLK), .D (signal_4168), .Q (signal_4169) ) ;
    buf_clk cell_2027 ( .C (CLK), .D (signal_4170), .Q (signal_4171) ) ;
    buf_clk cell_2029 ( .C (CLK), .D (signal_4172), .Q (signal_4173) ) ;
    buf_clk cell_2031 ( .C (CLK), .D (signal_4174), .Q (signal_4175) ) ;
    buf_clk cell_2033 ( .C (CLK), .D (signal_4176), .Q (signal_4177) ) ;
    buf_clk cell_2035 ( .C (CLK), .D (signal_4178), .Q (signal_4179) ) ;
    buf_clk cell_2037 ( .C (CLK), .D (signal_4180), .Q (signal_4181) ) ;
    buf_clk cell_2039 ( .C (CLK), .D (signal_4182), .Q (signal_4183) ) ;
    buf_clk cell_2041 ( .C (CLK), .D (signal_4184), .Q (signal_4185) ) ;
    buf_clk cell_2043 ( .C (CLK), .D (signal_4186), .Q (signal_4187) ) ;
    buf_clk cell_2045 ( .C (CLK), .D (signal_4188), .Q (signal_4189) ) ;
    buf_clk cell_2047 ( .C (CLK), .D (signal_4190), .Q (signal_4191) ) ;
    buf_clk cell_2049 ( .C (CLK), .D (signal_4192), .Q (signal_4193) ) ;
    buf_clk cell_2051 ( .C (CLK), .D (signal_4194), .Q (signal_4195) ) ;
    buf_clk cell_2053 ( .C (CLK), .D (signal_4196), .Q (signal_4197) ) ;
    buf_clk cell_2055 ( .C (CLK), .D (signal_4198), .Q (signal_4199) ) ;
    buf_clk cell_2057 ( .C (CLK), .D (signal_4200), .Q (signal_4201) ) ;
    buf_clk cell_2059 ( .C (CLK), .D (signal_4202), .Q (signal_4203) ) ;
    buf_clk cell_2061 ( .C (CLK), .D (signal_4204), .Q (signal_4205) ) ;
    buf_clk cell_2063 ( .C (CLK), .D (signal_4206), .Q (signal_4207) ) ;
    buf_clk cell_2065 ( .C (CLK), .D (signal_4208), .Q (signal_4209) ) ;
    buf_clk cell_2067 ( .C (CLK), .D (signal_4210), .Q (signal_4211) ) ;
    buf_clk cell_2069 ( .C (CLK), .D (signal_4212), .Q (signal_4213) ) ;
    buf_clk cell_2071 ( .C (CLK), .D (signal_4214), .Q (signal_4215) ) ;
    buf_clk cell_2073 ( .C (CLK), .D (signal_4216), .Q (signal_4217) ) ;
    buf_clk cell_2075 ( .C (CLK), .D (signal_4218), .Q (signal_4219) ) ;
    buf_clk cell_2077 ( .C (CLK), .D (signal_4220), .Q (signal_4221) ) ;
    buf_clk cell_2079 ( .C (CLK), .D (signal_4222), .Q (signal_4223) ) ;
    buf_clk cell_2081 ( .C (CLK), .D (signal_4224), .Q (signal_4225) ) ;
    buf_clk cell_2083 ( .C (CLK), .D (signal_4226), .Q (signal_4227) ) ;
    buf_clk cell_2085 ( .C (CLK), .D (signal_4228), .Q (signal_4229) ) ;
    buf_clk cell_2087 ( .C (CLK), .D (signal_4230), .Q (signal_4231) ) ;
    buf_clk cell_2089 ( .C (CLK), .D (signal_4232), .Q (signal_4233) ) ;
    buf_clk cell_2091 ( .C (CLK), .D (signal_4234), .Q (signal_4235) ) ;
    buf_clk cell_2093 ( .C (CLK), .D (signal_4236), .Q (signal_4237) ) ;
    buf_clk cell_2095 ( .C (CLK), .D (signal_4238), .Q (signal_4239) ) ;
    buf_clk cell_2097 ( .C (CLK), .D (signal_4240), .Q (signal_4241) ) ;
    buf_clk cell_2099 ( .C (CLK), .D (signal_4242), .Q (signal_4243) ) ;
    buf_clk cell_2101 ( .C (CLK), .D (signal_4244), .Q (signal_4245) ) ;
    buf_clk cell_2103 ( .C (CLK), .D (signal_4246), .Q (signal_4247) ) ;
    buf_clk cell_2105 ( .C (CLK), .D (signal_4248), .Q (signal_4249) ) ;
    buf_clk cell_2107 ( .C (CLK), .D (signal_4250), .Q (signal_4251) ) ;
    buf_clk cell_2109 ( .C (CLK), .D (signal_4252), .Q (signal_4253) ) ;
    buf_clk cell_2111 ( .C (CLK), .D (signal_4254), .Q (signal_4255) ) ;
    buf_clk cell_2113 ( .C (CLK), .D (signal_4256), .Q (signal_4257) ) ;
    buf_clk cell_2115 ( .C (CLK), .D (signal_4258), .Q (signal_4259) ) ;
    buf_clk cell_2117 ( .C (CLK), .D (signal_4260), .Q (signal_4261) ) ;
    buf_clk cell_2119 ( .C (CLK), .D (signal_4262), .Q (signal_4263) ) ;
    buf_clk cell_2121 ( .C (CLK), .D (signal_4264), .Q (signal_4265) ) ;
    buf_clk cell_2123 ( .C (CLK), .D (signal_4266), .Q (signal_4267) ) ;
    buf_clk cell_2125 ( .C (CLK), .D (signal_4268), .Q (signal_4269) ) ;
    buf_clk cell_2127 ( .C (CLK), .D (signal_4270), .Q (signal_4271) ) ;
    buf_clk cell_2129 ( .C (CLK), .D (signal_4272), .Q (signal_4273) ) ;
    buf_clk cell_2131 ( .C (CLK), .D (signal_4274), .Q (signal_4275) ) ;
    buf_clk cell_2133 ( .C (CLK), .D (signal_4276), .Q (signal_4277) ) ;
    buf_clk cell_2135 ( .C (CLK), .D (signal_4278), .Q (signal_4279) ) ;
    buf_clk cell_2137 ( .C (CLK), .D (signal_4280), .Q (signal_4281) ) ;
    buf_clk cell_2139 ( .C (CLK), .D (signal_4282), .Q (signal_4283) ) ;
    buf_clk cell_2141 ( .C (CLK), .D (signal_4284), .Q (signal_4285) ) ;
    buf_clk cell_2143 ( .C (CLK), .D (signal_4286), .Q (signal_4287) ) ;
    buf_clk cell_2145 ( .C (CLK), .D (signal_4288), .Q (signal_4289) ) ;
    buf_clk cell_2147 ( .C (CLK), .D (signal_4290), .Q (signal_4291) ) ;
    buf_clk cell_2149 ( .C (CLK), .D (signal_4292), .Q (signal_4293) ) ;
    buf_clk cell_2151 ( .C (CLK), .D (signal_4294), .Q (signal_4295) ) ;
    buf_clk cell_2153 ( .C (CLK), .D (signal_4296), .Q (signal_4297) ) ;
    buf_clk cell_2155 ( .C (CLK), .D (signal_4298), .Q (signal_4299) ) ;
    buf_clk cell_2157 ( .C (CLK), .D (signal_4300), .Q (signal_4301) ) ;
    buf_clk cell_2161 ( .C (CLK), .D (signal_4304), .Q (signal_4305) ) ;
    buf_clk cell_2165 ( .C (CLK), .D (signal_4308), .Q (signal_4309) ) ;
    buf_clk cell_2167 ( .C (CLK), .D (signal_4310), .Q (signal_4311) ) ;
    buf_clk cell_2169 ( .C (CLK), .D (signal_4312), .Q (signal_4313) ) ;
    buf_clk cell_2171 ( .C (CLK), .D (signal_4314), .Q (signal_4315) ) ;
    buf_clk cell_2173 ( .C (CLK), .D (signal_4316), .Q (signal_4317) ) ;
    buf_clk cell_2177 ( .C (CLK), .D (signal_4320), .Q (signal_4321) ) ;
    buf_clk cell_2181 ( .C (CLK), .D (signal_4324), .Q (signal_4325) ) ;
    buf_clk cell_2183 ( .C (CLK), .D (signal_4326), .Q (signal_4327) ) ;
    buf_clk cell_2185 ( .C (CLK), .D (signal_4328), .Q (signal_4329) ) ;
    buf_clk cell_2187 ( .C (CLK), .D (signal_4330), .Q (signal_4331) ) ;
    buf_clk cell_2189 ( .C (CLK), .D (signal_4332), .Q (signal_4333) ) ;
    buf_clk cell_2193 ( .C (CLK), .D (signal_4336), .Q (signal_4337) ) ;
    buf_clk cell_2201 ( .C (CLK), .D (signal_4344), .Q (signal_4345) ) ;
    buf_clk cell_2209 ( .C (CLK), .D (signal_4352), .Q (signal_4353) ) ;
    buf_clk cell_2217 ( .C (CLK), .D (signal_4360), .Q (signal_4361) ) ;
    buf_clk cell_2225 ( .C (CLK), .D (signal_4368), .Q (signal_4369) ) ;
    buf_clk cell_2233 ( .C (CLK), .D (signal_4376), .Q (signal_4377) ) ;
    buf_clk cell_2241 ( .C (CLK), .D (signal_4384), .Q (signal_4385) ) ;
    buf_clk cell_2249 ( .C (CLK), .D (signal_4392), .Q (signal_4393) ) ;
    buf_clk cell_2257 ( .C (CLK), .D (signal_4400), .Q (signal_4401) ) ;
    buf_clk cell_2265 ( .C (CLK), .D (signal_4408), .Q (signal_4409) ) ;
    buf_clk cell_2281 ( .C (CLK), .D (signal_4424), .Q (signal_4425) ) ;
    buf_clk cell_2289 ( .C (CLK), .D (signal_4432), .Q (signal_4433) ) ;
    buf_clk cell_2313 ( .C (CLK), .D (signal_4456), .Q (signal_4457) ) ;
    buf_clk cell_2321 ( .C (CLK), .D (signal_4464), .Q (signal_4465) ) ;
    buf_clk cell_2329 ( .C (CLK), .D (signal_4472), .Q (signal_4473) ) ;
    buf_clk cell_2337 ( .C (CLK), .D (signal_4480), .Q (signal_4481) ) ;
    buf_clk cell_2353 ( .C (CLK), .D (signal_4496), .Q (signal_4497) ) ;
    buf_clk cell_2359 ( .C (CLK), .D (signal_4502), .Q (signal_4503) ) ;
    buf_clk cell_2365 ( .C (CLK), .D (signal_4508), .Q (signal_4509) ) ;
    buf_clk cell_2373 ( .C (CLK), .D (signal_4516), .Q (signal_4517) ) ;
    buf_clk cell_2381 ( .C (CLK), .D (signal_4524), .Q (signal_4525) ) ;
    buf_clk cell_2389 ( .C (CLK), .D (signal_4532), .Q (signal_4533) ) ;
    buf_clk cell_2397 ( .C (CLK), .D (signal_4540), .Q (signal_4541) ) ;
    buf_clk cell_2405 ( .C (CLK), .D (signal_4548), .Q (signal_4549) ) ;
    buf_clk cell_2413 ( .C (CLK), .D (signal_4556), .Q (signal_4557) ) ;
    buf_clk cell_2421 ( .C (CLK), .D (signal_4564), .Q (signal_4565) ) ;
    buf_clk cell_2429 ( .C (CLK), .D (signal_4572), .Q (signal_4573) ) ;
    buf_clk cell_2437 ( .C (CLK), .D (signal_4580), .Q (signal_4581) ) ;
    buf_clk cell_2445 ( .C (CLK), .D (signal_4588), .Q (signal_4589) ) ;
    buf_clk cell_2453 ( .C (CLK), .D (signal_4596), .Q (signal_4597) ) ;
    buf_clk cell_2461 ( .C (CLK), .D (signal_4604), .Q (signal_4605) ) ;
    buf_clk cell_2469 ( .C (CLK), .D (signal_4612), .Q (signal_4613) ) ;
    buf_clk cell_2477 ( .C (CLK), .D (signal_4620), .Q (signal_4621) ) ;
    buf_clk cell_2485 ( .C (CLK), .D (signal_4628), .Q (signal_4629) ) ;
    buf_clk cell_2493 ( .C (CLK), .D (signal_4636), .Q (signal_4637) ) ;
    buf_clk cell_2501 ( .C (CLK), .D (signal_4644), .Q (signal_4645) ) ;
    buf_clk cell_2509 ( .C (CLK), .D (signal_4652), .Q (signal_4653) ) ;
    buf_clk cell_2517 ( .C (CLK), .D (signal_4660), .Q (signal_4661) ) ;
    buf_clk cell_2525 ( .C (CLK), .D (signal_4668), .Q (signal_4669) ) ;
    buf_clk cell_2533 ( .C (CLK), .D (signal_4676), .Q (signal_4677) ) ;
    buf_clk cell_2541 ( .C (CLK), .D (signal_4684), .Q (signal_4685) ) ;
    buf_clk cell_2549 ( .C (CLK), .D (signal_4692), .Q (signal_4693) ) ;
    buf_clk cell_2557 ( .C (CLK), .D (signal_4700), .Q (signal_4701) ) ;
    buf_clk cell_2565 ( .C (CLK), .D (signal_4708), .Q (signal_4709) ) ;
    buf_clk cell_2589 ( .C (CLK), .D (signal_4732), .Q (signal_4733) ) ;
    buf_clk cell_2597 ( .C (CLK), .D (signal_4740), .Q (signal_4741) ) ;
    buf_clk cell_2605 ( .C (CLK), .D (signal_4748), .Q (signal_4749) ) ;
    buf_clk cell_2613 ( .C (CLK), .D (signal_4756), .Q (signal_4757) ) ;
    buf_clk cell_2627 ( .C (CLK), .D (signal_4770), .Q (signal_4771) ) ;
    buf_clk cell_2633 ( .C (CLK), .D (signal_4776), .Q (signal_4777) ) ;
    buf_clk cell_2641 ( .C (CLK), .D (signal_4784), .Q (signal_4785) ) ;
    buf_clk cell_2649 ( .C (CLK), .D (signal_4792), .Q (signal_4793) ) ;
    buf_clk cell_2657 ( .C (CLK), .D (signal_4800), .Q (signal_4801) ) ;
    buf_clk cell_2665 ( .C (CLK), .D (signal_4808), .Q (signal_4809) ) ;
    buf_clk cell_2671 ( .C (CLK), .D (signal_4814), .Q (signal_4815) ) ;
    buf_clk cell_2677 ( .C (CLK), .D (signal_4820), .Q (signal_4821) ) ;
    buf_clk cell_2693 ( .C (CLK), .D (signal_4836), .Q (signal_4837) ) ;
    buf_clk cell_2701 ( .C (CLK), .D (signal_4844), .Q (signal_4845) ) ;
    buf_clk cell_2709 ( .C (CLK), .D (signal_4852), .Q (signal_4853) ) ;
    buf_clk cell_2717 ( .C (CLK), .D (signal_4860), .Q (signal_4861) ) ;
    buf_clk cell_2725 ( .C (CLK), .D (signal_4868), .Q (signal_4869) ) ;
    buf_clk cell_2733 ( .C (CLK), .D (signal_4876), .Q (signal_4877) ) ;
    buf_clk cell_2741 ( .C (CLK), .D (signal_4884), .Q (signal_4885) ) ;
    buf_clk cell_2749 ( .C (CLK), .D (signal_4892), .Q (signal_4893) ) ;
    buf_clk cell_2757 ( .C (CLK), .D (signal_4900), .Q (signal_4901) ) ;
    buf_clk cell_2765 ( .C (CLK), .D (signal_4908), .Q (signal_4909) ) ;
    buf_clk cell_2773 ( .C (CLK), .D (signal_4916), .Q (signal_4917) ) ;
    buf_clk cell_2781 ( .C (CLK), .D (signal_4924), .Q (signal_4925) ) ;
    buf_clk cell_2789 ( .C (CLK), .D (signal_4932), .Q (signal_4933) ) ;
    buf_clk cell_2795 ( .C (CLK), .D (signal_4938), .Q (signal_4939) ) ;
    buf_clk cell_2801 ( .C (CLK), .D (signal_4944), .Q (signal_4945) ) ;
    buf_clk cell_2807 ( .C (CLK), .D (signal_4950), .Q (signal_4951) ) ;
    buf_clk cell_2813 ( .C (CLK), .D (signal_4956), .Q (signal_4957) ) ;
    buf_clk cell_2819 ( .C (CLK), .D (signal_4962), .Q (signal_4963) ) ;
    buf_clk cell_2825 ( .C (CLK), .D (signal_4968), .Q (signal_4969) ) ;
    buf_clk cell_2831 ( .C (CLK), .D (signal_4974), .Q (signal_4975) ) ;
    buf_clk cell_2837 ( .C (CLK), .D (signal_4980), .Q (signal_4981) ) ;
    buf_clk cell_2843 ( .C (CLK), .D (signal_4986), .Q (signal_4987) ) ;
    buf_clk cell_2849 ( .C (CLK), .D (signal_4992), .Q (signal_4993) ) ;
    buf_clk cell_2855 ( .C (CLK), .D (signal_4998), .Q (signal_4999) ) ;
    buf_clk cell_2861 ( .C (CLK), .D (signal_5004), .Q (signal_5005) ) ;
    buf_clk cell_2867 ( .C (CLK), .D (signal_5010), .Q (signal_5011) ) ;
    buf_clk cell_2935 ( .C (CLK), .D (signal_5078), .Q (signal_5079) ) ;
    buf_clk cell_2939 ( .C (CLK), .D (signal_5082), .Q (signal_5083) ) ;
    buf_clk cell_2973 ( .C (CLK), .D (signal_5116), .Q (signal_5117) ) ;
    buf_clk cell_2979 ( .C (CLK), .D (signal_5122), .Q (signal_5123) ) ;
    buf_clk cell_2983 ( .C (CLK), .D (signal_5126), .Q (signal_5127) ) ;
    buf_clk cell_2987 ( .C (CLK), .D (signal_5130), .Q (signal_5131) ) ;
    buf_clk cell_3015 ( .C (CLK), .D (signal_5158), .Q (signal_5159) ) ;
    buf_clk cell_3021 ( .C (CLK), .D (signal_5164), .Q (signal_5165) ) ;
    buf_clk cell_3057 ( .C (CLK), .D (signal_5200), .Q (signal_5201) ) ;
    buf_clk cell_3065 ( .C (CLK), .D (signal_5208), .Q (signal_5209) ) ;
    buf_clk cell_3195 ( .C (CLK), .D (signal_5338), .Q (signal_5339) ) ;
    buf_clk cell_3203 ( .C (CLK), .D (signal_5346), .Q (signal_5347) ) ;
    buf_clk cell_3449 ( .C (CLK), .D (signal_5592), .Q (signal_5593) ) ;
    buf_clk cell_3465 ( .C (CLK), .D (signal_5608), .Q (signal_5609) ) ;
    buf_clk cell_3489 ( .C (CLK), .D (signal_5632), .Q (signal_5633) ) ;
    buf_clk cell_3505 ( .C (CLK), .D (signal_5648), .Q (signal_5649) ) ;
    buf_clk cell_3529 ( .C (CLK), .D (signal_5672), .Q (signal_5673) ) ;
    buf_clk cell_3545 ( .C (CLK), .D (signal_5688), .Q (signal_5689) ) ;
    buf_clk cell_3561 ( .C (CLK), .D (signal_5704), .Q (signal_5705) ) ;
    buf_clk cell_3577 ( .C (CLK), .D (signal_5720), .Q (signal_5721) ) ;
    buf_clk cell_3637 ( .C (CLK), .D (signal_5780), .Q (signal_5781) ) ;
    buf_clk cell_3653 ( .C (CLK), .D (signal_5796), .Q (signal_5797) ) ;
    buf_clk cell_3669 ( .C (CLK), .D (signal_5812), .Q (signal_5813) ) ;
    buf_clk cell_3685 ( .C (CLK), .D (signal_5828), .Q (signal_5829) ) ;
    buf_clk cell_3701 ( .C (CLK), .D (signal_5844), .Q (signal_5845) ) ;
    buf_clk cell_3717 ( .C (CLK), .D (signal_5860), .Q (signal_5861) ) ;
    buf_clk cell_3733 ( .C (CLK), .D (signal_5876), .Q (signal_5877) ) ;
    buf_clk cell_3749 ( .C (CLK), .D (signal_5892), .Q (signal_5893) ) ;
    buf_clk cell_3765 ( .C (CLK), .D (signal_5908), .Q (signal_5909) ) ;
    buf_clk cell_3781 ( .C (CLK), .D (signal_5924), .Q (signal_5925) ) ;
    buf_clk cell_3889 ( .C (CLK), .D (signal_6032), .Q (signal_6033) ) ;
    buf_clk cell_3905 ( .C (CLK), .D (signal_6048), .Q (signal_6049) ) ;
    buf_clk cell_3921 ( .C (CLK), .D (signal_6064), .Q (signal_6065) ) ;
    buf_clk cell_3937 ( .C (CLK), .D (signal_6080), .Q (signal_6081) ) ;
    buf_clk cell_3953 ( .C (CLK), .D (signal_6096), .Q (signal_6097) ) ;
    buf_clk cell_3969 ( .C (CLK), .D (signal_6112), .Q (signal_6113) ) ;
    buf_clk cell_3985 ( .C (CLK), .D (signal_6128), .Q (signal_6129) ) ;
    buf_clk cell_4001 ( .C (CLK), .D (signal_6144), .Q (signal_6145) ) ;
    buf_clk cell_4017 ( .C (CLK), .D (signal_6160), .Q (signal_6161) ) ;
    buf_clk cell_4033 ( .C (CLK), .D (signal_6176), .Q (signal_6177) ) ;
    buf_clk cell_4049 ( .C (CLK), .D (signal_6192), .Q (signal_6193) ) ;
    buf_clk cell_4065 ( .C (CLK), .D (signal_6208), .Q (signal_6209) ) ;
    buf_clk cell_4081 ( .C (CLK), .D (signal_6224), .Q (signal_6225) ) ;
    buf_clk cell_4097 ( .C (CLK), .D (signal_6240), .Q (signal_6241) ) ;
    buf_clk cell_4181 ( .C (CLK), .D (signal_6324), .Q (signal_6325) ) ;
    buf_clk cell_4259 ( .C (CLK), .D (signal_6402), .Q (signal_6403) ) ;
    buf_clk cell_4273 ( .C (CLK), .D (signal_6416), .Q (signal_6417) ) ;
    buf_clk cell_4289 ( .C (CLK), .D (signal_6432), .Q (signal_6433) ) ;
    buf_clk cell_4305 ( .C (CLK), .D (signal_6448), .Q (signal_6449) ) ;
    buf_clk cell_4321 ( .C (CLK), .D (signal_6464), .Q (signal_6465) ) ;
    buf_clk cell_4337 ( .C (CLK), .D (signal_6480), .Q (signal_6481) ) ;
    buf_clk cell_4353 ( .C (CLK), .D (signal_6496), .Q (signal_6497) ) ;
    buf_clk cell_4369 ( .C (CLK), .D (signal_6512), .Q (signal_6513) ) ;
    buf_clk cell_4385 ( .C (CLK), .D (signal_6528), .Q (signal_6529) ) ;
    buf_clk cell_4401 ( .C (CLK), .D (signal_6544), .Q (signal_6545) ) ;
    buf_clk cell_4417 ( .C (CLK), .D (signal_6560), .Q (signal_6561) ) ;
    buf_clk cell_4433 ( .C (CLK), .D (signal_6576), .Q (signal_6577) ) ;
    buf_clk cell_4449 ( .C (CLK), .D (signal_6592), .Q (signal_6593) ) ;
    buf_clk cell_4465 ( .C (CLK), .D (signal_6608), .Q (signal_6609) ) ;
    buf_clk cell_4481 ( .C (CLK), .D (signal_6624), .Q (signal_6625) ) ;
    buf_clk cell_4497 ( .C (CLK), .D (signal_6640), .Q (signal_6641) ) ;
    buf_clk cell_4513 ( .C (CLK), .D (signal_6656), .Q (signal_6657) ) ;
    buf_clk cell_4529 ( .C (CLK), .D (signal_6672), .Q (signal_6673) ) ;
    buf_clk cell_4603 ( .C (CLK), .D (signal_6746), .Q (signal_6747) ) ;
    buf_clk cell_4617 ( .C (CLK), .D (signal_6760), .Q (signal_6761) ) ;
    buf_clk cell_4633 ( .C (CLK), .D (signal_6776), .Q (signal_6777) ) ;
    buf_clk cell_4649 ( .C (CLK), .D (signal_6792), .Q (signal_6793) ) ;
    buf_clk cell_4745 ( .C (CLK), .D (signal_6888), .Q (signal_6889) ) ;
    buf_clk cell_4761 ( .C (CLK), .D (signal_6904), .Q (signal_6905) ) ;
    buf_clk cell_4777 ( .C (CLK), .D (signal_6920), .Q (signal_6921) ) ;
    buf_clk cell_4793 ( .C (CLK), .D (signal_6936), .Q (signal_6937) ) ;
    buf_clk cell_4809 ( .C (CLK), .D (signal_6952), .Q (signal_6953) ) ;
    buf_clk cell_4825 ( .C (CLK), .D (signal_6968), .Q (signal_6969) ) ;
    buf_clk cell_4841 ( .C (CLK), .D (signal_6984), .Q (signal_6985) ) ;
    buf_clk cell_4857 ( .C (CLK), .D (signal_7000), .Q (signal_7001) ) ;
    buf_clk cell_4873 ( .C (CLK), .D (signal_7016), .Q (signal_7017) ) ;
    buf_clk cell_4889 ( .C (CLK), .D (signal_7032), .Q (signal_7033) ) ;
    buf_clk cell_4905 ( .C (CLK), .D (signal_7048), .Q (signal_7049) ) ;
    buf_clk cell_4921 ( .C (CLK), .D (signal_7064), .Q (signal_7065) ) ;
    buf_clk cell_4937 ( .C (CLK), .D (signal_7080), .Q (signal_7081) ) ;
    buf_clk cell_4953 ( .C (CLK), .D (signal_7096), .Q (signal_7097) ) ;
    buf_clk cell_4969 ( .C (CLK), .D (signal_7112), .Q (signal_7113) ) ;
    buf_clk cell_4985 ( .C (CLK), .D (signal_7128), .Q (signal_7129) ) ;
    buf_clk cell_5001 ( .C (CLK), .D (signal_7144), .Q (signal_7145) ) ;
    buf_clk cell_5017 ( .C (CLK), .D (signal_7160), .Q (signal_7161) ) ;
    buf_clk cell_5033 ( .C (CLK), .D (signal_7176), .Q (signal_7177) ) ;
    buf_clk cell_5049 ( .C (CLK), .D (signal_7192), .Q (signal_7193) ) ;
    buf_clk cell_5065 ( .C (CLK), .D (signal_7208), .Q (signal_7209) ) ;
    buf_clk cell_5081 ( .C (CLK), .D (signal_7224), .Q (signal_7225) ) ;
    buf_clk cell_5097 ( .C (CLK), .D (signal_7240), .Q (signal_7241) ) ;
    buf_clk cell_5113 ( .C (CLK), .D (signal_7256), .Q (signal_7257) ) ;
    buf_clk cell_5129 ( .C (CLK), .D (signal_7272), .Q (signal_7273) ) ;
    buf_clk cell_5145 ( .C (CLK), .D (signal_7288), .Q (signal_7289) ) ;
    buf_clk cell_5161 ( .C (CLK), .D (signal_7304), .Q (signal_7305) ) ;
    buf_clk cell_5177 ( .C (CLK), .D (signal_7320), .Q (signal_7321) ) ;
    buf_clk cell_5193 ( .C (CLK), .D (signal_7336), .Q (signal_7337) ) ;
    buf_clk cell_5209 ( .C (CLK), .D (signal_7352), .Q (signal_7353) ) ;
    buf_clk cell_5225 ( .C (CLK), .D (signal_7368), .Q (signal_7369) ) ;
    buf_clk cell_5241 ( .C (CLK), .D (signal_7384), .Q (signal_7385) ) ;
    buf_clk cell_5257 ( .C (CLK), .D (signal_7400), .Q (signal_7401) ) ;
    buf_clk cell_5273 ( .C (CLK), .D (signal_7416), .Q (signal_7417) ) ;
    buf_clk cell_5289 ( .C (CLK), .D (signal_7432), .Q (signal_7433) ) ;
    buf_clk cell_5305 ( .C (CLK), .D (signal_7448), .Q (signal_7449) ) ;
    buf_clk cell_5321 ( .C (CLK), .D (signal_7464), .Q (signal_7465) ) ;
    buf_clk cell_5337 ( .C (CLK), .D (signal_7480), .Q (signal_7481) ) ;
    buf_clk cell_5353 ( .C (CLK), .D (signal_7496), .Q (signal_7497) ) ;
    buf_clk cell_5369 ( .C (CLK), .D (signal_7512), .Q (signal_7513) ) ;
    buf_clk cell_5385 ( .C (CLK), .D (signal_7528), .Q (signal_7529) ) ;
    buf_clk cell_5401 ( .C (CLK), .D (signal_7544), .Q (signal_7545) ) ;
    buf_clk cell_5417 ( .C (CLK), .D (signal_7560), .Q (signal_7561) ) ;
    buf_clk cell_5433 ( .C (CLK), .D (signal_7576), .Q (signal_7577) ) ;
    buf_clk cell_5449 ( .C (CLK), .D (signal_7592), .Q (signal_7593) ) ;
    buf_clk cell_5465 ( .C (CLK), .D (signal_7608), .Q (signal_7609) ) ;
    buf_clk cell_5481 ( .C (CLK), .D (signal_7624), .Q (signal_7625) ) ;
    buf_clk cell_5497 ( .C (CLK), .D (signal_7640), .Q (signal_7641) ) ;
    buf_clk cell_5513 ( .C (CLK), .D (signal_7656), .Q (signal_7657) ) ;
    buf_clk cell_5529 ( .C (CLK), .D (signal_7672), .Q (signal_7673) ) ;
    buf_clk cell_5545 ( .C (CLK), .D (signal_7688), .Q (signal_7689) ) ;
    buf_clk cell_5561 ( .C (CLK), .D (signal_7704), .Q (signal_7705) ) ;
    buf_clk cell_5577 ( .C (CLK), .D (signal_7720), .Q (signal_7721) ) ;
    buf_clk cell_5593 ( .C (CLK), .D (signal_7736), .Q (signal_7737) ) ;
    buf_clk cell_5609 ( .C (CLK), .D (signal_7752), .Q (signal_7753) ) ;
    buf_clk cell_5625 ( .C (CLK), .D (signal_7768), .Q (signal_7769) ) ;
    buf_clk cell_5641 ( .C (CLK), .D (signal_7784), .Q (signal_7785) ) ;
    buf_clk cell_5657 ( .C (CLK), .D (signal_7800), .Q (signal_7801) ) ;
    buf_clk cell_5673 ( .C (CLK), .D (signal_7816), .Q (signal_7817) ) ;
    buf_clk cell_5689 ( .C (CLK), .D (signal_7832), .Q (signal_7833) ) ;
    buf_clk cell_5705 ( .C (CLK), .D (signal_7848), .Q (signal_7849) ) ;
    buf_clk cell_5721 ( .C (CLK), .D (signal_7864), .Q (signal_7865) ) ;
    buf_clk cell_5737 ( .C (CLK), .D (signal_7880), .Q (signal_7881) ) ;
    buf_clk cell_5753 ( .C (CLK), .D (signal_7896), .Q (signal_7897) ) ;
    buf_clk cell_5769 ( .C (CLK), .D (signal_7912), .Q (signal_7913) ) ;
    buf_clk cell_5785 ( .C (CLK), .D (signal_7928), .Q (signal_7929) ) ;
    buf_clk cell_5801 ( .C (CLK), .D (signal_7944), .Q (signal_7945) ) ;
    buf_clk cell_5817 ( .C (CLK), .D (signal_7960), .Q (signal_7961) ) ;
    buf_clk cell_5833 ( .C (CLK), .D (signal_7976), .Q (signal_7977) ) ;
    buf_clk cell_5849 ( .C (CLK), .D (signal_7992), .Q (signal_7993) ) ;
    buf_clk cell_5865 ( .C (CLK), .D (signal_8008), .Q (signal_8009) ) ;
    buf_clk cell_5881 ( .C (CLK), .D (signal_8024), .Q (signal_8025) ) ;
    buf_clk cell_5897 ( .C (CLK), .D (signal_8040), .Q (signal_8041) ) ;
    buf_clk cell_5913 ( .C (CLK), .D (signal_8056), .Q (signal_8057) ) ;
    buf_clk cell_5929 ( .C (CLK), .D (signal_8072), .Q (signal_8073) ) ;
    buf_clk cell_5945 ( .C (CLK), .D (signal_8088), .Q (signal_8089) ) ;
    buf_clk cell_5961 ( .C (CLK), .D (signal_8104), .Q (signal_8105) ) ;
    buf_clk cell_5977 ( .C (CLK), .D (signal_8120), .Q (signal_8121) ) ;
    buf_clk cell_5993 ( .C (CLK), .D (signal_8136), .Q (signal_8137) ) ;
    buf_clk cell_6009 ( .C (CLK), .D (signal_8152), .Q (signal_8153) ) ;
    buf_clk cell_6025 ( .C (CLK), .D (signal_8168), .Q (signal_8169) ) ;
    buf_clk cell_6041 ( .C (CLK), .D (signal_8184), .Q (signal_8185) ) ;
    buf_clk cell_6057 ( .C (CLK), .D (signal_8200), .Q (signal_8201) ) ;
    buf_clk cell_6073 ( .C (CLK), .D (signal_8216), .Q (signal_8217) ) ;
    buf_clk cell_6089 ( .C (CLK), .D (signal_8232), .Q (signal_8233) ) ;
    buf_clk cell_6105 ( .C (CLK), .D (signal_8248), .Q (signal_8249) ) ;
    buf_clk cell_6121 ( .C (CLK), .D (signal_8264), .Q (signal_8265) ) ;
    buf_clk cell_6137 ( .C (CLK), .D (signal_8280), .Q (signal_8281) ) ;
    buf_clk cell_6153 ( .C (CLK), .D (signal_8296), .Q (signal_8297) ) ;
    buf_clk cell_6169 ( .C (CLK), .D (signal_8312), .Q (signal_8313) ) ;
    buf_clk cell_6185 ( .C (CLK), .D (signal_8328), .Q (signal_8329) ) ;
    buf_clk cell_6201 ( .C (CLK), .D (signal_8344), .Q (signal_8345) ) ;
    buf_clk cell_6217 ( .C (CLK), .D (signal_8360), .Q (signal_8361) ) ;
    buf_clk cell_6233 ( .C (CLK), .D (signal_8376), .Q (signal_8377) ) ;
    buf_clk cell_6249 ( .C (CLK), .D (signal_8392), .Q (signal_8393) ) ;
    buf_clk cell_6265 ( .C (CLK), .D (signal_8408), .Q (signal_8409) ) ;
    buf_clk cell_6281 ( .C (CLK), .D (signal_8424), .Q (signal_8425) ) ;
    buf_clk cell_6297 ( .C (CLK), .D (signal_8440), .Q (signal_8441) ) ;
    buf_clk cell_6313 ( .C (CLK), .D (signal_8456), .Q (signal_8457) ) ;
    buf_clk cell_6329 ( .C (CLK), .D (signal_8472), .Q (signal_8473) ) ;
    buf_clk cell_6345 ( .C (CLK), .D (signal_8488), .Q (signal_8489) ) ;
    buf_clk cell_6361 ( .C (CLK), .D (signal_8504), .Q (signal_8505) ) ;
    buf_clk cell_6377 ( .C (CLK), .D (signal_8520), .Q (signal_8521) ) ;
    buf_clk cell_6393 ( .C (CLK), .D (signal_8536), .Q (signal_8537) ) ;
    buf_clk cell_7593 ( .C (CLK), .D (signal_9736), .Q (signal_9737) ) ;
    buf_clk cell_7609 ( .C (CLK), .D (signal_9752), .Q (signal_9753) ) ;
    buf_clk cell_7625 ( .C (CLK), .D (signal_9768), .Q (signal_9769) ) ;
    buf_clk cell_7641 ( .C (CLK), .D (signal_9784), .Q (signal_9785) ) ;
    buf_clk cell_7657 ( .C (CLK), .D (signal_9800), .Q (signal_9801) ) ;
    buf_clk cell_7673 ( .C (CLK), .D (signal_9816), .Q (signal_9817) ) ;
    buf_clk cell_7689 ( .C (CLK), .D (signal_9832), .Q (signal_9833) ) ;
    buf_clk cell_7705 ( .C (CLK), .D (signal_9848), .Q (signal_9849) ) ;
    buf_clk cell_7721 ( .C (CLK), .D (signal_9864), .Q (signal_9865) ) ;
    buf_clk cell_7737 ( .C (CLK), .D (signal_9880), .Q (signal_9881) ) ;
    buf_clk cell_7945 ( .C (CLK), .D (signal_10088), .Q (signal_10089) ) ;

    /* cells in depth 5 */
    buf_clk cell_2194 ( .C (CLK), .D (signal_4337), .Q (signal_4338) ) ;
    buf_clk cell_2202 ( .C (CLK), .D (signal_4345), .Q (signal_4346) ) ;
    buf_clk cell_2210 ( .C (CLK), .D (signal_4353), .Q (signal_4354) ) ;
    buf_clk cell_2218 ( .C (CLK), .D (signal_4361), .Q (signal_4362) ) ;
    buf_clk cell_2226 ( .C (CLK), .D (signal_4369), .Q (signal_4370) ) ;
    buf_clk cell_2234 ( .C (CLK), .D (signal_4377), .Q (signal_4378) ) ;
    buf_clk cell_2242 ( .C (CLK), .D (signal_4385), .Q (signal_4386) ) ;
    buf_clk cell_2250 ( .C (CLK), .D (signal_4393), .Q (signal_4394) ) ;
    buf_clk cell_2258 ( .C (CLK), .D (signal_4401), .Q (signal_4402) ) ;
    buf_clk cell_2266 ( .C (CLK), .D (signal_4409), .Q (signal_4410) ) ;
    buf_clk cell_2270 ( .C (CLK), .D (signal_3957), .Q (signal_4414) ) ;
    buf_clk cell_2274 ( .C (CLK), .D (signal_3961), .Q (signal_4418) ) ;
    buf_clk cell_2282 ( .C (CLK), .D (signal_4425), .Q (signal_4426) ) ;
    buf_clk cell_2290 ( .C (CLK), .D (signal_4433), .Q (signal_4434) ) ;
    buf_clk cell_2294 ( .C (CLK), .D (signal_3969), .Q (signal_4438) ) ;
    buf_clk cell_2298 ( .C (CLK), .D (signal_3973), .Q (signal_4442) ) ;
    buf_clk cell_2302 ( .C (CLK), .D (signal_4321), .Q (signal_4446) ) ;
    buf_clk cell_2306 ( .C (CLK), .D (signal_4325), .Q (signal_4450) ) ;
    buf_clk cell_2314 ( .C (CLK), .D (signal_4457), .Q (signal_4458) ) ;
    buf_clk cell_2322 ( .C (CLK), .D (signal_4465), .Q (signal_4466) ) ;
    buf_clk cell_2330 ( .C (CLK), .D (signal_4473), .Q (signal_4474) ) ;
    buf_clk cell_2338 ( .C (CLK), .D (signal_4481), .Q (signal_4482) ) ;
    buf_clk cell_2342 ( .C (CLK), .D (signal_3981), .Q (signal_4486) ) ;
    buf_clk cell_2346 ( .C (CLK), .D (signal_3985), .Q (signal_4490) ) ;
    buf_clk cell_2354 ( .C (CLK), .D (signal_4497), .Q (signal_4498) ) ;
    buf_clk cell_2360 ( .C (CLK), .D (signal_4503), .Q (signal_4504) ) ;
    buf_clk cell_2366 ( .C (CLK), .D (signal_4509), .Q (signal_4510) ) ;
    buf_clk cell_2374 ( .C (CLK), .D (signal_4517), .Q (signal_4518) ) ;
    buf_clk cell_2382 ( .C (CLK), .D (signal_4525), .Q (signal_4526) ) ;
    buf_clk cell_2390 ( .C (CLK), .D (signal_4533), .Q (signal_4534) ) ;
    buf_clk cell_2398 ( .C (CLK), .D (signal_4541), .Q (signal_4542) ) ;
    buf_clk cell_2406 ( .C (CLK), .D (signal_4549), .Q (signal_4550) ) ;
    buf_clk cell_2414 ( .C (CLK), .D (signal_4557), .Q (signal_4558) ) ;
    buf_clk cell_2422 ( .C (CLK), .D (signal_4565), .Q (signal_4566) ) ;
    buf_clk cell_2430 ( .C (CLK), .D (signal_4573), .Q (signal_4574) ) ;
    buf_clk cell_2438 ( .C (CLK), .D (signal_4581), .Q (signal_4582) ) ;
    buf_clk cell_2446 ( .C (CLK), .D (signal_4589), .Q (signal_4590) ) ;
    buf_clk cell_2454 ( .C (CLK), .D (signal_4597), .Q (signal_4598) ) ;
    buf_clk cell_2462 ( .C (CLK), .D (signal_4605), .Q (signal_4606) ) ;
    buf_clk cell_2470 ( .C (CLK), .D (signal_4613), .Q (signal_4614) ) ;
    buf_clk cell_2478 ( .C (CLK), .D (signal_4621), .Q (signal_4622) ) ;
    buf_clk cell_2486 ( .C (CLK), .D (signal_4629), .Q (signal_4630) ) ;
    buf_clk cell_2494 ( .C (CLK), .D (signal_4637), .Q (signal_4638) ) ;
    buf_clk cell_2502 ( .C (CLK), .D (signal_4645), .Q (signal_4646) ) ;
    buf_clk cell_2510 ( .C (CLK), .D (signal_4653), .Q (signal_4654) ) ;
    buf_clk cell_2518 ( .C (CLK), .D (signal_4661), .Q (signal_4662) ) ;
    buf_clk cell_2526 ( .C (CLK), .D (signal_4669), .Q (signal_4670) ) ;
    buf_clk cell_2534 ( .C (CLK), .D (signal_4677), .Q (signal_4678) ) ;
    buf_clk cell_2542 ( .C (CLK), .D (signal_4685), .Q (signal_4686) ) ;
    buf_clk cell_2550 ( .C (CLK), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_2558 ( .C (CLK), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_2566 ( .C (CLK), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_2570 ( .C (CLK), .D (signal_4053), .Q (signal_4714) ) ;
    buf_clk cell_2574 ( .C (CLK), .D (signal_4057), .Q (signal_4718) ) ;
    buf_clk cell_2578 ( .C (CLK), .D (signal_4315), .Q (signal_4722) ) ;
    buf_clk cell_2582 ( .C (CLK), .D (signal_4317), .Q (signal_4726) ) ;
    buf_clk cell_2590 ( .C (CLK), .D (signal_4733), .Q (signal_4734) ) ;
    buf_clk cell_2598 ( .C (CLK), .D (signal_4741), .Q (signal_4742) ) ;
    buf_clk cell_2606 ( .C (CLK), .D (signal_4749), .Q (signal_4750) ) ;
    buf_clk cell_2614 ( .C (CLK), .D (signal_4757), .Q (signal_4758) ) ;
    buf_clk cell_2618 ( .C (CLK), .D (signal_4085), .Q (signal_4762) ) ;
    buf_clk cell_2622 ( .C (CLK), .D (signal_4089), .Q (signal_4766) ) ;
    buf_clk cell_2628 ( .C (CLK), .D (signal_4771), .Q (signal_4772) ) ;
    buf_clk cell_2634 ( .C (CLK), .D (signal_4777), .Q (signal_4778) ) ;
    buf_clk cell_2642 ( .C (CLK), .D (signal_4785), .Q (signal_4786) ) ;
    buf_clk cell_2650 ( .C (CLK), .D (signal_4793), .Q (signal_4794) ) ;
    buf_clk cell_2658 ( .C (CLK), .D (signal_4801), .Q (signal_4802) ) ;
    buf_clk cell_2666 ( .C (CLK), .D (signal_4809), .Q (signal_4810) ) ;
    buf_clk cell_2672 ( .C (CLK), .D (signal_4815), .Q (signal_4816) ) ;
    buf_clk cell_2678 ( .C (CLK), .D (signal_4821), .Q (signal_4822) ) ;
    buf_clk cell_2682 ( .C (CLK), .D (signal_4129), .Q (signal_4826) ) ;
    buf_clk cell_2686 ( .C (CLK), .D (signal_4133), .Q (signal_4830) ) ;
    buf_clk cell_2694 ( .C (CLK), .D (signal_4837), .Q (signal_4838) ) ;
    buf_clk cell_2702 ( .C (CLK), .D (signal_4845), .Q (signal_4846) ) ;
    buf_clk cell_2710 ( .C (CLK), .D (signal_4853), .Q (signal_4854) ) ;
    buf_clk cell_2718 ( .C (CLK), .D (signal_4861), .Q (signal_4862) ) ;
    buf_clk cell_2726 ( .C (CLK), .D (signal_4869), .Q (signal_4870) ) ;
    buf_clk cell_2734 ( .C (CLK), .D (signal_4877), .Q (signal_4878) ) ;
    buf_clk cell_2742 ( .C (CLK), .D (signal_4885), .Q (signal_4886) ) ;
    buf_clk cell_2750 ( .C (CLK), .D (signal_4893), .Q (signal_4894) ) ;
    buf_clk cell_2758 ( .C (CLK), .D (signal_4901), .Q (signal_4902) ) ;
    buf_clk cell_2766 ( .C (CLK), .D (signal_4909), .Q (signal_4910) ) ;
    buf_clk cell_2774 ( .C (CLK), .D (signal_4917), .Q (signal_4918) ) ;
    buf_clk cell_2782 ( .C (CLK), .D (signal_4925), .Q (signal_4926) ) ;
    buf_clk cell_2790 ( .C (CLK), .D (signal_4933), .Q (signal_4934) ) ;
    buf_clk cell_2796 ( .C (CLK), .D (signal_4939), .Q (signal_4940) ) ;
    buf_clk cell_2802 ( .C (CLK), .D (signal_4945), .Q (signal_4946) ) ;
    buf_clk cell_2808 ( .C (CLK), .D (signal_4951), .Q (signal_4952) ) ;
    buf_clk cell_2814 ( .C (CLK), .D (signal_4957), .Q (signal_4958) ) ;
    buf_clk cell_2820 ( .C (CLK), .D (signal_4963), .Q (signal_4964) ) ;
    buf_clk cell_2826 ( .C (CLK), .D (signal_4969), .Q (signal_4970) ) ;
    buf_clk cell_2832 ( .C (CLK), .D (signal_4975), .Q (signal_4976) ) ;
    buf_clk cell_2838 ( .C (CLK), .D (signal_4981), .Q (signal_4982) ) ;
    buf_clk cell_2844 ( .C (CLK), .D (signal_4987), .Q (signal_4988) ) ;
    buf_clk cell_2850 ( .C (CLK), .D (signal_4993), .Q (signal_4994) ) ;
    buf_clk cell_2856 ( .C (CLK), .D (signal_4999), .Q (signal_5000) ) ;
    buf_clk cell_2862 ( .C (CLK), .D (signal_5005), .Q (signal_5006) ) ;
    buf_clk cell_2868 ( .C (CLK), .D (signal_5011), .Q (signal_5012) ) ;
    buf_clk cell_2870 ( .C (CLK), .D (signal_4005), .Q (signal_5014) ) ;
    buf_clk cell_2872 ( .C (CLK), .D (signal_4009), .Q (signal_5016) ) ;
    buf_clk cell_2874 ( .C (CLK), .D (signal_1443), .Q (signal_5018) ) ;
    buf_clk cell_2876 ( .C (CLK), .D (signal_2400), .Q (signal_5020) ) ;
    buf_clk cell_2878 ( .C (CLK), .D (signal_4227), .Q (signal_5022) ) ;
    buf_clk cell_2880 ( .C (CLK), .D (signal_4229), .Q (signal_5024) ) ;
    buf_clk cell_2882 ( .C (CLK), .D (signal_1412), .Q (signal_5026) ) ;
    buf_clk cell_2884 ( .C (CLK), .D (signal_2386), .Q (signal_5028) ) ;
    buf_clk cell_2886 ( .C (CLK), .D (signal_1445), .Q (signal_5030) ) ;
    buf_clk cell_2888 ( .C (CLK), .D (signal_2402), .Q (signal_5032) ) ;
    buf_clk cell_2890 ( .C (CLK), .D (signal_1446), .Q (signal_5034) ) ;
    buf_clk cell_2892 ( .C (CLK), .D (signal_2403), .Q (signal_5036) ) ;
    buf_clk cell_2894 ( .C (CLK), .D (signal_1447), .Q (signal_5038) ) ;
    buf_clk cell_2896 ( .C (CLK), .D (signal_2404), .Q (signal_5040) ) ;
    buf_clk cell_2898 ( .C (CLK), .D (signal_4099), .Q (signal_5042) ) ;
    buf_clk cell_2900 ( .C (CLK), .D (signal_4101), .Q (signal_5044) ) ;
    buf_clk cell_2902 ( .C (CLK), .D (signal_4239), .Q (signal_5046) ) ;
    buf_clk cell_2904 ( .C (CLK), .D (signal_4241), .Q (signal_5048) ) ;
    buf_clk cell_2906 ( .C (CLK), .D (signal_1476), .Q (signal_5050) ) ;
    buf_clk cell_2908 ( .C (CLK), .D (signal_2420), .Q (signal_5052) ) ;
    buf_clk cell_2910 ( .C (CLK), .D (signal_4291), .Q (signal_5054) ) ;
    buf_clk cell_2912 ( .C (CLK), .D (signal_4293), .Q (signal_5056) ) ;
    buf_clk cell_2914 ( .C (CLK), .D (signal_1477), .Q (signal_5058) ) ;
    buf_clk cell_2916 ( .C (CLK), .D (signal_2421), .Q (signal_5060) ) ;
    buf_clk cell_2918 ( .C (CLK), .D (signal_1478), .Q (signal_5062) ) ;
    buf_clk cell_2920 ( .C (CLK), .D (signal_2422), .Q (signal_5064) ) ;
    buf_clk cell_2922 ( .C (CLK), .D (signal_1480), .Q (signal_5066) ) ;
    buf_clk cell_2924 ( .C (CLK), .D (signal_2424), .Q (signal_5068) ) ;
    buf_clk cell_2926 ( .C (CLK), .D (signal_1481), .Q (signal_5070) ) ;
    buf_clk cell_2928 ( .C (CLK), .D (signal_2425), .Q (signal_5072) ) ;
    buf_clk cell_2930 ( .C (CLK), .D (signal_1482), .Q (signal_5074) ) ;
    buf_clk cell_2932 ( .C (CLK), .D (signal_2426), .Q (signal_5076) ) ;
    buf_clk cell_2936 ( .C (CLK), .D (signal_5079), .Q (signal_5080) ) ;
    buf_clk cell_2940 ( .C (CLK), .D (signal_5083), .Q (signal_5084) ) ;
    buf_clk cell_2942 ( .C (CLK), .D (signal_1487), .Q (signal_5086) ) ;
    buf_clk cell_2944 ( .C (CLK), .D (signal_2429), .Q (signal_5088) ) ;
    buf_clk cell_2946 ( .C (CLK), .D (signal_1488), .Q (signal_5090) ) ;
    buf_clk cell_2948 ( .C (CLK), .D (signal_2430), .Q (signal_5092) ) ;
    buf_clk cell_2950 ( .C (CLK), .D (signal_4145), .Q (signal_5094) ) ;
    buf_clk cell_2952 ( .C (CLK), .D (signal_4149), .Q (signal_5096) ) ;
    buf_clk cell_2954 ( .C (CLK), .D (signal_1491), .Q (signal_5098) ) ;
    buf_clk cell_2956 ( .C (CLK), .D (signal_2433), .Q (signal_5100) ) ;
    buf_clk cell_2958 ( .C (CLK), .D (signal_1493), .Q (signal_5102) ) ;
    buf_clk cell_2960 ( .C (CLK), .D (signal_2435), .Q (signal_5104) ) ;
    buf_clk cell_2962 ( .C (CLK), .D (signal_1494), .Q (signal_5106) ) ;
    buf_clk cell_2964 ( .C (CLK), .D (signal_2436), .Q (signal_5108) ) ;
    buf_clk cell_2966 ( .C (CLK), .D (signal_1495), .Q (signal_5110) ) ;
    buf_clk cell_2968 ( .C (CLK), .D (signal_2437), .Q (signal_5112) ) ;
    buf_clk cell_2974 ( .C (CLK), .D (signal_5117), .Q (signal_5118) ) ;
    buf_clk cell_2980 ( .C (CLK), .D (signal_5123), .Q (signal_5124) ) ;
    buf_clk cell_2984 ( .C (CLK), .D (signal_5127), .Q (signal_5128) ) ;
    buf_clk cell_2988 ( .C (CLK), .D (signal_5131), .Q (signal_5132) ) ;
    buf_clk cell_2990 ( .C (CLK), .D (signal_4327), .Q (signal_5134) ) ;
    buf_clk cell_2992 ( .C (CLK), .D (signal_4329), .Q (signal_5136) ) ;
    buf_clk cell_2994 ( .C (CLK), .D (signal_1500), .Q (signal_5138) ) ;
    buf_clk cell_2996 ( .C (CLK), .D (signal_2440), .Q (signal_5140) ) ;
    buf_clk cell_2998 ( .C (CLK), .D (signal_1501), .Q (signal_5142) ) ;
    buf_clk cell_3000 ( .C (CLK), .D (signal_2441), .Q (signal_5144) ) ;
    buf_clk cell_3002 ( .C (CLK), .D (signal_1504), .Q (signal_5146) ) ;
    buf_clk cell_3004 ( .C (CLK), .D (signal_2442), .Q (signal_5148) ) ;
    buf_clk cell_3006 ( .C (CLK), .D (signal_1444), .Q (signal_5150) ) ;
    buf_clk cell_3008 ( .C (CLK), .D (signal_2401), .Q (signal_5152) ) ;
    buf_clk cell_3016 ( .C (CLK), .D (signal_5159), .Q (signal_5160) ) ;
    buf_clk cell_3022 ( .C (CLK), .D (signal_5165), .Q (signal_5166) ) ;
    buf_clk cell_3058 ( .C (CLK), .D (signal_5201), .Q (signal_5202) ) ;
    buf_clk cell_3066 ( .C (CLK), .D (signal_5209), .Q (signal_5210) ) ;
    buf_clk cell_3086 ( .C (CLK), .D (signal_4041), .Q (signal_5230) ) ;
    buf_clk cell_3090 ( .C (CLK), .D (signal_4045), .Q (signal_5234) ) ;
    buf_clk cell_3196 ( .C (CLK), .D (signal_5339), .Q (signal_5340) ) ;
    buf_clk cell_3204 ( .C (CLK), .D (signal_5347), .Q (signal_5348) ) ;
    buf_clk cell_3318 ( .C (CLK), .D (signal_3993), .Q (signal_5462) ) ;
    buf_clk cell_3326 ( .C (CLK), .D (signal_3997), .Q (signal_5470) ) ;
    buf_clk cell_3354 ( .C (CLK), .D (signal_4069), .Q (signal_5498) ) ;
    buf_clk cell_3362 ( .C (CLK), .D (signal_4073), .Q (signal_5506) ) ;
    buf_clk cell_3450 ( .C (CLK), .D (signal_5593), .Q (signal_5594) ) ;
    buf_clk cell_3466 ( .C (CLK), .D (signal_5609), .Q (signal_5610) ) ;
    buf_clk cell_3490 ( .C (CLK), .D (signal_5633), .Q (signal_5634) ) ;
    buf_clk cell_3506 ( .C (CLK), .D (signal_5649), .Q (signal_5650) ) ;
    buf_clk cell_3530 ( .C (CLK), .D (signal_5673), .Q (signal_5674) ) ;
    buf_clk cell_3546 ( .C (CLK), .D (signal_5689), .Q (signal_5690) ) ;
    buf_clk cell_3562 ( .C (CLK), .D (signal_5705), .Q (signal_5706) ) ;
    buf_clk cell_3578 ( .C (CLK), .D (signal_5721), .Q (signal_5722) ) ;
    buf_clk cell_3638 ( .C (CLK), .D (signal_5781), .Q (signal_5782) ) ;
    buf_clk cell_3654 ( .C (CLK), .D (signal_5797), .Q (signal_5798) ) ;
    buf_clk cell_3670 ( .C (CLK), .D (signal_5813), .Q (signal_5814) ) ;
    buf_clk cell_3686 ( .C (CLK), .D (signal_5829), .Q (signal_5830) ) ;
    buf_clk cell_3702 ( .C (CLK), .D (signal_5845), .Q (signal_5846) ) ;
    buf_clk cell_3718 ( .C (CLK), .D (signal_5861), .Q (signal_5862) ) ;
    buf_clk cell_3734 ( .C (CLK), .D (signal_5877), .Q (signal_5878) ) ;
    buf_clk cell_3750 ( .C (CLK), .D (signal_5893), .Q (signal_5894) ) ;
    buf_clk cell_3766 ( .C (CLK), .D (signal_5909), .Q (signal_5910) ) ;
    buf_clk cell_3782 ( .C (CLK), .D (signal_5925), .Q (signal_5926) ) ;
    buf_clk cell_3890 ( .C (CLK), .D (signal_6033), .Q (signal_6034) ) ;
    buf_clk cell_3906 ( .C (CLK), .D (signal_6049), .Q (signal_6050) ) ;
    buf_clk cell_3922 ( .C (CLK), .D (signal_6065), .Q (signal_6066) ) ;
    buf_clk cell_3938 ( .C (CLK), .D (signal_6081), .Q (signal_6082) ) ;
    buf_clk cell_3954 ( .C (CLK), .D (signal_6097), .Q (signal_6098) ) ;
    buf_clk cell_3970 ( .C (CLK), .D (signal_6113), .Q (signal_6114) ) ;
    buf_clk cell_3986 ( .C (CLK), .D (signal_6129), .Q (signal_6130) ) ;
    buf_clk cell_4002 ( .C (CLK), .D (signal_6145), .Q (signal_6146) ) ;
    buf_clk cell_4018 ( .C (CLK), .D (signal_6161), .Q (signal_6162) ) ;
    buf_clk cell_4034 ( .C (CLK), .D (signal_6177), .Q (signal_6178) ) ;
    buf_clk cell_4050 ( .C (CLK), .D (signal_6193), .Q (signal_6194) ) ;
    buf_clk cell_4066 ( .C (CLK), .D (signal_6209), .Q (signal_6210) ) ;
    buf_clk cell_4082 ( .C (CLK), .D (signal_6225), .Q (signal_6226) ) ;
    buf_clk cell_4098 ( .C (CLK), .D (signal_6241), .Q (signal_6242) ) ;
    buf_clk cell_4182 ( .C (CLK), .D (signal_6325), .Q (signal_6326) ) ;
    buf_clk cell_4194 ( .C (CLK), .D (signal_4231), .Q (signal_6338) ) ;
    buf_clk cell_4206 ( .C (CLK), .D (signal_4233), .Q (signal_6350) ) ;
    buf_clk cell_4234 ( .C (CLK), .D (signal_4017), .Q (signal_6378) ) ;
    buf_clk cell_4246 ( .C (CLK), .D (signal_4021), .Q (signal_6390) ) ;
    buf_clk cell_4260 ( .C (CLK), .D (signal_6403), .Q (signal_6404) ) ;
    buf_clk cell_4274 ( .C (CLK), .D (signal_6417), .Q (signal_6418) ) ;
    buf_clk cell_4290 ( .C (CLK), .D (signal_6433), .Q (signal_6434) ) ;
    buf_clk cell_4306 ( .C (CLK), .D (signal_6449), .Q (signal_6450) ) ;
    buf_clk cell_4322 ( .C (CLK), .D (signal_6465), .Q (signal_6466) ) ;
    buf_clk cell_4338 ( .C (CLK), .D (signal_6481), .Q (signal_6482) ) ;
    buf_clk cell_4354 ( .C (CLK), .D (signal_6497), .Q (signal_6498) ) ;
    buf_clk cell_4370 ( .C (CLK), .D (signal_6513), .Q (signal_6514) ) ;
    buf_clk cell_4386 ( .C (CLK), .D (signal_6529), .Q (signal_6530) ) ;
    buf_clk cell_4402 ( .C (CLK), .D (signal_6545), .Q (signal_6546) ) ;
    buf_clk cell_4418 ( .C (CLK), .D (signal_6561), .Q (signal_6562) ) ;
    buf_clk cell_4434 ( .C (CLK), .D (signal_6577), .Q (signal_6578) ) ;
    buf_clk cell_4450 ( .C (CLK), .D (signal_6593), .Q (signal_6594) ) ;
    buf_clk cell_4466 ( .C (CLK), .D (signal_6609), .Q (signal_6610) ) ;
    buf_clk cell_4482 ( .C (CLK), .D (signal_6625), .Q (signal_6626) ) ;
    buf_clk cell_4498 ( .C (CLK), .D (signal_6641), .Q (signal_6642) ) ;
    buf_clk cell_4514 ( .C (CLK), .D (signal_6657), .Q (signal_6658) ) ;
    buf_clk cell_4530 ( .C (CLK), .D (signal_6673), .Q (signal_6674) ) ;
    buf_clk cell_4578 ( .C (CLK), .D (signal_4029), .Q (signal_6722) ) ;
    buf_clk cell_4590 ( .C (CLK), .D (signal_4033), .Q (signal_6734) ) ;
    buf_clk cell_4604 ( .C (CLK), .D (signal_6747), .Q (signal_6748) ) ;
    buf_clk cell_4618 ( .C (CLK), .D (signal_6761), .Q (signal_6762) ) ;
    buf_clk cell_4634 ( .C (CLK), .D (signal_6777), .Q (signal_6778) ) ;
    buf_clk cell_4650 ( .C (CLK), .D (signal_6793), .Q (signal_6794) ) ;
    buf_clk cell_4710 ( .C (CLK), .D (signal_4305), .Q (signal_6854) ) ;
    buf_clk cell_4722 ( .C (CLK), .D (signal_4309), .Q (signal_6866) ) ;
    buf_clk cell_4746 ( .C (CLK), .D (signal_6889), .Q (signal_6890) ) ;
    buf_clk cell_4762 ( .C (CLK), .D (signal_6905), .Q (signal_6906) ) ;
    buf_clk cell_4778 ( .C (CLK), .D (signal_6921), .Q (signal_6922) ) ;
    buf_clk cell_4794 ( .C (CLK), .D (signal_6937), .Q (signal_6938) ) ;
    buf_clk cell_4810 ( .C (CLK), .D (signal_6953), .Q (signal_6954) ) ;
    buf_clk cell_4826 ( .C (CLK), .D (signal_6969), .Q (signal_6970) ) ;
    buf_clk cell_4842 ( .C (CLK), .D (signal_6985), .Q (signal_6986) ) ;
    buf_clk cell_4858 ( .C (CLK), .D (signal_7001), .Q (signal_7002) ) ;
    buf_clk cell_4874 ( .C (CLK), .D (signal_7017), .Q (signal_7018) ) ;
    buf_clk cell_4890 ( .C (CLK), .D (signal_7033), .Q (signal_7034) ) ;
    buf_clk cell_4906 ( .C (CLK), .D (signal_7049), .Q (signal_7050) ) ;
    buf_clk cell_4922 ( .C (CLK), .D (signal_7065), .Q (signal_7066) ) ;
    buf_clk cell_4938 ( .C (CLK), .D (signal_7081), .Q (signal_7082) ) ;
    buf_clk cell_4954 ( .C (CLK), .D (signal_7097), .Q (signal_7098) ) ;
    buf_clk cell_4970 ( .C (CLK), .D (signal_7113), .Q (signal_7114) ) ;
    buf_clk cell_4986 ( .C (CLK), .D (signal_7129), .Q (signal_7130) ) ;
    buf_clk cell_5002 ( .C (CLK), .D (signal_7145), .Q (signal_7146) ) ;
    buf_clk cell_5018 ( .C (CLK), .D (signal_7161), .Q (signal_7162) ) ;
    buf_clk cell_5034 ( .C (CLK), .D (signal_7177), .Q (signal_7178) ) ;
    buf_clk cell_5050 ( .C (CLK), .D (signal_7193), .Q (signal_7194) ) ;
    buf_clk cell_5066 ( .C (CLK), .D (signal_7209), .Q (signal_7210) ) ;
    buf_clk cell_5082 ( .C (CLK), .D (signal_7225), .Q (signal_7226) ) ;
    buf_clk cell_5098 ( .C (CLK), .D (signal_7241), .Q (signal_7242) ) ;
    buf_clk cell_5114 ( .C (CLK), .D (signal_7257), .Q (signal_7258) ) ;
    buf_clk cell_5130 ( .C (CLK), .D (signal_7273), .Q (signal_7274) ) ;
    buf_clk cell_5146 ( .C (CLK), .D (signal_7289), .Q (signal_7290) ) ;
    buf_clk cell_5162 ( .C (CLK), .D (signal_7305), .Q (signal_7306) ) ;
    buf_clk cell_5178 ( .C (CLK), .D (signal_7321), .Q (signal_7322) ) ;
    buf_clk cell_5194 ( .C (CLK), .D (signal_7337), .Q (signal_7338) ) ;
    buf_clk cell_5210 ( .C (CLK), .D (signal_7353), .Q (signal_7354) ) ;
    buf_clk cell_5226 ( .C (CLK), .D (signal_7369), .Q (signal_7370) ) ;
    buf_clk cell_5242 ( .C (CLK), .D (signal_7385), .Q (signal_7386) ) ;
    buf_clk cell_5258 ( .C (CLK), .D (signal_7401), .Q (signal_7402) ) ;
    buf_clk cell_5274 ( .C (CLK), .D (signal_7417), .Q (signal_7418) ) ;
    buf_clk cell_5290 ( .C (CLK), .D (signal_7433), .Q (signal_7434) ) ;
    buf_clk cell_5306 ( .C (CLK), .D (signal_7449), .Q (signal_7450) ) ;
    buf_clk cell_5322 ( .C (CLK), .D (signal_7465), .Q (signal_7466) ) ;
    buf_clk cell_5338 ( .C (CLK), .D (signal_7481), .Q (signal_7482) ) ;
    buf_clk cell_5354 ( .C (CLK), .D (signal_7497), .Q (signal_7498) ) ;
    buf_clk cell_5370 ( .C (CLK), .D (signal_7513), .Q (signal_7514) ) ;
    buf_clk cell_5386 ( .C (CLK), .D (signal_7529), .Q (signal_7530) ) ;
    buf_clk cell_5402 ( .C (CLK), .D (signal_7545), .Q (signal_7546) ) ;
    buf_clk cell_5418 ( .C (CLK), .D (signal_7561), .Q (signal_7562) ) ;
    buf_clk cell_5434 ( .C (CLK), .D (signal_7577), .Q (signal_7578) ) ;
    buf_clk cell_5450 ( .C (CLK), .D (signal_7593), .Q (signal_7594) ) ;
    buf_clk cell_5466 ( .C (CLK), .D (signal_7609), .Q (signal_7610) ) ;
    buf_clk cell_5482 ( .C (CLK), .D (signal_7625), .Q (signal_7626) ) ;
    buf_clk cell_5498 ( .C (CLK), .D (signal_7641), .Q (signal_7642) ) ;
    buf_clk cell_5514 ( .C (CLK), .D (signal_7657), .Q (signal_7658) ) ;
    buf_clk cell_5530 ( .C (CLK), .D (signal_7673), .Q (signal_7674) ) ;
    buf_clk cell_5546 ( .C (CLK), .D (signal_7689), .Q (signal_7690) ) ;
    buf_clk cell_5562 ( .C (CLK), .D (signal_7705), .Q (signal_7706) ) ;
    buf_clk cell_5578 ( .C (CLK), .D (signal_7721), .Q (signal_7722) ) ;
    buf_clk cell_5594 ( .C (CLK), .D (signal_7737), .Q (signal_7738) ) ;
    buf_clk cell_5610 ( .C (CLK), .D (signal_7753), .Q (signal_7754) ) ;
    buf_clk cell_5626 ( .C (CLK), .D (signal_7769), .Q (signal_7770) ) ;
    buf_clk cell_5642 ( .C (CLK), .D (signal_7785), .Q (signal_7786) ) ;
    buf_clk cell_5658 ( .C (CLK), .D (signal_7801), .Q (signal_7802) ) ;
    buf_clk cell_5674 ( .C (CLK), .D (signal_7817), .Q (signal_7818) ) ;
    buf_clk cell_5690 ( .C (CLK), .D (signal_7833), .Q (signal_7834) ) ;
    buf_clk cell_5706 ( .C (CLK), .D (signal_7849), .Q (signal_7850) ) ;
    buf_clk cell_5722 ( .C (CLK), .D (signal_7865), .Q (signal_7866) ) ;
    buf_clk cell_5738 ( .C (CLK), .D (signal_7881), .Q (signal_7882) ) ;
    buf_clk cell_5754 ( .C (CLK), .D (signal_7897), .Q (signal_7898) ) ;
    buf_clk cell_5770 ( .C (CLK), .D (signal_7913), .Q (signal_7914) ) ;
    buf_clk cell_5786 ( .C (CLK), .D (signal_7929), .Q (signal_7930) ) ;
    buf_clk cell_5802 ( .C (CLK), .D (signal_7945), .Q (signal_7946) ) ;
    buf_clk cell_5818 ( .C (CLK), .D (signal_7961), .Q (signal_7962) ) ;
    buf_clk cell_5834 ( .C (CLK), .D (signal_7977), .Q (signal_7978) ) ;
    buf_clk cell_5850 ( .C (CLK), .D (signal_7993), .Q (signal_7994) ) ;
    buf_clk cell_5866 ( .C (CLK), .D (signal_8009), .Q (signal_8010) ) ;
    buf_clk cell_5882 ( .C (CLK), .D (signal_8025), .Q (signal_8026) ) ;
    buf_clk cell_5898 ( .C (CLK), .D (signal_8041), .Q (signal_8042) ) ;
    buf_clk cell_5914 ( .C (CLK), .D (signal_8057), .Q (signal_8058) ) ;
    buf_clk cell_5930 ( .C (CLK), .D (signal_8073), .Q (signal_8074) ) ;
    buf_clk cell_5946 ( .C (CLK), .D (signal_8089), .Q (signal_8090) ) ;
    buf_clk cell_5962 ( .C (CLK), .D (signal_8105), .Q (signal_8106) ) ;
    buf_clk cell_5978 ( .C (CLK), .D (signal_8121), .Q (signal_8122) ) ;
    buf_clk cell_5994 ( .C (CLK), .D (signal_8137), .Q (signal_8138) ) ;
    buf_clk cell_6010 ( .C (CLK), .D (signal_8153), .Q (signal_8154) ) ;
    buf_clk cell_6026 ( .C (CLK), .D (signal_8169), .Q (signal_8170) ) ;
    buf_clk cell_6042 ( .C (CLK), .D (signal_8185), .Q (signal_8186) ) ;
    buf_clk cell_6058 ( .C (CLK), .D (signal_8201), .Q (signal_8202) ) ;
    buf_clk cell_6074 ( .C (CLK), .D (signal_8217), .Q (signal_8218) ) ;
    buf_clk cell_6090 ( .C (CLK), .D (signal_8233), .Q (signal_8234) ) ;
    buf_clk cell_6106 ( .C (CLK), .D (signal_8249), .Q (signal_8250) ) ;
    buf_clk cell_6122 ( .C (CLK), .D (signal_8265), .Q (signal_8266) ) ;
    buf_clk cell_6138 ( .C (CLK), .D (signal_8281), .Q (signal_8282) ) ;
    buf_clk cell_6154 ( .C (CLK), .D (signal_8297), .Q (signal_8298) ) ;
    buf_clk cell_6170 ( .C (CLK), .D (signal_8313), .Q (signal_8314) ) ;
    buf_clk cell_6186 ( .C (CLK), .D (signal_8329), .Q (signal_8330) ) ;
    buf_clk cell_6202 ( .C (CLK), .D (signal_8345), .Q (signal_8346) ) ;
    buf_clk cell_6218 ( .C (CLK), .D (signal_8361), .Q (signal_8362) ) ;
    buf_clk cell_6234 ( .C (CLK), .D (signal_8377), .Q (signal_8378) ) ;
    buf_clk cell_6250 ( .C (CLK), .D (signal_8393), .Q (signal_8394) ) ;
    buf_clk cell_6266 ( .C (CLK), .D (signal_8409), .Q (signal_8410) ) ;
    buf_clk cell_6282 ( .C (CLK), .D (signal_8425), .Q (signal_8426) ) ;
    buf_clk cell_6298 ( .C (CLK), .D (signal_8441), .Q (signal_8442) ) ;
    buf_clk cell_6314 ( .C (CLK), .D (signal_8457), .Q (signal_8458) ) ;
    buf_clk cell_6330 ( .C (CLK), .D (signal_8473), .Q (signal_8474) ) ;
    buf_clk cell_6346 ( .C (CLK), .D (signal_8489), .Q (signal_8490) ) ;
    buf_clk cell_6362 ( .C (CLK), .D (signal_8505), .Q (signal_8506) ) ;
    buf_clk cell_6378 ( .C (CLK), .D (signal_8521), .Q (signal_8522) ) ;
    buf_clk cell_6394 ( .C (CLK), .D (signal_8537), .Q (signal_8538) ) ;
    buf_clk cell_7594 ( .C (CLK), .D (signal_9737), .Q (signal_9738) ) ;
    buf_clk cell_7610 ( .C (CLK), .D (signal_9753), .Q (signal_9754) ) ;
    buf_clk cell_7626 ( .C (CLK), .D (signal_9769), .Q (signal_9770) ) ;
    buf_clk cell_7642 ( .C (CLK), .D (signal_9785), .Q (signal_9786) ) ;
    buf_clk cell_7658 ( .C (CLK), .D (signal_9801), .Q (signal_9802) ) ;
    buf_clk cell_7674 ( .C (CLK), .D (signal_9817), .Q (signal_9818) ) ;
    buf_clk cell_7690 ( .C (CLK), .D (signal_9833), .Q (signal_9834) ) ;
    buf_clk cell_7706 ( .C (CLK), .D (signal_9849), .Q (signal_9850) ) ;
    buf_clk cell_7722 ( .C (CLK), .D (signal_9865), .Q (signal_9866) ) ;
    buf_clk cell_7738 ( .C (CLK), .D (signal_9881), .Q (signal_9882) ) ;
    buf_clk cell_7946 ( .C (CLK), .D (signal_10089), .Q (signal_10090) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1305 ( .s ({signal_3961, signal_3957}), .b ({signal_2321, signal_1383}), .a ({signal_2320, signal_1382}), .clk (CLK), .r (Fresh[177]), .c ({signal_2443, signal_1505}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1306 ( .s ({signal_3961, signal_3957}), .b ({signal_3965, signal_3963}), .a ({signal_2322, signal_1384}), .clk (CLK), .r (Fresh[178]), .c ({signal_2444, signal_1506}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1307 ( .s ({signal_3973, signal_3969}), .b ({signal_2324, signal_1386}), .a ({signal_2323, signal_1385}), .clk (CLK), .r (Fresh[179]), .c ({signal_2445, signal_1507}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1308 ( .s ({signal_3973, signal_3969}), .b ({signal_3977, signal_3975}), .a ({signal_2325, signal_1387}), .clk (CLK), .r (Fresh[180]), .c ({signal_2446, signal_1508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1309 ( .s ({signal_3985, signal_3981}), .b ({signal_2327, signal_1389}), .a ({signal_2326, signal_1388}), .clk (CLK), .r (Fresh[181]), .c ({signal_2447, signal_1509}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1310 ( .s ({signal_3985, signal_3981}), .b ({signal_2328, signal_1390}), .a ({signal_3989, signal_3987}), .clk (CLK), .r (Fresh[182]), .c ({signal_2448, signal_1510}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1311 ( .s ({signal_3997, signal_3993}), .b ({signal_2330, signal_1392}), .a ({signal_2329, signal_1391}), .clk (CLK), .r (Fresh[183]), .c ({signal_2449, signal_1511}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1312 ( .s ({signal_3997, signal_3993}), .b ({signal_4001, signal_3999}), .a ({signal_2331, signal_1393}), .clk (CLK), .r (Fresh[184]), .c ({signal_2450, signal_1512}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1313 ( .s ({signal_4009, signal_4005}), .b ({signal_2333, signal_1395}), .a ({signal_2332, signal_1394}), .clk (CLK), .r (Fresh[185]), .c ({signal_2451, signal_1513}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1314 ( .s ({signal_4009, signal_4005}), .b ({signal_4013, signal_4011}), .a ({signal_2334, signal_1396}), .clk (CLK), .r (Fresh[186]), .c ({signal_2452, signal_1514}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1315 ( .s ({signal_4021, signal_4017}), .b ({signal_2336, signal_1398}), .a ({signal_2335, signal_1397}), .clk (CLK), .r (Fresh[187]), .c ({signal_2453, signal_1515}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1316 ( .s ({signal_4021, signal_4017}), .b ({signal_4025, signal_4023}), .a ({signal_2337, signal_1399}), .clk (CLK), .r (Fresh[188]), .c ({signal_2454, signal_1516}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1317 ( .s ({signal_4033, signal_4029}), .b ({signal_2339, signal_1401}), .a ({signal_2338, signal_1400}), .clk (CLK), .r (Fresh[189]), .c ({signal_2455, signal_1517}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1318 ( .s ({signal_4033, signal_4029}), .b ({signal_4037, signal_4035}), .a ({signal_2340, signal_1402}), .clk (CLK), .r (Fresh[190]), .c ({signal_2456, signal_1518}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1319 ( .s ({signal_4045, signal_4041}), .b ({signal_2342, signal_1404}), .a ({signal_2341, signal_1403}), .clk (CLK), .r (Fresh[191]), .c ({signal_2457, signal_1519}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1320 ( .s ({signal_4045, signal_4041}), .b ({signal_4049, signal_4047}), .a ({signal_2343, signal_1405}), .clk (CLK), .r (Fresh[192]), .c ({signal_2458, signal_1520}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1321 ( .s ({signal_4057, signal_4053}), .b ({signal_2380, signal_1406}), .a ({signal_4061, signal_4059}), .clk (CLK), .r (Fresh[193]), .c ({signal_2499, signal_1521}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1322 ( .s ({signal_4057, signal_4053}), .b ({signal_2381, signal_1407}), .a ({signal_4065, signal_4063}), .clk (CLK), .r (Fresh[194]), .c ({signal_2500, signal_1522}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1323 ( .s ({signal_4073, signal_4069}), .b ({signal_2382, signal_1408}), .a ({signal_4077, signal_4075}), .clk (CLK), .r (Fresh[195]), .c ({signal_2501, signal_1523}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1324 ( .s ({signal_4073, signal_4069}), .b ({signal_4081, signal_4079}), .a ({signal_2383, signal_1409}), .clk (CLK), .r (Fresh[196]), .c ({signal_2502, signal_1524}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1325 ( .s ({signal_4089, signal_4085}), .b ({signal_2384, signal_1410}), .a ({signal_4093, signal_4091}), .clk (CLK), .r (Fresh[197]), .c ({signal_2503, signal_1525}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1326 ( .s ({signal_4089, signal_4085}), .b ({signal_2385, signal_1411}), .a ({signal_4097, signal_4095}), .clk (CLK), .r (Fresh[198]), .c ({signal_2504, signal_1526}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1327 ( .s ({signal_4101, signal_4099}), .b ({signal_2386, signal_1412}), .a ({signal_4105, signal_4103}), .clk (CLK), .r (Fresh[199]), .c ({signal_2505, signal_1527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1328 ( .s ({signal_4101, signal_4099}), .b ({signal_4109, signal_4107}), .a ({signal_2387, signal_1413}), .clk (CLK), .r (Fresh[200]), .c ({signal_2506, signal_1528}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1329 ( .s ({signal_4117, signal_4113}), .b ({signal_2388, signal_1414}), .a ({signal_4121, signal_4119}), .clk (CLK), .r (Fresh[201]), .c ({signal_2507, signal_1529}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1330 ( .s ({signal_4117, signal_4113}), .b ({signal_4125, signal_4123}), .a ({signal_2389, signal_1415}), .clk (CLK), .r (Fresh[202]), .c ({signal_2508, signal_1530}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1331 ( .s ({signal_4133, signal_4129}), .b ({signal_2390, signal_1416}), .a ({signal_4137, signal_4135}), .clk (CLK), .r (Fresh[203]), .c ({signal_2509, signal_1531}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1332 ( .s ({signal_4133, signal_4129}), .b ({signal_2391, signal_1417}), .a ({signal_4141, signal_4139}), .clk (CLK), .r (Fresh[204]), .c ({signal_2510, signal_1532}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1333 ( .s ({signal_4149, signal_4145}), .b ({signal_2392, signal_1418}), .a ({signal_4153, signal_4151}), .clk (CLK), .r (Fresh[205]), .c ({signal_2511, signal_1533}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1334 ( .s ({signal_4149, signal_4145}), .b ({signal_4157, signal_4155}), .a ({signal_2393, signal_1419}), .clk (CLK), .r (Fresh[206]), .c ({signal_2512, signal_1534}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1335 ( .s ({signal_4165, signal_4161}), .b ({signal_2394, signal_1420}), .a ({signal_4169, signal_4167}), .clk (CLK), .r (Fresh[207]), .c ({signal_2513, signal_1535}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1336 ( .s ({signal_4165, signal_4161}), .b ({signal_4173, signal_4171}), .a ({signal_2395, signal_1421}), .clk (CLK), .r (Fresh[208]), .c ({signal_2514, signal_1536}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1337 ( .s ({signal_4009, signal_4005}), .b ({signal_4177, signal_4175}), .a ({signal_2344, signal_1422}), .clk (CLK), .r (Fresh[209]), .c ({signal_2459, signal_1537}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1338 ( .s ({signal_4009, signal_4005}), .b ({signal_2346, signal_1424}), .a ({signal_2345, signal_1423}), .clk (CLK), .r (Fresh[210]), .c ({signal_2460, signal_1538}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1339 ( .s ({signal_4009, signal_4005}), .b ({signal_2344, signal_1422}), .a ({signal_4013, signal_4011}), .clk (CLK), .r (Fresh[211]), .c ({signal_2461, signal_1539}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1340 ( .s ({signal_4009, signal_4005}), .b ({signal_2334, signal_1396}), .a ({signal_4177, signal_4175}), .clk (CLK), .r (Fresh[212]), .c ({signal_2462, signal_1540}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1341 ( .s ({signal_4009, signal_4005}), .b ({signal_2348, signal_1426}), .a ({signal_2347, signal_1425}), .clk (CLK), .r (Fresh[213]), .c ({signal_2463, signal_1541}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1342 ( .s ({signal_4009, signal_4005}), .b ({signal_2344, signal_1422}), .a ({signal_4181, signal_4179}), .clk (CLK), .r (Fresh[214]), .c ({signal_2464, signal_1542}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1343 ( .s ({signal_4045, signal_4041}), .b ({signal_2350, signal_1428}), .a ({signal_2349, signal_1427}), .clk (CLK), .r (Fresh[215]), .c ({signal_2465, signal_1543}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1344 ( .s ({signal_4045, signal_4041}), .b ({signal_2351, signal_1429}), .a ({signal_4185, signal_4183}), .clk (CLK), .r (Fresh[216]), .c ({signal_2466, signal_1544}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1345 ( .s ({signal_4045, signal_4041}), .b ({signal_2351, signal_1429}), .a ({signal_4049, signal_4047}), .clk (CLK), .r (Fresh[217]), .c ({signal_2467, signal_1545}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1346 ( .s ({signal_4045, signal_4041}), .b ({signal_2343, signal_1405}), .a ({signal_4189, signal_4187}), .clk (CLK), .r (Fresh[218]), .c ({signal_2468, signal_1546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1347 ( .s ({signal_4021, signal_4017}), .b ({signal_2352, signal_1430}), .a ({signal_4025, signal_4023}), .clk (CLK), .r (Fresh[219]), .c ({signal_2469, signal_1547}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1348 ( .s ({signal_4021, signal_4017}), .b ({signal_2337, signal_1399}), .a ({signal_4193, signal_4191}), .clk (CLK), .r (Fresh[220]), .c ({signal_2470, signal_1548}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1349 ( .s ({signal_4021, signal_4017}), .b ({signal_2354, signal_1432}), .a ({signal_2353, signal_1431}), .clk (CLK), .r (Fresh[221]), .c ({signal_2471, signal_1549}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1350 ( .s ({signal_4021, signal_4017}), .b ({signal_2352, signal_1430}), .a ({signal_4197, signal_4195}), .clk (CLK), .r (Fresh[222]), .c ({signal_2472, signal_1550}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1351 ( .s ({signal_4149, signal_4145}), .b ({signal_2396, signal_1433}), .a ({signal_4157, signal_4155}), .clk (CLK), .r (Fresh[223]), .c ({signal_2515, signal_1551}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1352 ( .s ({signal_4149, signal_4145}), .b ({signal_2393, signal_1419}), .a ({signal_2397, signal_1434}), .clk (CLK), .r (Fresh[224]), .c ({signal_2516, signal_1552}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1353 ( .s ({signal_4021, signal_4017}), .b ({signal_4193, signal_4191}), .a ({signal_2352, signal_1430}), .clk (CLK), .r (Fresh[225]), .c ({signal_2473, signal_1553}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1354 ( .s ({signal_4021, signal_4017}), .b ({signal_2356, signal_1436}), .a ({signal_2355, signal_1435}), .clk (CLK), .r (Fresh[226]), .c ({signal_2474, signal_1554}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1355 ( .s ({signal_3997, signal_3993}), .b ({signal_4201, signal_4199}), .a ({signal_2357, signal_1437}), .clk (CLK), .r (Fresh[227]), .c ({signal_2475, signal_1555}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1356 ( .s ({signal_3997, signal_3993}), .b ({signal_2359, signal_1439}), .a ({signal_2358, signal_1438}), .clk (CLK), .r (Fresh[228]), .c ({signal_2476, signal_1556}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1357 ( .s ({signal_4117, signal_4113}), .b ({signal_2398, signal_1440}), .a ({signal_4125, signal_4123}), .clk (CLK), .r (Fresh[229]), .c ({signal_2517, signal_1557}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1358 ( .s ({signal_4117, signal_4113}), .b ({signal_2389, signal_1415}), .a ({signal_2399, signal_1441}), .clk (CLK), .r (Fresh[230]), .c ({signal_2518, signal_1558}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1359 ( .s ({signal_4133, signal_4129}), .b ({signal_4205, signal_4203}), .a ({signal_2391, signal_1417}), .clk (CLK), .r (Fresh[231]), .c ({signal_2519, signal_1559}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1360 ( .s ({signal_4133, signal_4129}), .b ({signal_4209, signal_4207}), .a ({signal_2390, signal_1416}), .clk (CLK), .r (Fresh[232]), .c ({signal_2520, signal_1560}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1361 ( .s ({signal_4089, signal_4085}), .b ({signal_4213, signal_4211}), .a ({signal_2385, signal_1411}), .clk (CLK), .r (Fresh[233]), .c ({signal_2521, signal_1561}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1362 ( .s ({signal_4089, signal_4085}), .b ({signal_4217, signal_4215}), .a ({signal_2384, signal_1410}), .clk (CLK), .r (Fresh[234]), .c ({signal_2522, signal_1562}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1363 ( .s ({signal_4033, signal_4029}), .b ({signal_2360, signal_1442}), .a ({signal_4037, signal_4035}), .clk (CLK), .r (Fresh[235]), .c ({signal_2477, signal_1563}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1364 ( .s ({signal_4033, signal_4029}), .b ({signal_2340, signal_1402}), .a ({signal_4221, signal_4219}), .clk (CLK), .r (Fresh[236]), .c ({signal_2478, signal_1564}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1365 ( .s ({signal_4101, signal_4099}), .b ({signal_2387, signal_1413}), .a ({signal_4105, signal_4103}), .clk (CLK), .r (Fresh[237]), .c ({signal_2523, signal_1565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1366 ( .s ({signal_4101, signal_4099}), .b ({signal_4225, signal_4223}), .a ({signal_2386, signal_1412}), .clk (CLK), .r (Fresh[238]), .c ({signal_2524, signal_1566}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1367 ( .s ({signal_4229, signal_4227}), .b ({signal_2401, signal_1444}), .a ({signal_2400, signal_1443}), .clk (CLK), .r (Fresh[239]), .c ({signal_2525, signal_1567}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1368 ( .s ({signal_4229, signal_4227}), .b ({signal_4225, signal_4223}), .a ({signal_2401, signal_1444}), .clk (CLK), .r (Fresh[240]), .c ({signal_2526, signal_1568}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1369 ( .s ({signal_4229, signal_4227}), .b ({signal_2400, signal_1443}), .a ({signal_4109, signal_4107}), .clk (CLK), .r (Fresh[241]), .c ({signal_2527, signal_1569}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1370 ( .s ({signal_4233, signal_4231}), .b ({signal_2402, signal_1445}), .a ({signal_2386, signal_1412}), .clk (CLK), .r (Fresh[242]), .c ({signal_2528, signal_1570}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1371 ( .s ({signal_4233, signal_4231}), .b ({signal_2386, signal_1412}), .a ({signal_2402, signal_1445}), .clk (CLK), .r (Fresh[243]), .c ({signal_2529, signal_1571}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1372 ( .s ({signal_4233, signal_4231}), .b ({signal_2404, signal_1447}), .a ({signal_2403, signal_1446}), .clk (CLK), .r (Fresh[244]), .c ({signal_2530, signal_1572}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1373 ( .s ({signal_4233, signal_4231}), .b ({signal_2403, signal_1446}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[245]), .c ({signal_2531, signal_1573}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1374 ( .s ({signal_4237, signal_4235}), .b ({signal_2406, signal_1449}), .a ({signal_2405, signal_1448}), .clk (CLK), .r (Fresh[246]), .c ({signal_2532, signal_1574}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1375 ( .s ({signal_4237, signal_4235}), .b ({signal_2405, signal_1448}), .a ({signal_2406, signal_1449}), .clk (CLK), .r (Fresh[247]), .c ({signal_2533, signal_1575}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1376 ( .s ({signal_4101, signal_4099}), .b ({signal_2406, signal_1449}), .a ({signal_2405, signal_1448}), .clk (CLK), .r (Fresh[248]), .c ({signal_2534, signal_1576}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1377 ( .s ({signal_4241, signal_4239}), .b ({signal_2406, signal_1449}), .a ({signal_2405, signal_1448}), .clk (CLK), .r (Fresh[249]), .c ({signal_2535, signal_1577}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1378 ( .s ({signal_4241, signal_4239}), .b ({signal_2405, signal_1448}), .a ({signal_2406, signal_1449}), .clk (CLK), .r (Fresh[250]), .c ({signal_2536, signal_1578}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1379 ( .s ({signal_4241, signal_4239}), .b ({signal_2403, signal_1446}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[251]), .c ({signal_2537, signal_1579}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1380 ( .s ({signal_4241, signal_4239}), .b ({signal_2404, signal_1447}), .a ({signal_2403, signal_1446}), .clk (CLK), .r (Fresh[252]), .c ({signal_2538, signal_1580}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1381 ( .s ({signal_4101, signal_4099}), .b ({signal_2408, signal_1451}), .a ({signal_2407, signal_1450}), .clk (CLK), .r (Fresh[253]), .c ({signal_2539, signal_1581}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1382 ( .s ({signal_4149, signal_4145}), .b ({signal_2393, signal_1419}), .a ({signal_4153, signal_4151}), .clk (CLK), .r (Fresh[254]), .c ({signal_2540, signal_1582}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1383 ( .s ({signal_4149, signal_4145}), .b ({signal_4245, signal_4243}), .a ({signal_2392, signal_1418}), .clk (CLK), .r (Fresh[255]), .c ({signal_2541, signal_1583}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1384 ( .s ({signal_3985, signal_3981}), .b ({signal_2361, signal_1452}), .a ({signal_4249, signal_4247}), .clk (CLK), .r (Fresh[256]), .c ({signal_2479, signal_1584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1385 ( .s ({signal_3985, signal_3981}), .b ({signal_2363, signal_1454}), .a ({signal_2362, signal_1453}), .clk (CLK), .r (Fresh[257]), .c ({signal_2480, signal_1585}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1386 ( .s ({signal_4149, signal_4145}), .b ({signal_4253, signal_4251}), .a ({signal_2396, signal_1433}), .clk (CLK), .r (Fresh[258]), .c ({signal_2542, signal_1586}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1387 ( .s ({signal_4149, signal_4145}), .b ({signal_4153, signal_4151}), .a ({signal_2409, signal_1455}), .clk (CLK), .r (Fresh[259]), .c ({signal_2543, signal_1587}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1388 ( .s ({signal_4073, signal_4069}), .b ({signal_2383, signal_1409}), .a ({signal_4077, signal_4075}), .clk (CLK), .r (Fresh[260]), .c ({signal_2544, signal_1588}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1389 ( .s ({signal_4073, signal_4069}), .b ({signal_4257, signal_4255}), .a ({signal_2382, signal_1408}), .clk (CLK), .r (Fresh[261]), .c ({signal_2545, signal_1589}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1390 ( .s ({signal_4117, signal_4113}), .b ({signal_2389, signal_1415}), .a ({signal_4121, signal_4119}), .clk (CLK), .r (Fresh[262]), .c ({signal_2546, signal_1590}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1391 ( .s ({signal_4117, signal_4113}), .b ({signal_4261, signal_4259}), .a ({signal_2388, signal_1414}), .clk (CLK), .r (Fresh[263]), .c ({signal_2547, signal_1591}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1392 ( .s ({signal_4165, signal_4161}), .b ({signal_2395, signal_1421}), .a ({signal_4169, signal_4167}), .clk (CLK), .r (Fresh[264]), .c ({signal_2548, signal_1592}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1393 ( .s ({signal_4165, signal_4161}), .b ({signal_4265, signal_4263}), .a ({signal_2394, signal_1420}), .clk (CLK), .r (Fresh[265]), .c ({signal_2549, signal_1593}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1394 ( .s ({signal_4117, signal_4113}), .b ({signal_4269, signal_4267}), .a ({signal_2398, signal_1440}), .clk (CLK), .r (Fresh[266]), .c ({signal_2550, signal_1594}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1395 ( .s ({signal_4117, signal_4113}), .b ({signal_4121, signal_4119}), .a ({signal_2410, signal_1456}), .clk (CLK), .r (Fresh[267]), .c ({signal_2551, signal_1595}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1396 ( .s ({signal_3961, signal_3957}), .b ({signal_2365, signal_1458}), .a ({signal_2364, signal_1457}), .clk (CLK), .r (Fresh[268]), .c ({signal_2481, signal_1596}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1397 ( .s ({signal_3961, signal_3957}), .b ({signal_2366, signal_1459}), .a ({signal_4273, signal_4271}), .clk (CLK), .r (Fresh[269]), .c ({signal_2482, signal_1597}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1398 ( .s ({signal_4165, signal_4161}), .b ({signal_2411, signal_1460}), .a ({signal_4173, signal_4171}), .clk (CLK), .r (Fresh[270]), .c ({signal_2552, signal_1598}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1399 ( .s ({signal_4165, signal_4161}), .b ({signal_2395, signal_1421}), .a ({signal_2412, signal_1461}), .clk (CLK), .r (Fresh[271]), .c ({signal_2553, signal_1599}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1400 ( .s ({signal_4117, signal_4113}), .b ({signal_2399, signal_1441}), .a ({signal_4269, signal_4267}), .clk (CLK), .r (Fresh[272]), .c ({signal_2554, signal_1600}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1401 ( .s ({signal_4117, signal_4113}), .b ({signal_4125, signal_4123}), .a ({signal_2413, signal_1462}), .clk (CLK), .r (Fresh[273]), .c ({signal_2555, signal_1601}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1402 ( .s ({signal_4165, signal_4161}), .b ({signal_4277, signal_4275}), .a ({signal_2411, signal_1460}), .clk (CLK), .r (Fresh[274]), .c ({signal_2556, signal_1602}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1403 ( .s ({signal_4165, signal_4161}), .b ({signal_4169, signal_4167}), .a ({signal_2414, signal_1463}), .clk (CLK), .r (Fresh[275]), .c ({signal_2557, signal_1603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1404 ( .s ({signal_3961, signal_3957}), .b ({signal_4281, signal_4279}), .a ({signal_2366, signal_1459}), .clk (CLK), .r (Fresh[276]), .c ({signal_2483, signal_1604}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1405 ( .s ({signal_3961, signal_3957}), .b ({signal_2368, signal_1465}), .a ({signal_2367, signal_1464}), .clk (CLK), .r (Fresh[277]), .c ({signal_2484, signal_1605}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1406 ( .s ({signal_4133, signal_4129}), .b ({signal_2416, signal_1467}), .a ({signal_2415, signal_1466}), .clk (CLK), .r (Fresh[278]), .c ({signal_2558, signal_1606}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1407 ( .s ({signal_4133, signal_4129}), .b ({signal_2415, signal_1466}), .a ({signal_2416, signal_1467}), .clk (CLK), .r (Fresh[279]), .c ({signal_2559, signal_1607}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1408 ( .s ({signal_3973, signal_3969}), .b ({signal_2370, signal_1469}), .a ({signal_2369, signal_1468}), .clk (CLK), .r (Fresh[280]), .c ({signal_2485, signal_1608}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1409 ( .s ({signal_3973, signal_3969}), .b ({signal_2371, signal_1470}), .a ({signal_4285, signal_4283}), .clk (CLK), .r (Fresh[281]), .c ({signal_2486, signal_1609}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1410 ( .s ({signal_4133, signal_4129}), .b ({signal_2417, signal_1471}), .a ({signal_4141, signal_4139}), .clk (CLK), .r (Fresh[282]), .c ({signal_2560, signal_1610}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1411 ( .s ({signal_4133, signal_4129}), .b ({signal_4205, signal_4203}), .a ({signal_2418, signal_1472}), .clk (CLK), .r (Fresh[283]), .c ({signal_2561, signal_1611}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1412 ( .s ({signal_4033, signal_4029}), .b ({signal_2373, signal_1474}), .a ({signal_2372, signal_1473}), .clk (CLK), .r (Fresh[284]), .c ({signal_2487, signal_1612}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1413 ( .s ({signal_4033, signal_4029}), .b ({signal_2360, signal_1442}), .a ({signal_4289, signal_4287}), .clk (CLK), .r (Fresh[285]), .c ({signal_2488, signal_1613}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1414 ( .s ({signal_4293, signal_4291}), .b ({signal_2419, signal_1475}), .a ({signal_4217, signal_4215}), .clk (CLK), .r (Fresh[286]), .c ({signal_2562, signal_1614}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1415 ( .s ({signal_4297, signal_4295}), .b ({signal_2421, signal_1477}), .a ({signal_2422, signal_1478}), .clk (CLK), .r (Fresh[287]), .c ({signal_2563, signal_1615}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1416 ( .s ({signal_4293, signal_4291}), .b ({signal_2421, signal_1477}), .a ({signal_2422, signal_1478}), .clk (CLK), .r (Fresh[288]), .c ({signal_2564, signal_1616}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1417 ( .s ({signal_4297, signal_4295}), .b ({signal_2422, signal_1478}), .a ({signal_2421, signal_1477}), .clk (CLK), .r (Fresh[289]), .c ({signal_2565, signal_1617}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1418 ( .s ({signal_4293, signal_4291}), .b ({signal_2422, signal_1478}), .a ({signal_2421, signal_1477}), .clk (CLK), .r (Fresh[290]), .c ({signal_2566, signal_1618}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1419 ( .s ({signal_4293, signal_4291}), .b ({signal_2423, signal_1479}), .a ({signal_4093, signal_4091}), .clk (CLK), .r (Fresh[291]), .c ({signal_2567, signal_1619}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1420 ( .s ({signal_4293, signal_4291}), .b ({signal_2425, signal_1481}), .a ({signal_4097, signal_4095}), .clk (CLK), .r (Fresh[292]), .c ({signal_2568, signal_1620}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1421 ( .s ({signal_4293, signal_4291}), .b ({signal_2426, signal_1482}), .a ({signal_4213, signal_4211}), .clk (CLK), .r (Fresh[293]), .c ({signal_2569, signal_1621}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1422 ( .s ({signal_4045, signal_4041}), .b ({signal_4189, signal_4187}), .a ({signal_2351, signal_1429}), .clk (CLK), .r (Fresh[294]), .c ({signal_2489, signal_1622}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1423 ( .s ({signal_4045, signal_4041}), .b ({signal_2375, signal_1484}), .a ({signal_2374, signal_1483}), .clk (CLK), .r (Fresh[295]), .c ({signal_2490, signal_1623}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1424 ( .s ({signal_4057, signal_4053}), .b ({signal_2427, signal_1485}), .a ({signal_4065, signal_4063}), .clk (CLK), .r (Fresh[296]), .c ({signal_2570, signal_1624}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1425 ( .s ({signal_4057, signal_4053}), .b ({signal_4301, signal_4299}), .a ({signal_2428, signal_1486}), .clk (CLK), .r (Fresh[297]), .c ({signal_2571, signal_1625}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1426 ( .s ({signal_4309, signal_4305}), .b ({signal_2430, signal_1488}), .a ({signal_2429, signal_1487}), .clk (CLK), .r (Fresh[298]), .c ({signal_2572, signal_1626}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1427 ( .s ({signal_4309, signal_4305}), .b ({signal_2429, signal_1487}), .a ({signal_2430, signal_1488}), .clk (CLK), .r (Fresh[299]), .c ({signal_2573, signal_1627}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1428 ( .s ({signal_4057, signal_4053}), .b ({signal_4301, signal_4299}), .a ({signal_2381, signal_1407}), .clk (CLK), .r (Fresh[300]), .c ({signal_2574, signal_1628}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1429 ( .s ({signal_4057, signal_4053}), .b ({signal_4313, signal_4311}), .a ({signal_2380, signal_1406}), .clk (CLK), .r (Fresh[301]), .c ({signal_2575, signal_1629}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1430 ( .s ({signal_4073, signal_4069}), .b ({signal_2431, signal_1489}), .a ({signal_4081, signal_4079}), .clk (CLK), .r (Fresh[302]), .c ({signal_2576, signal_1630}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1431 ( .s ({signal_4073, signal_4069}), .b ({signal_2383, signal_1409}), .a ({signal_2432, signal_1490}), .clk (CLK), .r (Fresh[303]), .c ({signal_2577, signal_1631}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1432 ( .s ({signal_4317, signal_4315}), .b ({signal_2397, signal_1434}), .a ({signal_2393, signal_1419}), .clk (CLK), .r (Fresh[304]), .c ({signal_2578, signal_1632}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1433 ( .s ({signal_4317, signal_4315}), .b ({signal_2434, signal_1492}), .a ({signal_2392, signal_1418}), .clk (CLK), .r (Fresh[305]), .c ({signal_2579, signal_1633}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1434 ( .s ({signal_4317, signal_4315}), .b ({signal_2393, signal_1419}), .a ({signal_2397, signal_1434}), .clk (CLK), .r (Fresh[306]), .c ({signal_2580, signal_1634}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1435 ( .s ({signal_4317, signal_4315}), .b ({signal_2392, signal_1418}), .a ({signal_2434, signal_1492}), .clk (CLK), .r (Fresh[307]), .c ({signal_2581, signal_1635}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1436 ( .s ({signal_4073, signal_4069}), .b ({signal_2438, signal_1496}), .a ({signal_4257, signal_4255}), .clk (CLK), .r (Fresh[308]), .c ({signal_2582, signal_1636}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1437 ( .s ({signal_4073, signal_4069}), .b ({signal_2432, signal_1490}), .a ({signal_2383, signal_1409}), .clk (CLK), .r (Fresh[309]), .c ({signal_2583, signal_1637}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1438 ( .s ({signal_4165, signal_4161}), .b ({signal_2412, signal_1461}), .a ({signal_4277, signal_4275}), .clk (CLK), .r (Fresh[310]), .c ({signal_2584, signal_1638}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1439 ( .s ({signal_4165, signal_4161}), .b ({signal_4173, signal_4171}), .a ({signal_2439, signal_1497}), .clk (CLK), .r (Fresh[311]), .c ({signal_2585, signal_1639}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1440 ( .s ({signal_3997, signal_3993}), .b ({signal_2357, signal_1437}), .a ({signal_4001, signal_3999}), .clk (CLK), .r (Fresh[312]), .c ({signal_2491, signal_1640}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1441 ( .s ({signal_3997, signal_3993}), .b ({signal_2331, signal_1393}), .a ({signal_4201, signal_4199}), .clk (CLK), .r (Fresh[313]), .c ({signal_2492, signal_1641}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1442 ( .s ({signal_4033, signal_4029}), .b ({signal_4221, signal_4219}), .a ({signal_2360, signal_1442}), .clk (CLK), .r (Fresh[314]), .c ({signal_2493, signal_1642}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1443 ( .s ({signal_4033, signal_4029}), .b ({signal_2377, signal_1499}), .a ({signal_2376, signal_1498}), .clk (CLK), .r (Fresh[315]), .c ({signal_2494, signal_1643}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1444 ( .s ({signal_4325, signal_4321}), .b ({signal_2441, signal_1501}), .a ({signal_2440, signal_1500}), .clk (CLK), .r (Fresh[316]), .c ({signal_2586, signal_1644}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1445 ( .s ({signal_4325, signal_4321}), .b ({signal_2440, signal_1500}), .a ({signal_2441, signal_1501}), .clk (CLK), .r (Fresh[317]), .c ({signal_2587, signal_1645}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1446 ( .s ({signal_4329, signal_4327}), .b ({signal_2441, signal_1501}), .a ({signal_2440, signal_1500}), .clk (CLK), .r (Fresh[318]), .c ({signal_2588, signal_1646}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1447 ( .s ({signal_4329, signal_4327}), .b ({signal_2440, signal_1500}), .a ({signal_2441, signal_1501}), .clk (CLK), .r (Fresh[319]), .c ({signal_2589, signal_1647}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1448 ( .s ({signal_3973, signal_3969}), .b ({signal_4333, signal_4331}), .a ({signal_2371, signal_1470}), .clk (CLK), .r (Fresh[320]), .c ({signal_2495, signal_1648}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1449 ( .s ({signal_3973, signal_3969}), .b ({signal_2379, signal_1503}), .a ({signal_2378, signal_1502}), .clk (CLK), .r (Fresh[321]), .c ({signal_2496, signal_1649}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1450 ( .s ({signal_4089, signal_4085}), .b ({signal_2441, signal_1501}), .a ({signal_2440, signal_1500}), .clk (CLK), .r (Fresh[322]), .c ({signal_2590, signal_1650}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1451 ( .s ({signal_4089, signal_4085}), .b ({signal_2440, signal_1500}), .a ({signal_2441, signal_1501}), .clk (CLK), .r (Fresh[323]), .c ({signal_2591, signal_1651}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1452 ( .s ({signal_4101, signal_4099}), .b ({signal_2403, signal_1446}), .a ({signal_2404, signal_1447}), .clk (CLK), .r (Fresh[324]), .c ({signal_2592, signal_1652}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1453 ( .s ({signal_4229, signal_4227}), .b ({signal_2400, signal_1443}), .a ({signal_2401, signal_1444}), .clk (CLK), .r (Fresh[325]), .c ({signal_2593, signal_1653}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1454 ( .s ({signal_3985, signal_3981}), .b ({signal_3989, signal_3987}), .a ({signal_2361, signal_1452}), .clk (CLK), .r (Fresh[326]), .c ({signal_2497, signal_1654}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1455 ( .s ({signal_3985, signal_3981}), .b ({signal_4249, signal_4247}), .a ({signal_2328, signal_1390}), .clk (CLK), .r (Fresh[327]), .c ({signal_2498, signal_1655}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1456 ( .s ({signal_4293, signal_4291}), .b ({signal_4097, signal_4095}), .a ({signal_2419, signal_1475}), .clk (CLK), .r (Fresh[328]), .c ({signal_2594, signal_1656}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1457 ( .s ({signal_4293, signal_4291}), .b ({signal_4217, signal_4215}), .a ({signal_2425, signal_1481}), .clk (CLK), .r (Fresh[329]), .c ({signal_2595, signal_1657}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1458 ( .s ({signal_4293, signal_4291}), .b ({signal_4213, signal_4211}), .a ({signal_2423, signal_1479}), .clk (CLK), .r (Fresh[330]), .c ({signal_2596, signal_1658}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1459 ( .s ({signal_4293, signal_4291}), .b ({signal_4093, signal_4091}), .a ({signal_2426, signal_1482}), .clk (CLK), .r (Fresh[331]), .c ({signal_2597, signal_1659}) ) ;
    buf_clk cell_2195 ( .C (CLK), .D (signal_4338), .Q (signal_4339) ) ;
    buf_clk cell_2203 ( .C (CLK), .D (signal_4346), .Q (signal_4347) ) ;
    buf_clk cell_2211 ( .C (CLK), .D (signal_4354), .Q (signal_4355) ) ;
    buf_clk cell_2219 ( .C (CLK), .D (signal_4362), .Q (signal_4363) ) ;
    buf_clk cell_2227 ( .C (CLK), .D (signal_4370), .Q (signal_4371) ) ;
    buf_clk cell_2235 ( .C (CLK), .D (signal_4378), .Q (signal_4379) ) ;
    buf_clk cell_2243 ( .C (CLK), .D (signal_4386), .Q (signal_4387) ) ;
    buf_clk cell_2251 ( .C (CLK), .D (signal_4394), .Q (signal_4395) ) ;
    buf_clk cell_2259 ( .C (CLK), .D (signal_4402), .Q (signal_4403) ) ;
    buf_clk cell_2267 ( .C (CLK), .D (signal_4410), .Q (signal_4411) ) ;
    buf_clk cell_2271 ( .C (CLK), .D (signal_4414), .Q (signal_4415) ) ;
    buf_clk cell_2275 ( .C (CLK), .D (signal_4418), .Q (signal_4419) ) ;
    buf_clk cell_2283 ( .C (CLK), .D (signal_4426), .Q (signal_4427) ) ;
    buf_clk cell_2291 ( .C (CLK), .D (signal_4434), .Q (signal_4435) ) ;
    buf_clk cell_2295 ( .C (CLK), .D (signal_4438), .Q (signal_4439) ) ;
    buf_clk cell_2299 ( .C (CLK), .D (signal_4442), .Q (signal_4443) ) ;
    buf_clk cell_2303 ( .C (CLK), .D (signal_4446), .Q (signal_4447) ) ;
    buf_clk cell_2307 ( .C (CLK), .D (signal_4450), .Q (signal_4451) ) ;
    buf_clk cell_2315 ( .C (CLK), .D (signal_4458), .Q (signal_4459) ) ;
    buf_clk cell_2323 ( .C (CLK), .D (signal_4466), .Q (signal_4467) ) ;
    buf_clk cell_2331 ( .C (CLK), .D (signal_4474), .Q (signal_4475) ) ;
    buf_clk cell_2339 ( .C (CLK), .D (signal_4482), .Q (signal_4483) ) ;
    buf_clk cell_2343 ( .C (CLK), .D (signal_4486), .Q (signal_4487) ) ;
    buf_clk cell_2347 ( .C (CLK), .D (signal_4490), .Q (signal_4491) ) ;
    buf_clk cell_2355 ( .C (CLK), .D (signal_4498), .Q (signal_4499) ) ;
    buf_clk cell_2361 ( .C (CLK), .D (signal_4504), .Q (signal_4505) ) ;
    buf_clk cell_2367 ( .C (CLK), .D (signal_4510), .Q (signal_4511) ) ;
    buf_clk cell_2375 ( .C (CLK), .D (signal_4518), .Q (signal_4519) ) ;
    buf_clk cell_2383 ( .C (CLK), .D (signal_4526), .Q (signal_4527) ) ;
    buf_clk cell_2391 ( .C (CLK), .D (signal_4534), .Q (signal_4535) ) ;
    buf_clk cell_2399 ( .C (CLK), .D (signal_4542), .Q (signal_4543) ) ;
    buf_clk cell_2407 ( .C (CLK), .D (signal_4550), .Q (signal_4551) ) ;
    buf_clk cell_2415 ( .C (CLK), .D (signal_4558), .Q (signal_4559) ) ;
    buf_clk cell_2423 ( .C (CLK), .D (signal_4566), .Q (signal_4567) ) ;
    buf_clk cell_2431 ( .C (CLK), .D (signal_4574), .Q (signal_4575) ) ;
    buf_clk cell_2439 ( .C (CLK), .D (signal_4582), .Q (signal_4583) ) ;
    buf_clk cell_2447 ( .C (CLK), .D (signal_4590), .Q (signal_4591) ) ;
    buf_clk cell_2455 ( .C (CLK), .D (signal_4598), .Q (signal_4599) ) ;
    buf_clk cell_2463 ( .C (CLK), .D (signal_4606), .Q (signal_4607) ) ;
    buf_clk cell_2471 ( .C (CLK), .D (signal_4614), .Q (signal_4615) ) ;
    buf_clk cell_2479 ( .C (CLK), .D (signal_4622), .Q (signal_4623) ) ;
    buf_clk cell_2487 ( .C (CLK), .D (signal_4630), .Q (signal_4631) ) ;
    buf_clk cell_2495 ( .C (CLK), .D (signal_4638), .Q (signal_4639) ) ;
    buf_clk cell_2503 ( .C (CLK), .D (signal_4646), .Q (signal_4647) ) ;
    buf_clk cell_2511 ( .C (CLK), .D (signal_4654), .Q (signal_4655) ) ;
    buf_clk cell_2519 ( .C (CLK), .D (signal_4662), .Q (signal_4663) ) ;
    buf_clk cell_2527 ( .C (CLK), .D (signal_4670), .Q (signal_4671) ) ;
    buf_clk cell_2535 ( .C (CLK), .D (signal_4678), .Q (signal_4679) ) ;
    buf_clk cell_2543 ( .C (CLK), .D (signal_4686), .Q (signal_4687) ) ;
    buf_clk cell_2551 ( .C (CLK), .D (signal_4694), .Q (signal_4695) ) ;
    buf_clk cell_2559 ( .C (CLK), .D (signal_4702), .Q (signal_4703) ) ;
    buf_clk cell_2567 ( .C (CLK), .D (signal_4710), .Q (signal_4711) ) ;
    buf_clk cell_2571 ( .C (CLK), .D (signal_4714), .Q (signal_4715) ) ;
    buf_clk cell_2575 ( .C (CLK), .D (signal_4718), .Q (signal_4719) ) ;
    buf_clk cell_2579 ( .C (CLK), .D (signal_4722), .Q (signal_4723) ) ;
    buf_clk cell_2583 ( .C (CLK), .D (signal_4726), .Q (signal_4727) ) ;
    buf_clk cell_2591 ( .C (CLK), .D (signal_4734), .Q (signal_4735) ) ;
    buf_clk cell_2599 ( .C (CLK), .D (signal_4742), .Q (signal_4743) ) ;
    buf_clk cell_2607 ( .C (CLK), .D (signal_4750), .Q (signal_4751) ) ;
    buf_clk cell_2615 ( .C (CLK), .D (signal_4758), .Q (signal_4759) ) ;
    buf_clk cell_2619 ( .C (CLK), .D (signal_4762), .Q (signal_4763) ) ;
    buf_clk cell_2623 ( .C (CLK), .D (signal_4766), .Q (signal_4767) ) ;
    buf_clk cell_2629 ( .C (CLK), .D (signal_4772), .Q (signal_4773) ) ;
    buf_clk cell_2635 ( .C (CLK), .D (signal_4778), .Q (signal_4779) ) ;
    buf_clk cell_2643 ( .C (CLK), .D (signal_4786), .Q (signal_4787) ) ;
    buf_clk cell_2651 ( .C (CLK), .D (signal_4794), .Q (signal_4795) ) ;
    buf_clk cell_2659 ( .C (CLK), .D (signal_4802), .Q (signal_4803) ) ;
    buf_clk cell_2667 ( .C (CLK), .D (signal_4810), .Q (signal_4811) ) ;
    buf_clk cell_2673 ( .C (CLK), .D (signal_4816), .Q (signal_4817) ) ;
    buf_clk cell_2679 ( .C (CLK), .D (signal_4822), .Q (signal_4823) ) ;
    buf_clk cell_2683 ( .C (CLK), .D (signal_4826), .Q (signal_4827) ) ;
    buf_clk cell_2687 ( .C (CLK), .D (signal_4830), .Q (signal_4831) ) ;
    buf_clk cell_2695 ( .C (CLK), .D (signal_4838), .Q (signal_4839) ) ;
    buf_clk cell_2703 ( .C (CLK), .D (signal_4846), .Q (signal_4847) ) ;
    buf_clk cell_2711 ( .C (CLK), .D (signal_4854), .Q (signal_4855) ) ;
    buf_clk cell_2719 ( .C (CLK), .D (signal_4862), .Q (signal_4863) ) ;
    buf_clk cell_2727 ( .C (CLK), .D (signal_4870), .Q (signal_4871) ) ;
    buf_clk cell_2735 ( .C (CLK), .D (signal_4878), .Q (signal_4879) ) ;
    buf_clk cell_2743 ( .C (CLK), .D (signal_4886), .Q (signal_4887) ) ;
    buf_clk cell_2751 ( .C (CLK), .D (signal_4894), .Q (signal_4895) ) ;
    buf_clk cell_2759 ( .C (CLK), .D (signal_4902), .Q (signal_4903) ) ;
    buf_clk cell_2767 ( .C (CLK), .D (signal_4910), .Q (signal_4911) ) ;
    buf_clk cell_2775 ( .C (CLK), .D (signal_4918), .Q (signal_4919) ) ;
    buf_clk cell_2783 ( .C (CLK), .D (signal_4926), .Q (signal_4927) ) ;
    buf_clk cell_2791 ( .C (CLK), .D (signal_4934), .Q (signal_4935) ) ;
    buf_clk cell_2797 ( .C (CLK), .D (signal_4940), .Q (signal_4941) ) ;
    buf_clk cell_2803 ( .C (CLK), .D (signal_4946), .Q (signal_4947) ) ;
    buf_clk cell_2809 ( .C (CLK), .D (signal_4952), .Q (signal_4953) ) ;
    buf_clk cell_2815 ( .C (CLK), .D (signal_4958), .Q (signal_4959) ) ;
    buf_clk cell_2821 ( .C (CLK), .D (signal_4964), .Q (signal_4965) ) ;
    buf_clk cell_2827 ( .C (CLK), .D (signal_4970), .Q (signal_4971) ) ;
    buf_clk cell_2833 ( .C (CLK), .D (signal_4976), .Q (signal_4977) ) ;
    buf_clk cell_2839 ( .C (CLK), .D (signal_4982), .Q (signal_4983) ) ;
    buf_clk cell_2845 ( .C (CLK), .D (signal_4988), .Q (signal_4989) ) ;
    buf_clk cell_2851 ( .C (CLK), .D (signal_4994), .Q (signal_4995) ) ;
    buf_clk cell_2857 ( .C (CLK), .D (signal_5000), .Q (signal_5001) ) ;
    buf_clk cell_2863 ( .C (CLK), .D (signal_5006), .Q (signal_5007) ) ;
    buf_clk cell_2869 ( .C (CLK), .D (signal_5012), .Q (signal_5013) ) ;
    buf_clk cell_2871 ( .C (CLK), .D (signal_5014), .Q (signal_5015) ) ;
    buf_clk cell_2873 ( .C (CLK), .D (signal_5016), .Q (signal_5017) ) ;
    buf_clk cell_2875 ( .C (CLK), .D (signal_5018), .Q (signal_5019) ) ;
    buf_clk cell_2877 ( .C (CLK), .D (signal_5020), .Q (signal_5021) ) ;
    buf_clk cell_2879 ( .C (CLK), .D (signal_5022), .Q (signal_5023) ) ;
    buf_clk cell_2881 ( .C (CLK), .D (signal_5024), .Q (signal_5025) ) ;
    buf_clk cell_2883 ( .C (CLK), .D (signal_5026), .Q (signal_5027) ) ;
    buf_clk cell_2885 ( .C (CLK), .D (signal_5028), .Q (signal_5029) ) ;
    buf_clk cell_2887 ( .C (CLK), .D (signal_5030), .Q (signal_5031) ) ;
    buf_clk cell_2889 ( .C (CLK), .D (signal_5032), .Q (signal_5033) ) ;
    buf_clk cell_2891 ( .C (CLK), .D (signal_5034), .Q (signal_5035) ) ;
    buf_clk cell_2893 ( .C (CLK), .D (signal_5036), .Q (signal_5037) ) ;
    buf_clk cell_2895 ( .C (CLK), .D (signal_5038), .Q (signal_5039) ) ;
    buf_clk cell_2897 ( .C (CLK), .D (signal_5040), .Q (signal_5041) ) ;
    buf_clk cell_2899 ( .C (CLK), .D (signal_5042), .Q (signal_5043) ) ;
    buf_clk cell_2901 ( .C (CLK), .D (signal_5044), .Q (signal_5045) ) ;
    buf_clk cell_2903 ( .C (CLK), .D (signal_5046), .Q (signal_5047) ) ;
    buf_clk cell_2905 ( .C (CLK), .D (signal_5048), .Q (signal_5049) ) ;
    buf_clk cell_2907 ( .C (CLK), .D (signal_5050), .Q (signal_5051) ) ;
    buf_clk cell_2909 ( .C (CLK), .D (signal_5052), .Q (signal_5053) ) ;
    buf_clk cell_2911 ( .C (CLK), .D (signal_5054), .Q (signal_5055) ) ;
    buf_clk cell_2913 ( .C (CLK), .D (signal_5056), .Q (signal_5057) ) ;
    buf_clk cell_2915 ( .C (CLK), .D (signal_5058), .Q (signal_5059) ) ;
    buf_clk cell_2917 ( .C (CLK), .D (signal_5060), .Q (signal_5061) ) ;
    buf_clk cell_2919 ( .C (CLK), .D (signal_5062), .Q (signal_5063) ) ;
    buf_clk cell_2921 ( .C (CLK), .D (signal_5064), .Q (signal_5065) ) ;
    buf_clk cell_2923 ( .C (CLK), .D (signal_5066), .Q (signal_5067) ) ;
    buf_clk cell_2925 ( .C (CLK), .D (signal_5068), .Q (signal_5069) ) ;
    buf_clk cell_2927 ( .C (CLK), .D (signal_5070), .Q (signal_5071) ) ;
    buf_clk cell_2929 ( .C (CLK), .D (signal_5072), .Q (signal_5073) ) ;
    buf_clk cell_2931 ( .C (CLK), .D (signal_5074), .Q (signal_5075) ) ;
    buf_clk cell_2933 ( .C (CLK), .D (signal_5076), .Q (signal_5077) ) ;
    buf_clk cell_2937 ( .C (CLK), .D (signal_5080), .Q (signal_5081) ) ;
    buf_clk cell_2941 ( .C (CLK), .D (signal_5084), .Q (signal_5085) ) ;
    buf_clk cell_2943 ( .C (CLK), .D (signal_5086), .Q (signal_5087) ) ;
    buf_clk cell_2945 ( .C (CLK), .D (signal_5088), .Q (signal_5089) ) ;
    buf_clk cell_2947 ( .C (CLK), .D (signal_5090), .Q (signal_5091) ) ;
    buf_clk cell_2949 ( .C (CLK), .D (signal_5092), .Q (signal_5093) ) ;
    buf_clk cell_2951 ( .C (CLK), .D (signal_5094), .Q (signal_5095) ) ;
    buf_clk cell_2953 ( .C (CLK), .D (signal_5096), .Q (signal_5097) ) ;
    buf_clk cell_2955 ( .C (CLK), .D (signal_5098), .Q (signal_5099) ) ;
    buf_clk cell_2957 ( .C (CLK), .D (signal_5100), .Q (signal_5101) ) ;
    buf_clk cell_2959 ( .C (CLK), .D (signal_5102), .Q (signal_5103) ) ;
    buf_clk cell_2961 ( .C (CLK), .D (signal_5104), .Q (signal_5105) ) ;
    buf_clk cell_2963 ( .C (CLK), .D (signal_5106), .Q (signal_5107) ) ;
    buf_clk cell_2965 ( .C (CLK), .D (signal_5108), .Q (signal_5109) ) ;
    buf_clk cell_2967 ( .C (CLK), .D (signal_5110), .Q (signal_5111) ) ;
    buf_clk cell_2969 ( .C (CLK), .D (signal_5112), .Q (signal_5113) ) ;
    buf_clk cell_2975 ( .C (CLK), .D (signal_5118), .Q (signal_5119) ) ;
    buf_clk cell_2981 ( .C (CLK), .D (signal_5124), .Q (signal_5125) ) ;
    buf_clk cell_2985 ( .C (CLK), .D (signal_5128), .Q (signal_5129) ) ;
    buf_clk cell_2989 ( .C (CLK), .D (signal_5132), .Q (signal_5133) ) ;
    buf_clk cell_2991 ( .C (CLK), .D (signal_5134), .Q (signal_5135) ) ;
    buf_clk cell_2993 ( .C (CLK), .D (signal_5136), .Q (signal_5137) ) ;
    buf_clk cell_2995 ( .C (CLK), .D (signal_5138), .Q (signal_5139) ) ;
    buf_clk cell_2997 ( .C (CLK), .D (signal_5140), .Q (signal_5141) ) ;
    buf_clk cell_2999 ( .C (CLK), .D (signal_5142), .Q (signal_5143) ) ;
    buf_clk cell_3001 ( .C (CLK), .D (signal_5144), .Q (signal_5145) ) ;
    buf_clk cell_3003 ( .C (CLK), .D (signal_5146), .Q (signal_5147) ) ;
    buf_clk cell_3005 ( .C (CLK), .D (signal_5148), .Q (signal_5149) ) ;
    buf_clk cell_3007 ( .C (CLK), .D (signal_5150), .Q (signal_5151) ) ;
    buf_clk cell_3009 ( .C (CLK), .D (signal_5152), .Q (signal_5153) ) ;
    buf_clk cell_3017 ( .C (CLK), .D (signal_5160), .Q (signal_5161) ) ;
    buf_clk cell_3023 ( .C (CLK), .D (signal_5166), .Q (signal_5167) ) ;
    buf_clk cell_3059 ( .C (CLK), .D (signal_5202), .Q (signal_5203) ) ;
    buf_clk cell_3067 ( .C (CLK), .D (signal_5210), .Q (signal_5211) ) ;
    buf_clk cell_3087 ( .C (CLK), .D (signal_5230), .Q (signal_5231) ) ;
    buf_clk cell_3091 ( .C (CLK), .D (signal_5234), .Q (signal_5235) ) ;
    buf_clk cell_3197 ( .C (CLK), .D (signal_5340), .Q (signal_5341) ) ;
    buf_clk cell_3205 ( .C (CLK), .D (signal_5348), .Q (signal_5349) ) ;
    buf_clk cell_3319 ( .C (CLK), .D (signal_5462), .Q (signal_5463) ) ;
    buf_clk cell_3327 ( .C (CLK), .D (signal_5470), .Q (signal_5471) ) ;
    buf_clk cell_3355 ( .C (CLK), .D (signal_5498), .Q (signal_5499) ) ;
    buf_clk cell_3363 ( .C (CLK), .D (signal_5506), .Q (signal_5507) ) ;
    buf_clk cell_3451 ( .C (CLK), .D (signal_5594), .Q (signal_5595) ) ;
    buf_clk cell_3467 ( .C (CLK), .D (signal_5610), .Q (signal_5611) ) ;
    buf_clk cell_3491 ( .C (CLK), .D (signal_5634), .Q (signal_5635) ) ;
    buf_clk cell_3507 ( .C (CLK), .D (signal_5650), .Q (signal_5651) ) ;
    buf_clk cell_3531 ( .C (CLK), .D (signal_5674), .Q (signal_5675) ) ;
    buf_clk cell_3547 ( .C (CLK), .D (signal_5690), .Q (signal_5691) ) ;
    buf_clk cell_3563 ( .C (CLK), .D (signal_5706), .Q (signal_5707) ) ;
    buf_clk cell_3579 ( .C (CLK), .D (signal_5722), .Q (signal_5723) ) ;
    buf_clk cell_3639 ( .C (CLK), .D (signal_5782), .Q (signal_5783) ) ;
    buf_clk cell_3655 ( .C (CLK), .D (signal_5798), .Q (signal_5799) ) ;
    buf_clk cell_3671 ( .C (CLK), .D (signal_5814), .Q (signal_5815) ) ;
    buf_clk cell_3687 ( .C (CLK), .D (signal_5830), .Q (signal_5831) ) ;
    buf_clk cell_3703 ( .C (CLK), .D (signal_5846), .Q (signal_5847) ) ;
    buf_clk cell_3719 ( .C (CLK), .D (signal_5862), .Q (signal_5863) ) ;
    buf_clk cell_3735 ( .C (CLK), .D (signal_5878), .Q (signal_5879) ) ;
    buf_clk cell_3751 ( .C (CLK), .D (signal_5894), .Q (signal_5895) ) ;
    buf_clk cell_3767 ( .C (CLK), .D (signal_5910), .Q (signal_5911) ) ;
    buf_clk cell_3783 ( .C (CLK), .D (signal_5926), .Q (signal_5927) ) ;
    buf_clk cell_3891 ( .C (CLK), .D (signal_6034), .Q (signal_6035) ) ;
    buf_clk cell_3907 ( .C (CLK), .D (signal_6050), .Q (signal_6051) ) ;
    buf_clk cell_3923 ( .C (CLK), .D (signal_6066), .Q (signal_6067) ) ;
    buf_clk cell_3939 ( .C (CLK), .D (signal_6082), .Q (signal_6083) ) ;
    buf_clk cell_3955 ( .C (CLK), .D (signal_6098), .Q (signal_6099) ) ;
    buf_clk cell_3971 ( .C (CLK), .D (signal_6114), .Q (signal_6115) ) ;
    buf_clk cell_3987 ( .C (CLK), .D (signal_6130), .Q (signal_6131) ) ;
    buf_clk cell_4003 ( .C (CLK), .D (signal_6146), .Q (signal_6147) ) ;
    buf_clk cell_4019 ( .C (CLK), .D (signal_6162), .Q (signal_6163) ) ;
    buf_clk cell_4035 ( .C (CLK), .D (signal_6178), .Q (signal_6179) ) ;
    buf_clk cell_4051 ( .C (CLK), .D (signal_6194), .Q (signal_6195) ) ;
    buf_clk cell_4067 ( .C (CLK), .D (signal_6210), .Q (signal_6211) ) ;
    buf_clk cell_4083 ( .C (CLK), .D (signal_6226), .Q (signal_6227) ) ;
    buf_clk cell_4099 ( .C (CLK), .D (signal_6242), .Q (signal_6243) ) ;
    buf_clk cell_4183 ( .C (CLK), .D (signal_6326), .Q (signal_6327) ) ;
    buf_clk cell_4195 ( .C (CLK), .D (signal_6338), .Q (signal_6339) ) ;
    buf_clk cell_4207 ( .C (CLK), .D (signal_6350), .Q (signal_6351) ) ;
    buf_clk cell_4235 ( .C (CLK), .D (signal_6378), .Q (signal_6379) ) ;
    buf_clk cell_4247 ( .C (CLK), .D (signal_6390), .Q (signal_6391) ) ;
    buf_clk cell_4261 ( .C (CLK), .D (signal_6404), .Q (signal_6405) ) ;
    buf_clk cell_4275 ( .C (CLK), .D (signal_6418), .Q (signal_6419) ) ;
    buf_clk cell_4291 ( .C (CLK), .D (signal_6434), .Q (signal_6435) ) ;
    buf_clk cell_4307 ( .C (CLK), .D (signal_6450), .Q (signal_6451) ) ;
    buf_clk cell_4323 ( .C (CLK), .D (signal_6466), .Q (signal_6467) ) ;
    buf_clk cell_4339 ( .C (CLK), .D (signal_6482), .Q (signal_6483) ) ;
    buf_clk cell_4355 ( .C (CLK), .D (signal_6498), .Q (signal_6499) ) ;
    buf_clk cell_4371 ( .C (CLK), .D (signal_6514), .Q (signal_6515) ) ;
    buf_clk cell_4387 ( .C (CLK), .D (signal_6530), .Q (signal_6531) ) ;
    buf_clk cell_4403 ( .C (CLK), .D (signal_6546), .Q (signal_6547) ) ;
    buf_clk cell_4419 ( .C (CLK), .D (signal_6562), .Q (signal_6563) ) ;
    buf_clk cell_4435 ( .C (CLK), .D (signal_6578), .Q (signal_6579) ) ;
    buf_clk cell_4451 ( .C (CLK), .D (signal_6594), .Q (signal_6595) ) ;
    buf_clk cell_4467 ( .C (CLK), .D (signal_6610), .Q (signal_6611) ) ;
    buf_clk cell_4483 ( .C (CLK), .D (signal_6626), .Q (signal_6627) ) ;
    buf_clk cell_4499 ( .C (CLK), .D (signal_6642), .Q (signal_6643) ) ;
    buf_clk cell_4515 ( .C (CLK), .D (signal_6658), .Q (signal_6659) ) ;
    buf_clk cell_4531 ( .C (CLK), .D (signal_6674), .Q (signal_6675) ) ;
    buf_clk cell_4579 ( .C (CLK), .D (signal_6722), .Q (signal_6723) ) ;
    buf_clk cell_4591 ( .C (CLK), .D (signal_6734), .Q (signal_6735) ) ;
    buf_clk cell_4605 ( .C (CLK), .D (signal_6748), .Q (signal_6749) ) ;
    buf_clk cell_4619 ( .C (CLK), .D (signal_6762), .Q (signal_6763) ) ;
    buf_clk cell_4635 ( .C (CLK), .D (signal_6778), .Q (signal_6779) ) ;
    buf_clk cell_4651 ( .C (CLK), .D (signal_6794), .Q (signal_6795) ) ;
    buf_clk cell_4711 ( .C (CLK), .D (signal_6854), .Q (signal_6855) ) ;
    buf_clk cell_4723 ( .C (CLK), .D (signal_6866), .Q (signal_6867) ) ;
    buf_clk cell_4747 ( .C (CLK), .D (signal_6890), .Q (signal_6891) ) ;
    buf_clk cell_4763 ( .C (CLK), .D (signal_6906), .Q (signal_6907) ) ;
    buf_clk cell_4779 ( .C (CLK), .D (signal_6922), .Q (signal_6923) ) ;
    buf_clk cell_4795 ( .C (CLK), .D (signal_6938), .Q (signal_6939) ) ;
    buf_clk cell_4811 ( .C (CLK), .D (signal_6954), .Q (signal_6955) ) ;
    buf_clk cell_4827 ( .C (CLK), .D (signal_6970), .Q (signal_6971) ) ;
    buf_clk cell_4843 ( .C (CLK), .D (signal_6986), .Q (signal_6987) ) ;
    buf_clk cell_4859 ( .C (CLK), .D (signal_7002), .Q (signal_7003) ) ;
    buf_clk cell_4875 ( .C (CLK), .D (signal_7018), .Q (signal_7019) ) ;
    buf_clk cell_4891 ( .C (CLK), .D (signal_7034), .Q (signal_7035) ) ;
    buf_clk cell_4907 ( .C (CLK), .D (signal_7050), .Q (signal_7051) ) ;
    buf_clk cell_4923 ( .C (CLK), .D (signal_7066), .Q (signal_7067) ) ;
    buf_clk cell_4939 ( .C (CLK), .D (signal_7082), .Q (signal_7083) ) ;
    buf_clk cell_4955 ( .C (CLK), .D (signal_7098), .Q (signal_7099) ) ;
    buf_clk cell_4971 ( .C (CLK), .D (signal_7114), .Q (signal_7115) ) ;
    buf_clk cell_4987 ( .C (CLK), .D (signal_7130), .Q (signal_7131) ) ;
    buf_clk cell_5003 ( .C (CLK), .D (signal_7146), .Q (signal_7147) ) ;
    buf_clk cell_5019 ( .C (CLK), .D (signal_7162), .Q (signal_7163) ) ;
    buf_clk cell_5035 ( .C (CLK), .D (signal_7178), .Q (signal_7179) ) ;
    buf_clk cell_5051 ( .C (CLK), .D (signal_7194), .Q (signal_7195) ) ;
    buf_clk cell_5067 ( .C (CLK), .D (signal_7210), .Q (signal_7211) ) ;
    buf_clk cell_5083 ( .C (CLK), .D (signal_7226), .Q (signal_7227) ) ;
    buf_clk cell_5099 ( .C (CLK), .D (signal_7242), .Q (signal_7243) ) ;
    buf_clk cell_5115 ( .C (CLK), .D (signal_7258), .Q (signal_7259) ) ;
    buf_clk cell_5131 ( .C (CLK), .D (signal_7274), .Q (signal_7275) ) ;
    buf_clk cell_5147 ( .C (CLK), .D (signal_7290), .Q (signal_7291) ) ;
    buf_clk cell_5163 ( .C (CLK), .D (signal_7306), .Q (signal_7307) ) ;
    buf_clk cell_5179 ( .C (CLK), .D (signal_7322), .Q (signal_7323) ) ;
    buf_clk cell_5195 ( .C (CLK), .D (signal_7338), .Q (signal_7339) ) ;
    buf_clk cell_5211 ( .C (CLK), .D (signal_7354), .Q (signal_7355) ) ;
    buf_clk cell_5227 ( .C (CLK), .D (signal_7370), .Q (signal_7371) ) ;
    buf_clk cell_5243 ( .C (CLK), .D (signal_7386), .Q (signal_7387) ) ;
    buf_clk cell_5259 ( .C (CLK), .D (signal_7402), .Q (signal_7403) ) ;
    buf_clk cell_5275 ( .C (CLK), .D (signal_7418), .Q (signal_7419) ) ;
    buf_clk cell_5291 ( .C (CLK), .D (signal_7434), .Q (signal_7435) ) ;
    buf_clk cell_5307 ( .C (CLK), .D (signal_7450), .Q (signal_7451) ) ;
    buf_clk cell_5323 ( .C (CLK), .D (signal_7466), .Q (signal_7467) ) ;
    buf_clk cell_5339 ( .C (CLK), .D (signal_7482), .Q (signal_7483) ) ;
    buf_clk cell_5355 ( .C (CLK), .D (signal_7498), .Q (signal_7499) ) ;
    buf_clk cell_5371 ( .C (CLK), .D (signal_7514), .Q (signal_7515) ) ;
    buf_clk cell_5387 ( .C (CLK), .D (signal_7530), .Q (signal_7531) ) ;
    buf_clk cell_5403 ( .C (CLK), .D (signal_7546), .Q (signal_7547) ) ;
    buf_clk cell_5419 ( .C (CLK), .D (signal_7562), .Q (signal_7563) ) ;
    buf_clk cell_5435 ( .C (CLK), .D (signal_7578), .Q (signal_7579) ) ;
    buf_clk cell_5451 ( .C (CLK), .D (signal_7594), .Q (signal_7595) ) ;
    buf_clk cell_5467 ( .C (CLK), .D (signal_7610), .Q (signal_7611) ) ;
    buf_clk cell_5483 ( .C (CLK), .D (signal_7626), .Q (signal_7627) ) ;
    buf_clk cell_5499 ( .C (CLK), .D (signal_7642), .Q (signal_7643) ) ;
    buf_clk cell_5515 ( .C (CLK), .D (signal_7658), .Q (signal_7659) ) ;
    buf_clk cell_5531 ( .C (CLK), .D (signal_7674), .Q (signal_7675) ) ;
    buf_clk cell_5547 ( .C (CLK), .D (signal_7690), .Q (signal_7691) ) ;
    buf_clk cell_5563 ( .C (CLK), .D (signal_7706), .Q (signal_7707) ) ;
    buf_clk cell_5579 ( .C (CLK), .D (signal_7722), .Q (signal_7723) ) ;
    buf_clk cell_5595 ( .C (CLK), .D (signal_7738), .Q (signal_7739) ) ;
    buf_clk cell_5611 ( .C (CLK), .D (signal_7754), .Q (signal_7755) ) ;
    buf_clk cell_5627 ( .C (CLK), .D (signal_7770), .Q (signal_7771) ) ;
    buf_clk cell_5643 ( .C (CLK), .D (signal_7786), .Q (signal_7787) ) ;
    buf_clk cell_5659 ( .C (CLK), .D (signal_7802), .Q (signal_7803) ) ;
    buf_clk cell_5675 ( .C (CLK), .D (signal_7818), .Q (signal_7819) ) ;
    buf_clk cell_5691 ( .C (CLK), .D (signal_7834), .Q (signal_7835) ) ;
    buf_clk cell_5707 ( .C (CLK), .D (signal_7850), .Q (signal_7851) ) ;
    buf_clk cell_5723 ( .C (CLK), .D (signal_7866), .Q (signal_7867) ) ;
    buf_clk cell_5739 ( .C (CLK), .D (signal_7882), .Q (signal_7883) ) ;
    buf_clk cell_5755 ( .C (CLK), .D (signal_7898), .Q (signal_7899) ) ;
    buf_clk cell_5771 ( .C (CLK), .D (signal_7914), .Q (signal_7915) ) ;
    buf_clk cell_5787 ( .C (CLK), .D (signal_7930), .Q (signal_7931) ) ;
    buf_clk cell_5803 ( .C (CLK), .D (signal_7946), .Q (signal_7947) ) ;
    buf_clk cell_5819 ( .C (CLK), .D (signal_7962), .Q (signal_7963) ) ;
    buf_clk cell_5835 ( .C (CLK), .D (signal_7978), .Q (signal_7979) ) ;
    buf_clk cell_5851 ( .C (CLK), .D (signal_7994), .Q (signal_7995) ) ;
    buf_clk cell_5867 ( .C (CLK), .D (signal_8010), .Q (signal_8011) ) ;
    buf_clk cell_5883 ( .C (CLK), .D (signal_8026), .Q (signal_8027) ) ;
    buf_clk cell_5899 ( .C (CLK), .D (signal_8042), .Q (signal_8043) ) ;
    buf_clk cell_5915 ( .C (CLK), .D (signal_8058), .Q (signal_8059) ) ;
    buf_clk cell_5931 ( .C (CLK), .D (signal_8074), .Q (signal_8075) ) ;
    buf_clk cell_5947 ( .C (CLK), .D (signal_8090), .Q (signal_8091) ) ;
    buf_clk cell_5963 ( .C (CLK), .D (signal_8106), .Q (signal_8107) ) ;
    buf_clk cell_5979 ( .C (CLK), .D (signal_8122), .Q (signal_8123) ) ;
    buf_clk cell_5995 ( .C (CLK), .D (signal_8138), .Q (signal_8139) ) ;
    buf_clk cell_6011 ( .C (CLK), .D (signal_8154), .Q (signal_8155) ) ;
    buf_clk cell_6027 ( .C (CLK), .D (signal_8170), .Q (signal_8171) ) ;
    buf_clk cell_6043 ( .C (CLK), .D (signal_8186), .Q (signal_8187) ) ;
    buf_clk cell_6059 ( .C (CLK), .D (signal_8202), .Q (signal_8203) ) ;
    buf_clk cell_6075 ( .C (CLK), .D (signal_8218), .Q (signal_8219) ) ;
    buf_clk cell_6091 ( .C (CLK), .D (signal_8234), .Q (signal_8235) ) ;
    buf_clk cell_6107 ( .C (CLK), .D (signal_8250), .Q (signal_8251) ) ;
    buf_clk cell_6123 ( .C (CLK), .D (signal_8266), .Q (signal_8267) ) ;
    buf_clk cell_6139 ( .C (CLK), .D (signal_8282), .Q (signal_8283) ) ;
    buf_clk cell_6155 ( .C (CLK), .D (signal_8298), .Q (signal_8299) ) ;
    buf_clk cell_6171 ( .C (CLK), .D (signal_8314), .Q (signal_8315) ) ;
    buf_clk cell_6187 ( .C (CLK), .D (signal_8330), .Q (signal_8331) ) ;
    buf_clk cell_6203 ( .C (CLK), .D (signal_8346), .Q (signal_8347) ) ;
    buf_clk cell_6219 ( .C (CLK), .D (signal_8362), .Q (signal_8363) ) ;
    buf_clk cell_6235 ( .C (CLK), .D (signal_8378), .Q (signal_8379) ) ;
    buf_clk cell_6251 ( .C (CLK), .D (signal_8394), .Q (signal_8395) ) ;
    buf_clk cell_6267 ( .C (CLK), .D (signal_8410), .Q (signal_8411) ) ;
    buf_clk cell_6283 ( .C (CLK), .D (signal_8426), .Q (signal_8427) ) ;
    buf_clk cell_6299 ( .C (CLK), .D (signal_8442), .Q (signal_8443) ) ;
    buf_clk cell_6315 ( .C (CLK), .D (signal_8458), .Q (signal_8459) ) ;
    buf_clk cell_6331 ( .C (CLK), .D (signal_8474), .Q (signal_8475) ) ;
    buf_clk cell_6347 ( .C (CLK), .D (signal_8490), .Q (signal_8491) ) ;
    buf_clk cell_6363 ( .C (CLK), .D (signal_8506), .Q (signal_8507) ) ;
    buf_clk cell_6379 ( .C (CLK), .D (signal_8522), .Q (signal_8523) ) ;
    buf_clk cell_6395 ( .C (CLK), .D (signal_8538), .Q (signal_8539) ) ;
    buf_clk cell_7595 ( .C (CLK), .D (signal_9738), .Q (signal_9739) ) ;
    buf_clk cell_7611 ( .C (CLK), .D (signal_9754), .Q (signal_9755) ) ;
    buf_clk cell_7627 ( .C (CLK), .D (signal_9770), .Q (signal_9771) ) ;
    buf_clk cell_7643 ( .C (CLK), .D (signal_9786), .Q (signal_9787) ) ;
    buf_clk cell_7659 ( .C (CLK), .D (signal_9802), .Q (signal_9803) ) ;
    buf_clk cell_7675 ( .C (CLK), .D (signal_9818), .Q (signal_9819) ) ;
    buf_clk cell_7691 ( .C (CLK), .D (signal_9834), .Q (signal_9835) ) ;
    buf_clk cell_7707 ( .C (CLK), .D (signal_9850), .Q (signal_9851) ) ;
    buf_clk cell_7723 ( .C (CLK), .D (signal_9866), .Q (signal_9867) ) ;
    buf_clk cell_7739 ( .C (CLK), .D (signal_9882), .Q (signal_9883) ) ;
    buf_clk cell_7947 ( .C (CLK), .D (signal_10090), .Q (signal_10091) ) ;

    /* cells in depth 7 */
    buf_clk cell_2196 ( .C (CLK), .D (signal_4339), .Q (signal_4340) ) ;
    buf_clk cell_2204 ( .C (CLK), .D (signal_4347), .Q (signal_4348) ) ;
    buf_clk cell_2212 ( .C (CLK), .D (signal_4355), .Q (signal_4356) ) ;
    buf_clk cell_2220 ( .C (CLK), .D (signal_4363), .Q (signal_4364) ) ;
    buf_clk cell_2228 ( .C (CLK), .D (signal_4371), .Q (signal_4372) ) ;
    buf_clk cell_2236 ( .C (CLK), .D (signal_4379), .Q (signal_4380) ) ;
    buf_clk cell_2244 ( .C (CLK), .D (signal_4387), .Q (signal_4388) ) ;
    buf_clk cell_2252 ( .C (CLK), .D (signal_4395), .Q (signal_4396) ) ;
    buf_clk cell_2260 ( .C (CLK), .D (signal_4403), .Q (signal_4404) ) ;
    buf_clk cell_2268 ( .C (CLK), .D (signal_4411), .Q (signal_4412) ) ;
    buf_clk cell_2272 ( .C (CLK), .D (signal_4415), .Q (signal_4416) ) ;
    buf_clk cell_2276 ( .C (CLK), .D (signal_4419), .Q (signal_4420) ) ;
    buf_clk cell_2284 ( .C (CLK), .D (signal_4427), .Q (signal_4428) ) ;
    buf_clk cell_2292 ( .C (CLK), .D (signal_4435), .Q (signal_4436) ) ;
    buf_clk cell_2296 ( .C (CLK), .D (signal_4439), .Q (signal_4440) ) ;
    buf_clk cell_2300 ( .C (CLK), .D (signal_4443), .Q (signal_4444) ) ;
    buf_clk cell_2304 ( .C (CLK), .D (signal_4447), .Q (signal_4448) ) ;
    buf_clk cell_2308 ( .C (CLK), .D (signal_4451), .Q (signal_4452) ) ;
    buf_clk cell_2316 ( .C (CLK), .D (signal_4459), .Q (signal_4460) ) ;
    buf_clk cell_2324 ( .C (CLK), .D (signal_4467), .Q (signal_4468) ) ;
    buf_clk cell_2332 ( .C (CLK), .D (signal_4475), .Q (signal_4476) ) ;
    buf_clk cell_2340 ( .C (CLK), .D (signal_4483), .Q (signal_4484) ) ;
    buf_clk cell_2344 ( .C (CLK), .D (signal_4487), .Q (signal_4488) ) ;
    buf_clk cell_2348 ( .C (CLK), .D (signal_4491), .Q (signal_4492) ) ;
    buf_clk cell_2356 ( .C (CLK), .D (signal_4499), .Q (signal_4500) ) ;
    buf_clk cell_2362 ( .C (CLK), .D (signal_4505), .Q (signal_4506) ) ;
    buf_clk cell_2368 ( .C (CLK), .D (signal_4511), .Q (signal_4512) ) ;
    buf_clk cell_2376 ( .C (CLK), .D (signal_4519), .Q (signal_4520) ) ;
    buf_clk cell_2384 ( .C (CLK), .D (signal_4527), .Q (signal_4528) ) ;
    buf_clk cell_2392 ( .C (CLK), .D (signal_4535), .Q (signal_4536) ) ;
    buf_clk cell_2400 ( .C (CLK), .D (signal_4543), .Q (signal_4544) ) ;
    buf_clk cell_2408 ( .C (CLK), .D (signal_4551), .Q (signal_4552) ) ;
    buf_clk cell_2416 ( .C (CLK), .D (signal_4559), .Q (signal_4560) ) ;
    buf_clk cell_2424 ( .C (CLK), .D (signal_4567), .Q (signal_4568) ) ;
    buf_clk cell_2432 ( .C (CLK), .D (signal_4575), .Q (signal_4576) ) ;
    buf_clk cell_2440 ( .C (CLK), .D (signal_4583), .Q (signal_4584) ) ;
    buf_clk cell_2448 ( .C (CLK), .D (signal_4591), .Q (signal_4592) ) ;
    buf_clk cell_2456 ( .C (CLK), .D (signal_4599), .Q (signal_4600) ) ;
    buf_clk cell_2464 ( .C (CLK), .D (signal_4607), .Q (signal_4608) ) ;
    buf_clk cell_2472 ( .C (CLK), .D (signal_4615), .Q (signal_4616) ) ;
    buf_clk cell_2480 ( .C (CLK), .D (signal_4623), .Q (signal_4624) ) ;
    buf_clk cell_2488 ( .C (CLK), .D (signal_4631), .Q (signal_4632) ) ;
    buf_clk cell_2496 ( .C (CLK), .D (signal_4639), .Q (signal_4640) ) ;
    buf_clk cell_2504 ( .C (CLK), .D (signal_4647), .Q (signal_4648) ) ;
    buf_clk cell_2512 ( .C (CLK), .D (signal_4655), .Q (signal_4656) ) ;
    buf_clk cell_2520 ( .C (CLK), .D (signal_4663), .Q (signal_4664) ) ;
    buf_clk cell_2528 ( .C (CLK), .D (signal_4671), .Q (signal_4672) ) ;
    buf_clk cell_2536 ( .C (CLK), .D (signal_4679), .Q (signal_4680) ) ;
    buf_clk cell_2544 ( .C (CLK), .D (signal_4687), .Q (signal_4688) ) ;
    buf_clk cell_2552 ( .C (CLK), .D (signal_4695), .Q (signal_4696) ) ;
    buf_clk cell_2560 ( .C (CLK), .D (signal_4703), .Q (signal_4704) ) ;
    buf_clk cell_2568 ( .C (CLK), .D (signal_4711), .Q (signal_4712) ) ;
    buf_clk cell_2572 ( .C (CLK), .D (signal_4715), .Q (signal_4716) ) ;
    buf_clk cell_2576 ( .C (CLK), .D (signal_4719), .Q (signal_4720) ) ;
    buf_clk cell_2580 ( .C (CLK), .D (signal_4723), .Q (signal_4724) ) ;
    buf_clk cell_2584 ( .C (CLK), .D (signal_4727), .Q (signal_4728) ) ;
    buf_clk cell_2592 ( .C (CLK), .D (signal_4735), .Q (signal_4736) ) ;
    buf_clk cell_2600 ( .C (CLK), .D (signal_4743), .Q (signal_4744) ) ;
    buf_clk cell_2608 ( .C (CLK), .D (signal_4751), .Q (signal_4752) ) ;
    buf_clk cell_2616 ( .C (CLK), .D (signal_4759), .Q (signal_4760) ) ;
    buf_clk cell_2620 ( .C (CLK), .D (signal_4763), .Q (signal_4764) ) ;
    buf_clk cell_2624 ( .C (CLK), .D (signal_4767), .Q (signal_4768) ) ;
    buf_clk cell_2630 ( .C (CLK), .D (signal_4773), .Q (signal_4774) ) ;
    buf_clk cell_2636 ( .C (CLK), .D (signal_4779), .Q (signal_4780) ) ;
    buf_clk cell_2644 ( .C (CLK), .D (signal_4787), .Q (signal_4788) ) ;
    buf_clk cell_2652 ( .C (CLK), .D (signal_4795), .Q (signal_4796) ) ;
    buf_clk cell_2660 ( .C (CLK), .D (signal_4803), .Q (signal_4804) ) ;
    buf_clk cell_2668 ( .C (CLK), .D (signal_4811), .Q (signal_4812) ) ;
    buf_clk cell_2674 ( .C (CLK), .D (signal_4817), .Q (signal_4818) ) ;
    buf_clk cell_2680 ( .C (CLK), .D (signal_4823), .Q (signal_4824) ) ;
    buf_clk cell_2684 ( .C (CLK), .D (signal_4827), .Q (signal_4828) ) ;
    buf_clk cell_2688 ( .C (CLK), .D (signal_4831), .Q (signal_4832) ) ;
    buf_clk cell_2696 ( .C (CLK), .D (signal_4839), .Q (signal_4840) ) ;
    buf_clk cell_2704 ( .C (CLK), .D (signal_4847), .Q (signal_4848) ) ;
    buf_clk cell_2712 ( .C (CLK), .D (signal_4855), .Q (signal_4856) ) ;
    buf_clk cell_2720 ( .C (CLK), .D (signal_4863), .Q (signal_4864) ) ;
    buf_clk cell_2728 ( .C (CLK), .D (signal_4871), .Q (signal_4872) ) ;
    buf_clk cell_2736 ( .C (CLK), .D (signal_4879), .Q (signal_4880) ) ;
    buf_clk cell_2744 ( .C (CLK), .D (signal_4887), .Q (signal_4888) ) ;
    buf_clk cell_2752 ( .C (CLK), .D (signal_4895), .Q (signal_4896) ) ;
    buf_clk cell_2760 ( .C (CLK), .D (signal_4903), .Q (signal_4904) ) ;
    buf_clk cell_2768 ( .C (CLK), .D (signal_4911), .Q (signal_4912) ) ;
    buf_clk cell_2776 ( .C (CLK), .D (signal_4919), .Q (signal_4920) ) ;
    buf_clk cell_2784 ( .C (CLK), .D (signal_4927), .Q (signal_4928) ) ;
    buf_clk cell_3010 ( .C (CLK), .D (signal_5119), .Q (signal_5154) ) ;
    buf_clk cell_3012 ( .C (CLK), .D (signal_5125), .Q (signal_5156) ) ;
    buf_clk cell_3018 ( .C (CLK), .D (signal_5161), .Q (signal_5162) ) ;
    buf_clk cell_3024 ( .C (CLK), .D (signal_5167), .Q (signal_5168) ) ;
    buf_clk cell_3026 ( .C (CLK), .D (signal_5015), .Q (signal_5170) ) ;
    buf_clk cell_3028 ( .C (CLK), .D (signal_5017), .Q (signal_5172) ) ;
    buf_clk cell_3030 ( .C (CLK), .D (signal_1570), .Q (signal_5174) ) ;
    buf_clk cell_3032 ( .C (CLK), .D (signal_2528), .Q (signal_5176) ) ;
    buf_clk cell_3034 ( .C (CLK), .D (signal_1572), .Q (signal_5178) ) ;
    buf_clk cell_3036 ( .C (CLK), .D (signal_2530), .Q (signal_5180) ) ;
    buf_clk cell_3038 ( .C (CLK), .D (signal_1571), .Q (signal_5182) ) ;
    buf_clk cell_3040 ( .C (CLK), .D (signal_2529), .Q (signal_5184) ) ;
    buf_clk cell_3042 ( .C (CLK), .D (signal_5043), .Q (signal_5186) ) ;
    buf_clk cell_3044 ( .C (CLK), .D (signal_5045), .Q (signal_5188) ) ;
    buf_clk cell_3046 ( .C (CLK), .D (signal_1576), .Q (signal_5190) ) ;
    buf_clk cell_3048 ( .C (CLK), .D (signal_2534), .Q (signal_5192) ) ;
    buf_clk cell_3050 ( .C (CLK), .D (signal_1581), .Q (signal_5194) ) ;
    buf_clk cell_3052 ( .C (CLK), .D (signal_2539), .Q (signal_5196) ) ;
    buf_clk cell_3060 ( .C (CLK), .D (signal_5203), .Q (signal_5204) ) ;
    buf_clk cell_3068 ( .C (CLK), .D (signal_5211), .Q (signal_5212) ) ;
    buf_clk cell_3070 ( .C (CLK), .D (signal_1616), .Q (signal_5214) ) ;
    buf_clk cell_3072 ( .C (CLK), .D (signal_2564), .Q (signal_5216) ) ;
    buf_clk cell_3074 ( .C (CLK), .D (signal_1618), .Q (signal_5218) ) ;
    buf_clk cell_3076 ( .C (CLK), .D (signal_2566), .Q (signal_5220) ) ;
    buf_clk cell_3078 ( .C (CLK), .D (signal_1617), .Q (signal_5222) ) ;
    buf_clk cell_3080 ( .C (CLK), .D (signal_2565), .Q (signal_5224) ) ;
    buf_clk cell_3082 ( .C (CLK), .D (signal_1615), .Q (signal_5226) ) ;
    buf_clk cell_3084 ( .C (CLK), .D (signal_2563), .Q (signal_5228) ) ;
    buf_clk cell_3088 ( .C (CLK), .D (signal_5231), .Q (signal_5232) ) ;
    buf_clk cell_3092 ( .C (CLK), .D (signal_5235), .Q (signal_5236) ) ;
    buf_clk cell_3094 ( .C (CLK), .D (signal_1626), .Q (signal_5238) ) ;
    buf_clk cell_3096 ( .C (CLK), .D (signal_2572), .Q (signal_5240) ) ;
    buf_clk cell_3098 ( .C (CLK), .D (signal_1627), .Q (signal_5242) ) ;
    buf_clk cell_3100 ( .C (CLK), .D (signal_2573), .Q (signal_5244) ) ;
    buf_clk cell_3102 ( .C (CLK), .D (signal_4995), .Q (signal_5246) ) ;
    buf_clk cell_3104 ( .C (CLK), .D (signal_5001), .Q (signal_5248) ) ;
    buf_clk cell_3106 ( .C (CLK), .D (signal_5129), .Q (signal_5250) ) ;
    buf_clk cell_3108 ( .C (CLK), .D (signal_5133), .Q (signal_5252) ) ;
    buf_clk cell_3110 ( .C (CLK), .D (signal_1640), .Q (signal_5254) ) ;
    buf_clk cell_3112 ( .C (CLK), .D (signal_2491), .Q (signal_5256) ) ;
    buf_clk cell_3114 ( .C (CLK), .D (signal_1641), .Q (signal_5258) ) ;
    buf_clk cell_3116 ( .C (CLK), .D (signal_2492), .Q (signal_5260) ) ;
    buf_clk cell_3118 ( .C (CLK), .D (signal_1646), .Q (signal_5262) ) ;
    buf_clk cell_3120 ( .C (CLK), .D (signal_2588), .Q (signal_5264) ) ;
    buf_clk cell_3122 ( .C (CLK), .D (signal_1647), .Q (signal_5266) ) ;
    buf_clk cell_3124 ( .C (CLK), .D (signal_2589), .Q (signal_5268) ) ;
    buf_clk cell_3126 ( .C (CLK), .D (signal_1573), .Q (signal_5270) ) ;
    buf_clk cell_3128 ( .C (CLK), .D (signal_2531), .Q (signal_5272) ) ;
    buf_clk cell_3198 ( .C (CLK), .D (signal_5341), .Q (signal_5342) ) ;
    buf_clk cell_3206 ( .C (CLK), .D (signal_5349), .Q (signal_5350) ) ;
    buf_clk cell_3230 ( .C (CLK), .D (signal_5135), .Q (signal_5374) ) ;
    buf_clk cell_3234 ( .C (CLK), .D (signal_5137), .Q (signal_5378) ) ;
    buf_clk cell_3298 ( .C (CLK), .D (signal_4959), .Q (signal_5442) ) ;
    buf_clk cell_3304 ( .C (CLK), .D (signal_4965), .Q (signal_5448) ) ;
    buf_clk cell_3320 ( .C (CLK), .D (signal_5463), .Q (signal_5464) ) ;
    buf_clk cell_3328 ( .C (CLK), .D (signal_5471), .Q (signal_5472) ) ;
    buf_clk cell_3338 ( .C (CLK), .D (signal_4947), .Q (signal_5482) ) ;
    buf_clk cell_3344 ( .C (CLK), .D (signal_4953), .Q (signal_5488) ) ;
    buf_clk cell_3356 ( .C (CLK), .D (signal_5499), .Q (signal_5500) ) ;
    buf_clk cell_3364 ( .C (CLK), .D (signal_5507), .Q (signal_5508) ) ;
    buf_clk cell_3452 ( .C (CLK), .D (signal_5595), .Q (signal_5596) ) ;
    buf_clk cell_3468 ( .C (CLK), .D (signal_5611), .Q (signal_5612) ) ;
    buf_clk cell_3492 ( .C (CLK), .D (signal_5635), .Q (signal_5636) ) ;
    buf_clk cell_3508 ( .C (CLK), .D (signal_5651), .Q (signal_5652) ) ;
    buf_clk cell_3532 ( .C (CLK), .D (signal_5675), .Q (signal_5676) ) ;
    buf_clk cell_3548 ( .C (CLK), .D (signal_5691), .Q (signal_5692) ) ;
    buf_clk cell_3564 ( .C (CLK), .D (signal_5707), .Q (signal_5708) ) ;
    buf_clk cell_3580 ( .C (CLK), .D (signal_5723), .Q (signal_5724) ) ;
    buf_clk cell_3640 ( .C (CLK), .D (signal_5783), .Q (signal_5784) ) ;
    buf_clk cell_3656 ( .C (CLK), .D (signal_5799), .Q (signal_5800) ) ;
    buf_clk cell_3672 ( .C (CLK), .D (signal_5815), .Q (signal_5816) ) ;
    buf_clk cell_3688 ( .C (CLK), .D (signal_5831), .Q (signal_5832) ) ;
    buf_clk cell_3704 ( .C (CLK), .D (signal_5847), .Q (signal_5848) ) ;
    buf_clk cell_3720 ( .C (CLK), .D (signal_5863), .Q (signal_5864) ) ;
    buf_clk cell_3736 ( .C (CLK), .D (signal_5879), .Q (signal_5880) ) ;
    buf_clk cell_3752 ( .C (CLK), .D (signal_5895), .Q (signal_5896) ) ;
    buf_clk cell_3768 ( .C (CLK), .D (signal_5911), .Q (signal_5912) ) ;
    buf_clk cell_3784 ( .C (CLK), .D (signal_5927), .Q (signal_5928) ) ;
    buf_clk cell_3892 ( .C (CLK), .D (signal_6035), .Q (signal_6036) ) ;
    buf_clk cell_3908 ( .C (CLK), .D (signal_6051), .Q (signal_6052) ) ;
    buf_clk cell_3924 ( .C (CLK), .D (signal_6067), .Q (signal_6068) ) ;
    buf_clk cell_3940 ( .C (CLK), .D (signal_6083), .Q (signal_6084) ) ;
    buf_clk cell_3956 ( .C (CLK), .D (signal_6099), .Q (signal_6100) ) ;
    buf_clk cell_3972 ( .C (CLK), .D (signal_6115), .Q (signal_6116) ) ;
    buf_clk cell_3988 ( .C (CLK), .D (signal_6131), .Q (signal_6132) ) ;
    buf_clk cell_4004 ( .C (CLK), .D (signal_6147), .Q (signal_6148) ) ;
    buf_clk cell_4020 ( .C (CLK), .D (signal_6163), .Q (signal_6164) ) ;
    buf_clk cell_4036 ( .C (CLK), .D (signal_6179), .Q (signal_6180) ) ;
    buf_clk cell_4052 ( .C (CLK), .D (signal_6195), .Q (signal_6196) ) ;
    buf_clk cell_4068 ( .C (CLK), .D (signal_6211), .Q (signal_6212) ) ;
    buf_clk cell_4084 ( .C (CLK), .D (signal_6227), .Q (signal_6228) ) ;
    buf_clk cell_4100 ( .C (CLK), .D (signal_6243), .Q (signal_6244) ) ;
    buf_clk cell_4110 ( .C (CLK), .D (signal_4983), .Q (signal_6254) ) ;
    buf_clk cell_4120 ( .C (CLK), .D (signal_4989), .Q (signal_6264) ) ;
    buf_clk cell_4158 ( .C (CLK), .D (signal_5023), .Q (signal_6302) ) ;
    buf_clk cell_4168 ( .C (CLK), .D (signal_5025), .Q (signal_6312) ) ;
    buf_clk cell_4184 ( .C (CLK), .D (signal_6327), .Q (signal_6328) ) ;
    buf_clk cell_4196 ( .C (CLK), .D (signal_6339), .Q (signal_6340) ) ;
    buf_clk cell_4208 ( .C (CLK), .D (signal_6351), .Q (signal_6352) ) ;
    buf_clk cell_4236 ( .C (CLK), .D (signal_6379), .Q (signal_6380) ) ;
    buf_clk cell_4248 ( .C (CLK), .D (signal_6391), .Q (signal_6392) ) ;
    buf_clk cell_4262 ( .C (CLK), .D (signal_6405), .Q (signal_6406) ) ;
    buf_clk cell_4276 ( .C (CLK), .D (signal_6419), .Q (signal_6420) ) ;
    buf_clk cell_4292 ( .C (CLK), .D (signal_6435), .Q (signal_6436) ) ;
    buf_clk cell_4308 ( .C (CLK), .D (signal_6451), .Q (signal_6452) ) ;
    buf_clk cell_4324 ( .C (CLK), .D (signal_6467), .Q (signal_6468) ) ;
    buf_clk cell_4340 ( .C (CLK), .D (signal_6483), .Q (signal_6484) ) ;
    buf_clk cell_4356 ( .C (CLK), .D (signal_6499), .Q (signal_6500) ) ;
    buf_clk cell_4372 ( .C (CLK), .D (signal_6515), .Q (signal_6516) ) ;
    buf_clk cell_4388 ( .C (CLK), .D (signal_6531), .Q (signal_6532) ) ;
    buf_clk cell_4404 ( .C (CLK), .D (signal_6547), .Q (signal_6548) ) ;
    buf_clk cell_4420 ( .C (CLK), .D (signal_6563), .Q (signal_6564) ) ;
    buf_clk cell_4436 ( .C (CLK), .D (signal_6579), .Q (signal_6580) ) ;
    buf_clk cell_4452 ( .C (CLK), .D (signal_6595), .Q (signal_6596) ) ;
    buf_clk cell_4468 ( .C (CLK), .D (signal_6611), .Q (signal_6612) ) ;
    buf_clk cell_4484 ( .C (CLK), .D (signal_6627), .Q (signal_6628) ) ;
    buf_clk cell_4500 ( .C (CLK), .D (signal_6643), .Q (signal_6644) ) ;
    buf_clk cell_4516 ( .C (CLK), .D (signal_6659), .Q (signal_6660) ) ;
    buf_clk cell_4532 ( .C (CLK), .D (signal_6675), .Q (signal_6676) ) ;
    buf_clk cell_4542 ( .C (CLK), .D (signal_5007), .Q (signal_6686) ) ;
    buf_clk cell_4552 ( .C (CLK), .D (signal_5013), .Q (signal_6696) ) ;
    buf_clk cell_4580 ( .C (CLK), .D (signal_6723), .Q (signal_6724) ) ;
    buf_clk cell_4592 ( .C (CLK), .D (signal_6735), .Q (signal_6736) ) ;
    buf_clk cell_4606 ( .C (CLK), .D (signal_6749), .Q (signal_6750) ) ;
    buf_clk cell_4620 ( .C (CLK), .D (signal_6763), .Q (signal_6764) ) ;
    buf_clk cell_4636 ( .C (CLK), .D (signal_6779), .Q (signal_6780) ) ;
    buf_clk cell_4652 ( .C (CLK), .D (signal_6795), .Q (signal_6796) ) ;
    buf_clk cell_4690 ( .C (CLK), .D (signal_5081), .Q (signal_6834) ) ;
    buf_clk cell_4700 ( .C (CLK), .D (signal_5085), .Q (signal_6844) ) ;
    buf_clk cell_4712 ( .C (CLK), .D (signal_6855), .Q (signal_6856) ) ;
    buf_clk cell_4724 ( .C (CLK), .D (signal_6867), .Q (signal_6868) ) ;
    buf_clk cell_4748 ( .C (CLK), .D (signal_6891), .Q (signal_6892) ) ;
    buf_clk cell_4764 ( .C (CLK), .D (signal_6907), .Q (signal_6908) ) ;
    buf_clk cell_4780 ( .C (CLK), .D (signal_6923), .Q (signal_6924) ) ;
    buf_clk cell_4796 ( .C (CLK), .D (signal_6939), .Q (signal_6940) ) ;
    buf_clk cell_4812 ( .C (CLK), .D (signal_6955), .Q (signal_6956) ) ;
    buf_clk cell_4828 ( .C (CLK), .D (signal_6971), .Q (signal_6972) ) ;
    buf_clk cell_4844 ( .C (CLK), .D (signal_6987), .Q (signal_6988) ) ;
    buf_clk cell_4860 ( .C (CLK), .D (signal_7003), .Q (signal_7004) ) ;
    buf_clk cell_4876 ( .C (CLK), .D (signal_7019), .Q (signal_7020) ) ;
    buf_clk cell_4892 ( .C (CLK), .D (signal_7035), .Q (signal_7036) ) ;
    buf_clk cell_4908 ( .C (CLK), .D (signal_7051), .Q (signal_7052) ) ;
    buf_clk cell_4924 ( .C (CLK), .D (signal_7067), .Q (signal_7068) ) ;
    buf_clk cell_4940 ( .C (CLK), .D (signal_7083), .Q (signal_7084) ) ;
    buf_clk cell_4956 ( .C (CLK), .D (signal_7099), .Q (signal_7100) ) ;
    buf_clk cell_4972 ( .C (CLK), .D (signal_7115), .Q (signal_7116) ) ;
    buf_clk cell_4988 ( .C (CLK), .D (signal_7131), .Q (signal_7132) ) ;
    buf_clk cell_5004 ( .C (CLK), .D (signal_7147), .Q (signal_7148) ) ;
    buf_clk cell_5020 ( .C (CLK), .D (signal_7163), .Q (signal_7164) ) ;
    buf_clk cell_5036 ( .C (CLK), .D (signal_7179), .Q (signal_7180) ) ;
    buf_clk cell_5052 ( .C (CLK), .D (signal_7195), .Q (signal_7196) ) ;
    buf_clk cell_5068 ( .C (CLK), .D (signal_7211), .Q (signal_7212) ) ;
    buf_clk cell_5084 ( .C (CLK), .D (signal_7227), .Q (signal_7228) ) ;
    buf_clk cell_5100 ( .C (CLK), .D (signal_7243), .Q (signal_7244) ) ;
    buf_clk cell_5116 ( .C (CLK), .D (signal_7259), .Q (signal_7260) ) ;
    buf_clk cell_5132 ( .C (CLK), .D (signal_7275), .Q (signal_7276) ) ;
    buf_clk cell_5148 ( .C (CLK), .D (signal_7291), .Q (signal_7292) ) ;
    buf_clk cell_5164 ( .C (CLK), .D (signal_7307), .Q (signal_7308) ) ;
    buf_clk cell_5180 ( .C (CLK), .D (signal_7323), .Q (signal_7324) ) ;
    buf_clk cell_5196 ( .C (CLK), .D (signal_7339), .Q (signal_7340) ) ;
    buf_clk cell_5212 ( .C (CLK), .D (signal_7355), .Q (signal_7356) ) ;
    buf_clk cell_5228 ( .C (CLK), .D (signal_7371), .Q (signal_7372) ) ;
    buf_clk cell_5244 ( .C (CLK), .D (signal_7387), .Q (signal_7388) ) ;
    buf_clk cell_5260 ( .C (CLK), .D (signal_7403), .Q (signal_7404) ) ;
    buf_clk cell_5276 ( .C (CLK), .D (signal_7419), .Q (signal_7420) ) ;
    buf_clk cell_5292 ( .C (CLK), .D (signal_7435), .Q (signal_7436) ) ;
    buf_clk cell_5308 ( .C (CLK), .D (signal_7451), .Q (signal_7452) ) ;
    buf_clk cell_5324 ( .C (CLK), .D (signal_7467), .Q (signal_7468) ) ;
    buf_clk cell_5340 ( .C (CLK), .D (signal_7483), .Q (signal_7484) ) ;
    buf_clk cell_5356 ( .C (CLK), .D (signal_7499), .Q (signal_7500) ) ;
    buf_clk cell_5372 ( .C (CLK), .D (signal_7515), .Q (signal_7516) ) ;
    buf_clk cell_5388 ( .C (CLK), .D (signal_7531), .Q (signal_7532) ) ;
    buf_clk cell_5404 ( .C (CLK), .D (signal_7547), .Q (signal_7548) ) ;
    buf_clk cell_5420 ( .C (CLK), .D (signal_7563), .Q (signal_7564) ) ;
    buf_clk cell_5436 ( .C (CLK), .D (signal_7579), .Q (signal_7580) ) ;
    buf_clk cell_5452 ( .C (CLK), .D (signal_7595), .Q (signal_7596) ) ;
    buf_clk cell_5468 ( .C (CLK), .D (signal_7611), .Q (signal_7612) ) ;
    buf_clk cell_5484 ( .C (CLK), .D (signal_7627), .Q (signal_7628) ) ;
    buf_clk cell_5500 ( .C (CLK), .D (signal_7643), .Q (signal_7644) ) ;
    buf_clk cell_5516 ( .C (CLK), .D (signal_7659), .Q (signal_7660) ) ;
    buf_clk cell_5532 ( .C (CLK), .D (signal_7675), .Q (signal_7676) ) ;
    buf_clk cell_5548 ( .C (CLK), .D (signal_7691), .Q (signal_7692) ) ;
    buf_clk cell_5564 ( .C (CLK), .D (signal_7707), .Q (signal_7708) ) ;
    buf_clk cell_5580 ( .C (CLK), .D (signal_7723), .Q (signal_7724) ) ;
    buf_clk cell_5596 ( .C (CLK), .D (signal_7739), .Q (signal_7740) ) ;
    buf_clk cell_5612 ( .C (CLK), .D (signal_7755), .Q (signal_7756) ) ;
    buf_clk cell_5628 ( .C (CLK), .D (signal_7771), .Q (signal_7772) ) ;
    buf_clk cell_5644 ( .C (CLK), .D (signal_7787), .Q (signal_7788) ) ;
    buf_clk cell_5660 ( .C (CLK), .D (signal_7803), .Q (signal_7804) ) ;
    buf_clk cell_5676 ( .C (CLK), .D (signal_7819), .Q (signal_7820) ) ;
    buf_clk cell_5692 ( .C (CLK), .D (signal_7835), .Q (signal_7836) ) ;
    buf_clk cell_5708 ( .C (CLK), .D (signal_7851), .Q (signal_7852) ) ;
    buf_clk cell_5724 ( .C (CLK), .D (signal_7867), .Q (signal_7868) ) ;
    buf_clk cell_5740 ( .C (CLK), .D (signal_7883), .Q (signal_7884) ) ;
    buf_clk cell_5756 ( .C (CLK), .D (signal_7899), .Q (signal_7900) ) ;
    buf_clk cell_5772 ( .C (CLK), .D (signal_7915), .Q (signal_7916) ) ;
    buf_clk cell_5788 ( .C (CLK), .D (signal_7931), .Q (signal_7932) ) ;
    buf_clk cell_5804 ( .C (CLK), .D (signal_7947), .Q (signal_7948) ) ;
    buf_clk cell_5820 ( .C (CLK), .D (signal_7963), .Q (signal_7964) ) ;
    buf_clk cell_5836 ( .C (CLK), .D (signal_7979), .Q (signal_7980) ) ;
    buf_clk cell_5852 ( .C (CLK), .D (signal_7995), .Q (signal_7996) ) ;
    buf_clk cell_5868 ( .C (CLK), .D (signal_8011), .Q (signal_8012) ) ;
    buf_clk cell_5884 ( .C (CLK), .D (signal_8027), .Q (signal_8028) ) ;
    buf_clk cell_5900 ( .C (CLK), .D (signal_8043), .Q (signal_8044) ) ;
    buf_clk cell_5916 ( .C (CLK), .D (signal_8059), .Q (signal_8060) ) ;
    buf_clk cell_5932 ( .C (CLK), .D (signal_8075), .Q (signal_8076) ) ;
    buf_clk cell_5948 ( .C (CLK), .D (signal_8091), .Q (signal_8092) ) ;
    buf_clk cell_5964 ( .C (CLK), .D (signal_8107), .Q (signal_8108) ) ;
    buf_clk cell_5980 ( .C (CLK), .D (signal_8123), .Q (signal_8124) ) ;
    buf_clk cell_5996 ( .C (CLK), .D (signal_8139), .Q (signal_8140) ) ;
    buf_clk cell_6012 ( .C (CLK), .D (signal_8155), .Q (signal_8156) ) ;
    buf_clk cell_6028 ( .C (CLK), .D (signal_8171), .Q (signal_8172) ) ;
    buf_clk cell_6044 ( .C (CLK), .D (signal_8187), .Q (signal_8188) ) ;
    buf_clk cell_6060 ( .C (CLK), .D (signal_8203), .Q (signal_8204) ) ;
    buf_clk cell_6076 ( .C (CLK), .D (signal_8219), .Q (signal_8220) ) ;
    buf_clk cell_6092 ( .C (CLK), .D (signal_8235), .Q (signal_8236) ) ;
    buf_clk cell_6108 ( .C (CLK), .D (signal_8251), .Q (signal_8252) ) ;
    buf_clk cell_6124 ( .C (CLK), .D (signal_8267), .Q (signal_8268) ) ;
    buf_clk cell_6140 ( .C (CLK), .D (signal_8283), .Q (signal_8284) ) ;
    buf_clk cell_6156 ( .C (CLK), .D (signal_8299), .Q (signal_8300) ) ;
    buf_clk cell_6172 ( .C (CLK), .D (signal_8315), .Q (signal_8316) ) ;
    buf_clk cell_6188 ( .C (CLK), .D (signal_8331), .Q (signal_8332) ) ;
    buf_clk cell_6204 ( .C (CLK), .D (signal_8347), .Q (signal_8348) ) ;
    buf_clk cell_6220 ( .C (CLK), .D (signal_8363), .Q (signal_8364) ) ;
    buf_clk cell_6236 ( .C (CLK), .D (signal_8379), .Q (signal_8380) ) ;
    buf_clk cell_6252 ( .C (CLK), .D (signal_8395), .Q (signal_8396) ) ;
    buf_clk cell_6268 ( .C (CLK), .D (signal_8411), .Q (signal_8412) ) ;
    buf_clk cell_6284 ( .C (CLK), .D (signal_8427), .Q (signal_8428) ) ;
    buf_clk cell_6300 ( .C (CLK), .D (signal_8443), .Q (signal_8444) ) ;
    buf_clk cell_6316 ( .C (CLK), .D (signal_8459), .Q (signal_8460) ) ;
    buf_clk cell_6332 ( .C (CLK), .D (signal_8475), .Q (signal_8476) ) ;
    buf_clk cell_6348 ( .C (CLK), .D (signal_8491), .Q (signal_8492) ) ;
    buf_clk cell_6364 ( .C (CLK), .D (signal_8507), .Q (signal_8508) ) ;
    buf_clk cell_6380 ( .C (CLK), .D (signal_8523), .Q (signal_8524) ) ;
    buf_clk cell_6396 ( .C (CLK), .D (signal_8539), .Q (signal_8540) ) ;
    buf_clk cell_7562 ( .C (CLK), .D (signal_4935), .Q (signal_9706) ) ;
    buf_clk cell_7570 ( .C (CLK), .D (signal_4941), .Q (signal_9714) ) ;
    buf_clk cell_7596 ( .C (CLK), .D (signal_9739), .Q (signal_9740) ) ;
    buf_clk cell_7612 ( .C (CLK), .D (signal_9755), .Q (signal_9756) ) ;
    buf_clk cell_7628 ( .C (CLK), .D (signal_9771), .Q (signal_9772) ) ;
    buf_clk cell_7644 ( .C (CLK), .D (signal_9787), .Q (signal_9788) ) ;
    buf_clk cell_7660 ( .C (CLK), .D (signal_9803), .Q (signal_9804) ) ;
    buf_clk cell_7676 ( .C (CLK), .D (signal_9819), .Q (signal_9820) ) ;
    buf_clk cell_7692 ( .C (CLK), .D (signal_9835), .Q (signal_9836) ) ;
    buf_clk cell_7708 ( .C (CLK), .D (signal_9851), .Q (signal_9852) ) ;
    buf_clk cell_7724 ( .C (CLK), .D (signal_9867), .Q (signal_9868) ) ;
    buf_clk cell_7740 ( .C (CLK), .D (signal_9883), .Q (signal_9884) ) ;
    buf_clk cell_7948 ( .C (CLK), .D (signal_10091), .Q (signal_10092) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_40 ( .s (signal_4341), .b ({signal_2960, signal_1326}), .a ({signal_4357, signal_4349}), .c ({signal_2984, signal_1262}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_42 ( .s (signal_4365), .b ({signal_2922, signal_1324}), .a ({signal_4381, signal_4373}), .c ({signal_2949, signal_1260}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_44 ( .s (signal_4365), .b ({signal_2965, signal_1322}), .a ({signal_4397, signal_4389}), .c ({signal_2986, signal_1258}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_46 ( .s (signal_4365), .b ({signal_2882, signal_1320}), .a ({signal_4413, signal_4405}), .c ({signal_2918, signal_1256}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_48 ( .s (signal_4365), .b ({signal_2932, signal_1318}), .a ({signal_4421, signal_4417}), .c ({signal_2951, signal_1254}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_50 ( .s (signal_4365), .b ({signal_2885, signal_1316}), .a ({signal_4437, signal_4429}), .c ({signal_2919, signal_1252}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_52 ( .s (signal_4365), .b ({signal_2935, signal_1314}), .a ({signal_4445, signal_4441}), .c ({signal_2952, signal_1250}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_54 ( .s (signal_4365), .b ({signal_2936, signal_1312}), .a ({signal_4453, signal_4449}), .c ({signal_2953, signal_1248}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_57 ( .s (signal_4341), .b ({signal_3041, signal_1309}), .a ({signal_4469, signal_4461}), .c ({signal_3059, signal_1245}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_61 ( .s (signal_4341), .b ({signal_3045, signal_1305}), .a ({signal_4485, signal_4477}), .c ({signal_3060, signal_1241}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_65 ( .s (signal_4341), .b ({signal_3010, signal_1301}), .a ({signal_4493, signal_4489}), .c ({signal_3022, signal_1237}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_69 ( .s (signal_4501), .b ({signal_3014, signal_1297}), .a ({signal_4513, signal_4507}), .c ({signal_3024, signal_1233}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_104 ( .s (signal_4521), .b ({signal_2984, signal_1262}), .a ({signal_4537, signal_4529}), .c ({signal_3028, signal_1198}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_106 ( .s (signal_4521), .b ({signal_2949, signal_1260}), .a ({signal_4553, signal_4545}), .c ({signal_2992, signal_1196}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_108 ( .s (signal_4521), .b ({signal_2986, signal_1258}), .a ({signal_4569, signal_4561}), .c ({signal_3032, signal_1194}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_110 ( .s (signal_4521), .b ({signal_2918, signal_1256}), .a ({signal_4585, signal_4577}), .c ({signal_2955, signal_1192}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_112 ( .s (signal_4521), .b ({signal_2951, signal_1254}), .a ({signal_4601, signal_4593}), .c ({signal_2996, signal_1190}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_114 ( .s (signal_4521), .b ({signal_2919, signal_1252}), .a ({signal_4617, signal_4609}), .c ({signal_2957, signal_1188}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_116 ( .s (signal_4521), .b ({signal_2952, signal_1250}), .a ({signal_4633, signal_4625}), .c ({signal_2998, signal_1186}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_118 ( .s (signal_4521), .b ({signal_2953, signal_1248}), .a ({signal_4649, signal_4641}), .c ({signal_3000, signal_1184}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_121 ( .s (signal_4521), .b ({signal_3059, signal_1245}), .a ({signal_4665, signal_4657}), .c ({signal_3112, signal_1181}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_125 ( .s (signal_4521), .b ({signal_3060, signal_1241}), .a ({signal_4681, signal_4673}), .c ({signal_3114, signal_1177}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_129 ( .s (signal_4521), .b ({signal_3022, signal_1237}), .a ({signal_4697, signal_4689}), .c ({signal_3073, signal_1173}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_133 ( .s (signal_4521), .b ({signal_3024, signal_1233}), .a ({signal_4713, signal_4705}), .c ({signal_3077, signal_1169}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_412 ( .a ({signal_4721, signal_4717}), .b ({signal_2641, signal_356}), .c ({signal_2734, signal_940}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_435 ( .a ({signal_4729, signal_4725}), .b ({signal_2642, signal_375}), .c ({signal_2735, signal_936}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_458 ( .a ({signal_4745, signal_4737}), .b ({signal_2598, signal_394}), .c ({signal_2633, signal_932}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_481 ( .a ({signal_4761, signal_4753}), .b ({signal_2599, signal_413}), .c ({signal_2634, signal_928}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_504 ( .a ({signal_4769, signal_4765}), .b ({signal_2643, signal_432}), .c ({signal_2736, signal_924}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_527 ( .a ({signal_4781, signal_4775}), .b ({signal_2644, signal_451}), .c ({signal_2737, signal_920}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_550 ( .a ({signal_4797, signal_4789}), .b ({signal_2600, signal_470}), .c ({signal_2635, signal_916}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_573 ( .a ({signal_4813, signal_4805}), .b ({signal_2601, signal_489}), .c ({signal_2636, signal_912}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_596 ( .a ({signal_4825, signal_4819}), .b ({signal_2645, signal_508}), .c ({signal_2738, signal_908}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_619 ( .a ({signal_4833, signal_4829}), .b ({signal_2646, signal_527}), .c ({signal_2739, signal_904}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_642 ( .a ({signal_4849, signal_4841}), .b ({signal_2602, signal_546}), .c ({signal_2637, signal_900}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_665 ( .a ({signal_4865, signal_4857}), .b ({signal_2603, signal_565}), .c ({signal_2638, signal_896}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_688 ( .a ({signal_4881, signal_4873}), .b ({signal_2647, signal_584}), .c ({signal_2740, signal_892}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_711 ( .a ({signal_4897, signal_4889}), .b ({signal_2648, signal_603}), .c ({signal_2741, signal_888}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_734 ( .a ({signal_4913, signal_4905}), .b ({signal_2604, signal_622}), .c ({signal_2639, signal_884}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_757 ( .a ({signal_4929, signal_4921}), .b ({signal_2605, signal_641}), .c ({signal_2640, signal_880}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_763 ( .a ({signal_2922, signal_1324}), .b ({signal_2622, signal_882}), .c ({signal_2958, signal_657}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_766 ( .a ({signal_2609, signal_881}), .b ({signal_2879, signal_660}), .c ({signal_2920, signal_658}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_771 ( .a ({signal_2640, signal_880}), .b ({signal_2960, signal_1326}), .c ({signal_3001, signal_665}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_774 ( .a ({signal_2608, signal_901}), .b ({signal_2922, signal_1324}), .c ({signal_2959, signal_668}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_780 ( .a ({signal_2640, signal_880}), .b ({signal_2606, signal_902}), .c ({signal_2742, signal_671}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_782 ( .a ({signal_3002, signal_672}), .b ({signal_2878, signal_673}), .c ({signal_3041, signal_1309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_783 ( .a ({signal_2816, signal_674}), .b ({signal_2622, signal_882}), .c ({signal_2878, signal_673}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_784 ( .a ({signal_2960, signal_1326}), .b ({signal_2712, signal_923}), .c ({signal_3002, signal_672}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_785 ( .a ({signal_2921, signal_675}), .b ({signal_2743, signal_676}), .c ({signal_2960, signal_1326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_786 ( .a ({signal_2607, signal_903}), .b ({signal_2637, signal_900}), .c ({signal_2743, signal_676}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_787 ( .a ({signal_2746, signal_677}), .b ({signal_2879, signal_660}), .c ({signal_2921, signal_675}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_788 ( .a ({signal_2815, signal_678}), .b ({signal_2688, signal_941}), .c ({signal_2879, signal_660}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_789 ( .a ({signal_2653, signal_922}), .b ({signal_2734, signal_940}), .c ({signal_2815, signal_678}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_793 ( .a ({signal_2608, signal_901}), .b ({signal_2637, signal_900}), .c ({signal_2744, signal_681}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_796 ( .a ({signal_2922, signal_1324}), .b ({signal_2640, signal_880}), .c ({signal_2961, signal_684}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_799 ( .a ({signal_2609, signal_881}), .b ({signal_2637, signal_900}), .c ({signal_2745, signal_686}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_809 ( .a ({signal_2640, signal_880}), .b ({signal_2610, signal_883}), .c ({signal_2746, signal_677}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_811 ( .a ({signal_2640, signal_880}), .b ({signal_2637, signal_900}), .c ({signal_2747, signal_692}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_813 ( .a ({signal_2880, signal_693}), .b ({signal_2609, signal_881}), .c ({signal_2922, signal_1324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_814 ( .a ({signal_2816, signal_674}), .b ({signal_2695, signal_942}), .c ({signal_2880, signal_693}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_815 ( .a ({signal_2608, signal_901}), .b ({signal_2737, signal_920}), .c ({signal_2816, signal_674}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_817 ( .a ({signal_2882, signal_1320}), .b ({signal_2671, signal_894}), .c ({signal_2923, signal_695}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_820 ( .a ({signal_2649, signal_893}), .b ({signal_2881, signal_698}), .c ({signal_2924, signal_696}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_825 ( .a ({signal_2740, signal_892}), .b ({signal_2965, signal_1322}), .c ({signal_3006, signal_703}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_828 ( .a ({signal_2612, signal_897}), .b ({signal_2882, signal_1320}), .c ({signal_2925, signal_706}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_834 ( .a ({signal_2740, signal_892}), .b ({signal_2613, signal_898}), .c ({signal_2817, signal_709}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_836 ( .a ({signal_3007, signal_710}), .b ({signal_2818, signal_711}), .c ({signal_3045, signal_1305}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_837 ( .a ({signal_2751, signal_712}), .b ({signal_2671, signal_894}), .c ({signal_2818, signal_711}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_838 ( .a ({signal_2965, signal_1322}), .b ({signal_2632, signal_919}), .c ({signal_3007, signal_710}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_839 ( .a ({signal_2926, signal_713}), .b ({signal_2748, signal_714}), .c ({signal_2965, signal_1322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_840 ( .a ({signal_2611, signal_899}), .b ({signal_2638, signal_896}), .c ({signal_2748, signal_714}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_841 ( .a ({signal_2820, signal_715}), .b ({signal_2881, signal_698}), .c ({signal_2926, signal_713}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_842 ( .a ({signal_2819, signal_716}), .b ({signal_2696, signal_937}), .c ({signal_2881, signal_698}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_843 ( .a ({signal_2617, signal_918}), .b ({signal_2735, signal_936}), .c ({signal_2819, signal_716}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_847 ( .a ({signal_2612, signal_897}), .b ({signal_2638, signal_896}), .c ({signal_2749, signal_719}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_850 ( .a ({signal_2882, signal_1320}), .b ({signal_2740, signal_892}), .c ({signal_2927, signal_722}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_853 ( .a ({signal_2649, signal_893}), .b ({signal_2638, signal_896}), .c ({signal_2750, signal_724}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_863 ( .a ({signal_2740, signal_892}), .b ({signal_2672, signal_895}), .c ({signal_2820, signal_715}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_865 ( .a ({signal_2740, signal_892}), .b ({signal_2638, signal_896}), .c ({signal_2821, signal_730}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_867 ( .a ({signal_2822, signal_731}), .b ({signal_2649, signal_893}), .c ({signal_2882, signal_1320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_868 ( .a ({signal_2751, signal_712}), .b ({signal_2673, signal_938}), .c ({signal_2822, signal_731}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_869 ( .a ({signal_2612, signal_897}), .b ({signal_2635, signal_916}), .c ({signal_2751, signal_712}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_871 ( .a ({signal_2885, signal_1316}), .b ({signal_2675, signal_890}), .c ({signal_2930, signal_733}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_874 ( .a ({signal_2677, signal_889}), .b ({signal_2826, signal_736}), .c ({signal_2883, signal_734}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_879 ( .a ({signal_2741, signal_888}), .b ({signal_2932, signal_1318}), .c ({signal_2969, signal_741}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_882 ( .a ({signal_2650, signal_909}), .b ({signal_2885, signal_1316}), .c ({signal_2931, signal_744}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_888 ( .a ({signal_2741, signal_888}), .b ({signal_2674, signal_910}), .c ({signal_2823, signal_747}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_890 ( .a ({signal_2970, signal_748}), .b ({signal_2824, signal_749}), .c ({signal_3010, signal_1301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_891 ( .a ({signal_2753, signal_750}), .b ({signal_2675, signal_890}), .c ({signal_2824, signal_749}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_892 ( .a ({signal_2932, signal_1318}), .b ({signal_2631, signal_915}), .c ({signal_2970, signal_748}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_893 ( .a ({signal_2884, signal_751}), .b ({signal_2825, signal_752}), .c ({signal_2932, signal_1318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_894 ( .a ({signal_2676, signal_911}), .b ({signal_2738, signal_908}), .c ({signal_2825, signal_752}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_895 ( .a ({signal_2829, signal_753}), .b ({signal_2826, signal_736}), .c ({signal_2884, signal_751}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_896 ( .a ({signal_2752, signal_754}), .b ({signal_2618, signal_933}), .c ({signal_2826, signal_736}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_897 ( .a ({signal_2615, signal_914}), .b ({signal_2633, signal_932}), .c ({signal_2752, signal_754}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_901 ( .a ({signal_2650, signal_909}), .b ({signal_2738, signal_908}), .c ({signal_2827, signal_757}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_904 ( .a ({signal_2885, signal_1316}), .b ({signal_2741, signal_888}), .c ({signal_2933, signal_760}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_907 ( .a ({signal_2677, signal_889}), .b ({signal_2738, signal_908}), .c ({signal_2828, signal_762}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_917 ( .a ({signal_2741, signal_888}), .b ({signal_2679, signal_891}), .c ({signal_2829, signal_753}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_919 ( .a ({signal_2741, signal_888}), .b ({signal_2738, signal_908}), .c ({signal_2830, signal_768}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_921 ( .a ({signal_2831, signal_769}), .b ({signal_2677, signal_889}), .c ({signal_2885, signal_1316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_922 ( .a ({signal_2753, signal_750}), .b ({signal_2619, signal_934}), .c ({signal_2831, signal_769}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_923 ( .a ({signal_2650, signal_909}), .b ({signal_2636, signal_912}), .c ({signal_2753, signal_750}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_925 ( .a ({signal_2936, signal_1312}), .b ({signal_2627, signal_886}), .c ({signal_2975, signal_771}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_928 ( .a ({signal_2621, signal_885}), .b ({signal_2833, signal_774}), .c ({signal_2886, signal_772}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_933 ( .a ({signal_2639, signal_884}), .b ({signal_2935, signal_1314}), .c ({signal_2976, signal_779}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_936 ( .a ({signal_2681, signal_905}), .b ({signal_2936, signal_1312}), .c ({signal_2977, signal_782}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_942 ( .a ({signal_2639, signal_884}), .b ({signal_2651, signal_906}), .c ({signal_2754, signal_785}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_944 ( .a ({signal_2978, signal_786}), .b ({signal_2887, signal_787}), .c ({signal_3014, signal_1297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_945 ( .a ({signal_2837, signal_788}), .b ({signal_2627, signal_886}), .c ({signal_2887, signal_787}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_946 ( .a ({signal_2935, signal_1314}), .b ({signal_2711, signal_927}), .c ({signal_2978, signal_786}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_947 ( .a ({signal_2888, signal_789}), .b ({signal_2832, signal_790}), .c ({signal_2935, signal_1314}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_948 ( .a ({signal_2680, signal_907}), .b ({signal_2739, signal_904}), .c ({signal_2832, signal_790}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_949 ( .a ({signal_2756, signal_791}), .b ({signal_2833, signal_774}), .c ({signal_2888, signal_789}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_950 ( .a ({signal_2755, signal_792}), .b ({signal_2620, signal_929}), .c ({signal_2833, signal_774}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_951 ( .a ({signal_2652, signal_926}), .b ({signal_2634, signal_928}), .c ({signal_2755, signal_792}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_955 ( .a ({signal_2681, signal_905}), .b ({signal_2739, signal_904}), .c ({signal_2834, signal_795}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_958 ( .a ({signal_2936, signal_1312}), .b ({signal_2639, signal_884}), .c ({signal_2979, signal_798}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_961 ( .a ({signal_2621, signal_885}), .b ({signal_2739, signal_904}), .c ({signal_2835, signal_800}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_971 ( .a ({signal_2639, signal_884}), .b ({signal_2616, signal_887}), .c ({signal_2756, signal_791}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_973 ( .a ({signal_2639, signal_884}), .b ({signal_2739, signal_904}), .c ({signal_2836, signal_806}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_975 ( .a ({signal_2889, signal_807}), .b ({signal_2621, signal_885}), .c ({signal_2936, signal_1312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_976 ( .a ({signal_2837, signal_788}), .b ({signal_2629, signal_930}), .c ({signal_2889, signal_807}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_977 ( .a ({signal_2681, signal_905}), .b ({signal_2736, signal_924}), .c ({signal_2837, signal_788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1460 ( .s ({signal_4743, signal_4735}), .b ({signal_2444, signal_1506}), .a ({signal_2443, signal_1505}), .clk (CLK), .r (Fresh[332]), .c ({signal_2598, signal_394}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1461 ( .s ({signal_4759, signal_4751}), .b ({signal_2446, signal_1508}), .a ({signal_2445, signal_1507}), .clk (CLK), .r (Fresh[333]), .c ({signal_2599, signal_413}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1462 ( .s ({signal_4795, signal_4787}), .b ({signal_2448, signal_1510}), .a ({signal_2447, signal_1509}), .clk (CLK), .r (Fresh[334]), .c ({signal_2600, signal_470}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1463 ( .s ({signal_4811, signal_4803}), .b ({signal_2450, signal_1512}), .a ({signal_2449, signal_1511}), .clk (CLK), .r (Fresh[335]), .c ({signal_2601, signal_489}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1464 ( .s ({signal_4847, signal_4839}), .b ({signal_2452, signal_1514}), .a ({signal_2451, signal_1513}), .clk (CLK), .r (Fresh[336]), .c ({signal_2602, signal_546}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1465 ( .s ({signal_4863, signal_4855}), .b ({signal_2454, signal_1516}), .a ({signal_2453, signal_1515}), .clk (CLK), .r (Fresh[337]), .c ({signal_2603, signal_565}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1466 ( .s ({signal_4911, signal_4903}), .b ({signal_2456, signal_1518}), .a ({signal_2455, signal_1517}), .clk (CLK), .r (Fresh[338]), .c ({signal_2604, signal_622}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1467 ( .s ({signal_4927, signal_4919}), .b ({signal_2458, signal_1520}), .a ({signal_2457, signal_1519}), .clk (CLK), .r (Fresh[339]), .c ({signal_2605, signal_641}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1468 ( .s ({signal_4941, signal_4935}), .b ({signal_2500, signal_1522}), .a ({signal_2499, signal_1521}), .clk (CLK), .r (Fresh[340]), .c ({signal_2641, signal_356}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1469 ( .s ({signal_4411, signal_4403}), .b ({signal_2502, signal_1524}), .a ({signal_2501, signal_1523}), .clk (CLK), .r (Fresh[341]), .c ({signal_2642, signal_375}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1470 ( .s ({signal_4953, signal_4947}), .b ({signal_2504, signal_1526}), .a ({signal_2503, signal_1525}), .clk (CLK), .r (Fresh[342]), .c ({signal_2643, signal_432}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1471 ( .s ({signal_4965, signal_4959}), .b ({signal_2506, signal_1528}), .a ({signal_2505, signal_1527}), .clk (CLK), .r (Fresh[343]), .c ({signal_2644, signal_451}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1472 ( .s ({signal_4977, signal_4971}), .b ({signal_2508, signal_1530}), .a ({signal_2507, signal_1529}), .clk (CLK), .r (Fresh[344]), .c ({signal_2645, signal_508}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1473 ( .s ({signal_4989, signal_4983}), .b ({signal_2510, signal_1532}), .a ({signal_2509, signal_1531}), .clk (CLK), .r (Fresh[345]), .c ({signal_2646, signal_527}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1474 ( .s ({signal_5001, signal_4995}), .b ({signal_2512, signal_1534}), .a ({signal_2511, signal_1533}), .clk (CLK), .r (Fresh[346]), .c ({signal_2647, signal_584}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1475 ( .s ({signal_5013, signal_5007}), .b ({signal_2514, signal_1536}), .a ({signal_2513, signal_1535}), .clk (CLK), .r (Fresh[347]), .c ({signal_2648, signal_603}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1476 ( .s ({signal_4847, signal_4839}), .b ({signal_2460, signal_1538}), .a ({signal_2459, signal_1537}), .clk (CLK), .r (Fresh[348]), .c ({signal_2606, signal_902}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1477 ( .s ({signal_4847, signal_4839}), .b ({signal_2462, signal_1540}), .a ({signal_2461, signal_1539}), .clk (CLK), .r (Fresh[349]), .c ({signal_2607, signal_903}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1478 ( .s ({signal_4847, signal_4839}), .b ({signal_2464, signal_1542}), .a ({signal_2463, signal_1541}), .clk (CLK), .r (Fresh[350]), .c ({signal_2608, signal_901}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1479 ( .s ({signal_4927, signal_4919}), .b ({signal_2466, signal_1544}), .a ({signal_2465, signal_1543}), .clk (CLK), .r (Fresh[351]), .c ({signal_2609, signal_881}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1480 ( .s ({signal_4927, signal_4919}), .b ({signal_2468, signal_1546}), .a ({signal_2467, signal_1545}), .clk (CLK), .r (Fresh[352]), .c ({signal_2610, signal_883}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1481 ( .s ({signal_4863, signal_4855}), .b ({signal_2470, signal_1548}), .a ({signal_2469, signal_1547}), .clk (CLK), .r (Fresh[353]), .c ({signal_2611, signal_899}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1482 ( .s ({signal_4863, signal_4855}), .b ({signal_2472, signal_1550}), .a ({signal_2471, signal_1549}), .clk (CLK), .r (Fresh[354]), .c ({signal_2612, signal_897}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1483 ( .s ({signal_5001, signal_4995}), .b ({signal_2516, signal_1552}), .a ({signal_2515, signal_1551}), .clk (CLK), .r (Fresh[355]), .c ({signal_2649, signal_893}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1484 ( .s ({signal_4863, signal_4855}), .b ({signal_2474, signal_1554}), .a ({signal_2473, signal_1553}), .clk (CLK), .r (Fresh[356]), .c ({signal_2613, signal_898}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1485 ( .s ({signal_4863, signal_4855}), .b ({signal_2453, signal_1515}), .a ({signal_2454, signal_1516}), .clk (CLK), .r (Fresh[357]), .c ({signal_2614, signal_1660}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1486 ( .s ({signal_4811, signal_4803}), .b ({signal_2476, signal_1556}), .a ({signal_2475, signal_1555}), .clk (CLK), .r (Fresh[358]), .c ({signal_2615, signal_914}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1487 ( .s ({signal_4977, signal_4971}), .b ({signal_2518, signal_1558}), .a ({signal_2517, signal_1557}), .clk (CLK), .r (Fresh[359]), .c ({signal_2650, signal_909}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1488 ( .s ({signal_4989, signal_4983}), .b ({signal_2520, signal_1560}), .a ({signal_2519, signal_1559}), .clk (CLK), .r (Fresh[360]), .c ({signal_2651, signal_906}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1489 ( .s ({signal_4953, signal_4947}), .b ({signal_2522, signal_1562}), .a ({signal_2521, signal_1561}), .clk (CLK), .r (Fresh[361]), .c ({signal_2652, signal_926}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1490 ( .s ({signal_4911, signal_4903}), .b ({signal_2478, signal_1564}), .a ({signal_2477, signal_1563}), .clk (CLK), .r (Fresh[362]), .c ({signal_2616, signal_887}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1491 ( .s ({signal_4965, signal_4959}), .b ({signal_2524, signal_1566}), .a ({signal_2523, signal_1565}), .clk (CLK), .r (Fresh[363]), .c ({signal_2653, signal_922}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1492 ( .s ({signal_5017, signal_5015}), .b ({signal_5021, signal_5019}), .a ({signal_2525, signal_1567}), .clk (CLK), .r (Fresh[364]), .c ({signal_2654, signal_1661}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1493 ( .s ({signal_5017, signal_5015}), .b ({signal_2527, signal_1569}), .a ({signal_2526, signal_1568}), .clk (CLK), .r (Fresh[365]), .c ({signal_2655, signal_1662}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1494 ( .s ({signal_5025, signal_5023}), .b ({signal_2529, signal_1571}), .a ({signal_2528, signal_1570}), .clk (CLK), .r (Fresh[366]), .c ({signal_2656, signal_1663}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1495 ( .s ({signal_5025, signal_5023}), .b ({signal_5029, signal_5027}), .a ({signal_2529, signal_1571}), .clk (CLK), .r (Fresh[367]), .c ({signal_2657, signal_1664}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1496 ( .s ({signal_5025, signal_5023}), .b ({signal_2528, signal_1570}), .a ({signal_5033, signal_5031}), .clk (CLK), .r (Fresh[368]), .c ({signal_2658, signal_1665}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1497 ( .s ({signal_5025, signal_5023}), .b ({signal_2531, signal_1573}), .a ({signal_2530, signal_1572}), .clk (CLK), .r (Fresh[369]), .c ({signal_2659, signal_1666}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1498 ( .s ({signal_5025, signal_5023}), .b ({signal_5037, signal_5035}), .a ({signal_2531, signal_1573}), .clk (CLK), .r (Fresh[370]), .c ({signal_2660, signal_1667}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1499 ( .s ({signal_5025, signal_5023}), .b ({signal_2530, signal_1572}), .a ({signal_5041, signal_5039}), .clk (CLK), .r (Fresh[371]), .c ({signal_2661, signal_1668}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1500 ( .s ({signal_5025, signal_5023}), .b ({signal_2528, signal_1570}), .a ({signal_2529, signal_1571}), .clk (CLK), .r (Fresh[372]), .c ({signal_2662, signal_1669}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1501 ( .s ({signal_5025, signal_5023}), .b ({signal_5033, signal_5031}), .a ({signal_2528, signal_1570}), .clk (CLK), .r (Fresh[373]), .c ({signal_2663, signal_1670}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1502 ( .s ({signal_5025, signal_5023}), .b ({signal_2529, signal_1571}), .a ({signal_5029, signal_5027}), .clk (CLK), .r (Fresh[374]), .c ({signal_2664, signal_1671}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1503 ( .s ({signal_5045, signal_5043}), .b ({signal_2533, signal_1575}), .a ({signal_2532, signal_1574}), .clk (CLK), .r (Fresh[375]), .c ({signal_2665, signal_1672}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1504 ( .s ({signal_5049, signal_5047}), .b ({signal_2533, signal_1575}), .a ({signal_2532, signal_1574}), .clk (CLK), .r (Fresh[376]), .c ({signal_2666, signal_1673}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1505 ( .s ({signal_5049, signal_5047}), .b ({signal_2532, signal_1574}), .a ({signal_2533, signal_1575}), .clk (CLK), .r (Fresh[377]), .c ({signal_2667, signal_1674}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1506 ( .s ({signal_5045, signal_5043}), .b ({signal_2536, signal_1578}), .a ({signal_2535, signal_1577}), .clk (CLK), .r (Fresh[378]), .c ({signal_2668, signal_1675}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1507 ( .s ({signal_5045, signal_5043}), .b ({signal_2538, signal_1580}), .a ({signal_2537, signal_1579}), .clk (CLK), .r (Fresh[379]), .c ({signal_2669, signal_1676}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1508 ( .s ({signal_5045, signal_5043}), .b ({signal_2535, signal_1577}), .a ({signal_2536, signal_1578}), .clk (CLK), .r (Fresh[380]), .c ({signal_2670, signal_1677}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1509 ( .s ({signal_5001, signal_4995}), .b ({signal_2541, signal_1583}), .a ({signal_2540, signal_1582}), .clk (CLK), .r (Fresh[381]), .c ({signal_2671, signal_894}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1510 ( .s ({signal_4795, signal_4787}), .b ({signal_2480, signal_1585}), .a ({signal_2479, signal_1584}), .clk (CLK), .r (Fresh[382]), .c ({signal_2617, signal_918}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1511 ( .s ({signal_5001, signal_4995}), .b ({signal_2543, signal_1587}), .a ({signal_2542, signal_1586}), .clk (CLK), .r (Fresh[383]), .c ({signal_2672, signal_895}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1512 ( .s ({signal_4411, signal_4403}), .b ({signal_2545, signal_1589}), .a ({signal_2544, signal_1588}), .clk (CLK), .r (Fresh[384]), .c ({signal_2673, signal_938}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1513 ( .s ({signal_4977, signal_4971}), .b ({signal_2547, signal_1591}), .a ({signal_2546, signal_1590}), .clk (CLK), .r (Fresh[385]), .c ({signal_2674, signal_910}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1514 ( .s ({signal_5013, signal_5007}), .b ({signal_2549, signal_1593}), .a ({signal_2548, signal_1592}), .clk (CLK), .r (Fresh[386]), .c ({signal_2675, signal_890}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1515 ( .s ({signal_4977, signal_4971}), .b ({signal_2551, signal_1595}), .a ({signal_2550, signal_1594}), .clk (CLK), .r (Fresh[387]), .c ({signal_2676, signal_911}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1516 ( .s ({signal_4743, signal_4735}), .b ({signal_2482, signal_1597}), .a ({signal_2481, signal_1596}), .clk (CLK), .r (Fresh[388]), .c ({signal_2618, signal_933}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1517 ( .s ({signal_5013, signal_5007}), .b ({signal_2553, signal_1599}), .a ({signal_2552, signal_1598}), .clk (CLK), .r (Fresh[389]), .c ({signal_2677, signal_889}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1518 ( .s ({signal_4977, signal_4971}), .b ({signal_2555, signal_1601}), .a ({signal_2554, signal_1600}), .clk (CLK), .r (Fresh[390]), .c ({signal_2678, signal_1678}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1519 ( .s ({signal_5013, signal_5007}), .b ({signal_2557, signal_1603}), .a ({signal_2556, signal_1602}), .clk (CLK), .r (Fresh[391]), .c ({signal_2679, signal_891}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1520 ( .s ({signal_4743, signal_4735}), .b ({signal_2484, signal_1605}), .a ({signal_2483, signal_1604}), .clk (CLK), .r (Fresh[392]), .c ({signal_2619, signal_934}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1521 ( .s ({signal_4989, signal_4983}), .b ({signal_2559, signal_1607}), .a ({signal_2558, signal_1606}), .clk (CLK), .r (Fresh[393]), .c ({signal_2680, signal_907}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1522 ( .s ({signal_4759, signal_4751}), .b ({signal_2486, signal_1609}), .a ({signal_2485, signal_1608}), .clk (CLK), .r (Fresh[394]), .c ({signal_2620, signal_929}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1523 ( .s ({signal_4989, signal_4983}), .b ({signal_2561, signal_1611}), .a ({signal_2560, signal_1610}), .clk (CLK), .r (Fresh[395]), .c ({signal_2681, signal_905}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1524 ( .s ({signal_4911, signal_4903}), .b ({signal_2488, signal_1613}), .a ({signal_2487, signal_1612}), .clk (CLK), .r (Fresh[396]), .c ({signal_2621, signal_885}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1525 ( .s ({signal_4831, signal_4827}), .b ({signal_5053, signal_5051}), .a ({signal_2562, signal_1614}), .clk (CLK), .r (Fresh[397]), .c ({signal_2682, signal_1679}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1526 ( .s ({signal_5057, signal_5055}), .b ({signal_2563, signal_1615}), .a ({signal_5061, signal_5059}), .clk (CLK), .r (Fresh[398]), .c ({signal_2683, signal_1680}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1527 ( .s ({signal_5057, signal_5055}), .b ({signal_2565, signal_1617}), .a ({signal_5065, signal_5063}), .clk (CLK), .r (Fresh[399]), .c ({signal_2684, signal_1681}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1528 ( .s ({signal_4831, signal_4827}), .b ({signal_5069, signal_5067}), .a ({signal_2567, signal_1619}), .clk (CLK), .r (Fresh[400]), .c ({signal_2685, signal_1682}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1529 ( .s ({signal_4831, signal_4827}), .b ({signal_5073, signal_5071}), .a ({signal_2568, signal_1620}), .clk (CLK), .r (Fresh[401]), .c ({signal_2686, signal_1683}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1530 ( .s ({signal_4831, signal_4827}), .b ({signal_5077, signal_5075}), .a ({signal_2569, signal_1621}), .clk (CLK), .r (Fresh[402]), .c ({signal_2687, signal_1684}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1531 ( .s ({signal_4927, signal_4919}), .b ({signal_2490, signal_1623}), .a ({signal_2489, signal_1622}), .clk (CLK), .r (Fresh[403]), .c ({signal_2622, signal_882}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1532 ( .s ({signal_4941, signal_4935}), .b ({signal_2571, signal_1625}), .a ({signal_2570, signal_1624}), .clk (CLK), .r (Fresh[404]), .c ({signal_2688, signal_941}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1533 ( .s ({signal_5085, signal_5081}), .b ({signal_2573, signal_1627}), .a ({signal_2572, signal_1626}), .clk (CLK), .r (Fresh[405]), .c ({signal_2689, signal_1685}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1534 ( .s ({signal_5085, signal_5081}), .b ({signal_5089, signal_5087}), .a ({signal_2573, signal_1627}), .clk (CLK), .r (Fresh[406]), .c ({signal_2690, signal_1686}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1535 ( .s ({signal_5085, signal_5081}), .b ({signal_2572, signal_1626}), .a ({signal_5093, signal_5091}), .clk (CLK), .r (Fresh[407]), .c ({signal_2691, signal_1687}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1536 ( .s ({signal_5085, signal_5081}), .b ({signal_2572, signal_1626}), .a ({signal_2573, signal_1627}), .clk (CLK), .r (Fresh[408]), .c ({signal_2692, signal_1688}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1537 ( .s ({signal_5085, signal_5081}), .b ({signal_5093, signal_5091}), .a ({signal_2572, signal_1626}), .clk (CLK), .r (Fresh[409]), .c ({signal_2693, signal_1689}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1538 ( .s ({signal_5085, signal_5081}), .b ({signal_2573, signal_1627}), .a ({signal_5089, signal_5087}), .clk (CLK), .r (Fresh[410]), .c ({signal_2694, signal_1690}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1539 ( .s ({signal_4941, signal_4935}), .b ({signal_2575, signal_1629}), .a ({signal_2574, signal_1628}), .clk (CLK), .r (Fresh[411]), .c ({signal_2695, signal_942}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1540 ( .s ({signal_4411, signal_4403}), .b ({signal_2577, signal_1631}), .a ({signal_2576, signal_1630}), .clk (CLK), .r (Fresh[412]), .c ({signal_2696, signal_937}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1541 ( .s ({signal_5097, signal_5095}), .b ({signal_2578, signal_1632}), .a ({signal_5101, signal_5099}), .clk (CLK), .r (Fresh[413]), .c ({signal_2697, signal_1691}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1542 ( .s ({signal_5097, signal_5095}), .b ({signal_5105, signal_5103}), .a ({signal_2579, signal_1633}), .clk (CLK), .r (Fresh[414]), .c ({signal_2698, signal_1692}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1543 ( .s ({signal_5097, signal_5095}), .b ({signal_2580, signal_1634}), .a ({signal_5109, signal_5107}), .clk (CLK), .r (Fresh[415]), .c ({signal_2699, signal_1693}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1544 ( .s ({signal_5097, signal_5095}), .b ({signal_5113, signal_5111}), .a ({signal_2581, signal_1635}), .clk (CLK), .r (Fresh[416]), .c ({signal_2700, signal_1694}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1545 ( .s ({signal_5125, signal_5119}), .b ({signal_2582, signal_1636}), .a ({signal_2576, signal_1630}), .clk (CLK), .r (Fresh[417]), .c ({signal_2701, signal_1695}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1546 ( .s ({signal_5125, signal_5119}), .b ({signal_2576, signal_1630}), .a ({signal_2582, signal_1636}), .clk (CLK), .r (Fresh[418]), .c ({signal_2702, signal_1696}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1547 ( .s ({signal_5125, signal_5119}), .b ({signal_2583, signal_1637}), .a ({signal_2577, signal_1631}), .clk (CLK), .r (Fresh[419]), .c ({signal_2703, signal_1697}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1548 ( .s ({signal_5125, signal_5119}), .b ({signal_2577, signal_1631}), .a ({signal_2583, signal_1637}), .clk (CLK), .r (Fresh[420]), .c ({signal_2704, signal_1698}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1549 ( .s ({signal_5013, signal_5007}), .b ({signal_2585, signal_1639}), .a ({signal_2584, signal_1638}), .clk (CLK), .r (Fresh[421]), .c ({signal_2705, signal_1699}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1550 ( .s ({signal_4435, signal_4427}), .b ({signal_2492, signal_1641}), .a ({signal_2491, signal_1640}), .clk (CLK), .r (Fresh[422]), .c ({signal_2623, signal_1700}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1551 ( .s ({signal_4435, signal_4427}), .b ({signal_2491, signal_1640}), .a ({signal_2492, signal_1641}), .clk (CLK), .r (Fresh[423]), .c ({signal_2624, signal_1701}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1552 ( .s ({signal_5133, signal_5129}), .b ({signal_2492, signal_1641}), .a ({signal_2491, signal_1640}), .clk (CLK), .r (Fresh[424]), .c ({signal_2625, signal_1702}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1553 ( .s ({signal_5133, signal_5129}), .b ({signal_2491, signal_1640}), .a ({signal_2492, signal_1641}), .clk (CLK), .r (Fresh[425]), .c ({signal_2626, signal_1703}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1554 ( .s ({signal_4911, signal_4903}), .b ({signal_2494, signal_1643}), .a ({signal_2493, signal_1642}), .clk (CLK), .r (Fresh[426]), .c ({signal_2627, signal_886}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1555 ( .s ({signal_4911, signal_4903}), .b ({signal_2455, signal_1517}), .a ({signal_2456, signal_1518}), .clk (CLK), .r (Fresh[427]), .c ({signal_2628, signal_1704}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1556 ( .s ({signal_5137, signal_5135}), .b ({signal_5141, signal_5139}), .a ({signal_2586, signal_1644}), .clk (CLK), .r (Fresh[428]), .c ({signal_2706, signal_1705}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1557 ( .s ({signal_5137, signal_5135}), .b ({signal_5145, signal_5143}), .a ({signal_2587, signal_1645}), .clk (CLK), .r (Fresh[429]), .c ({signal_2707, signal_1706}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1558 ( .s ({signal_5137, signal_5135}), .b ({signal_2586, signal_1644}), .a ({signal_2587, signal_1645}), .clk (CLK), .r (Fresh[430]), .c ({signal_2708, signal_1707}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1559 ( .s ({signal_5137, signal_5135}), .b ({signal_2587, signal_1645}), .a ({signal_2586, signal_1644}), .clk (CLK), .r (Fresh[431]), .c ({signal_2709, signal_1708}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1560 ( .s ({signal_4759, signal_4751}), .b ({signal_2496, signal_1649}), .a ({signal_2495, signal_1648}), .clk (CLK), .r (Fresh[432]), .c ({signal_2629, signal_930}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1561 ( .s ({signal_4863, signal_4855}), .b ({signal_2469, signal_1547}), .a ({signal_2470, signal_1548}), .clk (CLK), .r (Fresh[433]), .c ({signal_2630, signal_1709}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1562 ( .s ({signal_4811, signal_4803}), .b ({signal_2492, signal_1641}), .a ({signal_2491, signal_1640}), .clk (CLK), .r (Fresh[434]), .c ({signal_2631, signal_915}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1563 ( .s ({signal_4977, signal_4971}), .b ({signal_2550, signal_1594}), .a ({signal_2551, signal_1595}), .clk (CLK), .r (Fresh[435]), .c ({signal_2710, signal_1710}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1564 ( .s ({signal_4953, signal_4947}), .b ({signal_2591, signal_1651}), .a ({signal_2590, signal_1650}), .clk (CLK), .r (Fresh[436]), .c ({signal_2711, signal_927}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1565 ( .s ({signal_4965, signal_4959}), .b ({signal_5149, signal_5147}), .a ({signal_2592, signal_1652}), .clk (CLK), .r (Fresh[437]), .c ({signal_2712, signal_923}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1566 ( .s ({signal_5017, signal_5015}), .b ({signal_2525, signal_1567}), .a ({signal_5153, signal_5151}), .clk (CLK), .r (Fresh[438]), .c ({signal_2713, signal_1711}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1567 ( .s ({signal_5017, signal_5015}), .b ({signal_2593, signal_1653}), .a ({signal_5021, signal_5019}), .clk (CLK), .r (Fresh[439]), .c ({signal_2714, signal_1712}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1568 ( .s ({signal_5025, signal_5023}), .b ({signal_2530, signal_1572}), .a ({signal_2531, signal_1573}), .clk (CLK), .r (Fresh[440]), .c ({signal_2715, signal_1713}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1569 ( .s ({signal_4795, signal_4787}), .b ({signal_2498, signal_1655}), .a ({signal_2497, signal_1654}), .clk (CLK), .r (Fresh[441]), .c ({signal_2632, signal_919}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1570 ( .s ({signal_4831, signal_4827}), .b ({signal_2595, signal_1657}), .a ({signal_2594, signal_1656}), .clk (CLK), .r (Fresh[442]), .c ({signal_2716, signal_1714}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1571 ( .s ({signal_5057, signal_5055}), .b ({signal_5065, signal_5063}), .a ({signal_2563, signal_1615}), .clk (CLK), .r (Fresh[443]), .c ({signal_2717, signal_1715}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1572 ( .s ({signal_5057, signal_5055}), .b ({signal_5061, signal_5059}), .a ({signal_2565, signal_1617}), .clk (CLK), .r (Fresh[444]), .c ({signal_2718, signal_1716}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1573 ( .s ({signal_4831, signal_4827}), .b ({signal_2597, signal_1659}), .a ({signal_2596, signal_1658}), .clk (CLK), .r (Fresh[445]), .c ({signal_2719, signal_1717}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1574 ( .s ({signal_4831, signal_4827}), .b ({signal_2594, signal_1656}), .a ({signal_2595, signal_1657}), .clk (CLK), .r (Fresh[446]), .c ({signal_2720, signal_1718}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1575 ( .s ({signal_4831, signal_4827}), .b ({signal_2596, signal_1658}), .a ({signal_2597, signal_1659}), .clk (CLK), .r (Fresh[447]), .c ({signal_2721, signal_1719}) ) ;
    buf_clk cell_2197 ( .C (CLK), .D (signal_4340), .Q (signal_4341) ) ;
    buf_clk cell_2205 ( .C (CLK), .D (signal_4348), .Q (signal_4349) ) ;
    buf_clk cell_2213 ( .C (CLK), .D (signal_4356), .Q (signal_4357) ) ;
    buf_clk cell_2221 ( .C (CLK), .D (signal_4364), .Q (signal_4365) ) ;
    buf_clk cell_2229 ( .C (CLK), .D (signal_4372), .Q (signal_4373) ) ;
    buf_clk cell_2237 ( .C (CLK), .D (signal_4380), .Q (signal_4381) ) ;
    buf_clk cell_2245 ( .C (CLK), .D (signal_4388), .Q (signal_4389) ) ;
    buf_clk cell_2253 ( .C (CLK), .D (signal_4396), .Q (signal_4397) ) ;
    buf_clk cell_2261 ( .C (CLK), .D (signal_4404), .Q (signal_4405) ) ;
    buf_clk cell_2269 ( .C (CLK), .D (signal_4412), .Q (signal_4413) ) ;
    buf_clk cell_2273 ( .C (CLK), .D (signal_4416), .Q (signal_4417) ) ;
    buf_clk cell_2277 ( .C (CLK), .D (signal_4420), .Q (signal_4421) ) ;
    buf_clk cell_2285 ( .C (CLK), .D (signal_4428), .Q (signal_4429) ) ;
    buf_clk cell_2293 ( .C (CLK), .D (signal_4436), .Q (signal_4437) ) ;
    buf_clk cell_2297 ( .C (CLK), .D (signal_4440), .Q (signal_4441) ) ;
    buf_clk cell_2301 ( .C (CLK), .D (signal_4444), .Q (signal_4445) ) ;
    buf_clk cell_2305 ( .C (CLK), .D (signal_4448), .Q (signal_4449) ) ;
    buf_clk cell_2309 ( .C (CLK), .D (signal_4452), .Q (signal_4453) ) ;
    buf_clk cell_2317 ( .C (CLK), .D (signal_4460), .Q (signal_4461) ) ;
    buf_clk cell_2325 ( .C (CLK), .D (signal_4468), .Q (signal_4469) ) ;
    buf_clk cell_2333 ( .C (CLK), .D (signal_4476), .Q (signal_4477) ) ;
    buf_clk cell_2341 ( .C (CLK), .D (signal_4484), .Q (signal_4485) ) ;
    buf_clk cell_2345 ( .C (CLK), .D (signal_4488), .Q (signal_4489) ) ;
    buf_clk cell_2349 ( .C (CLK), .D (signal_4492), .Q (signal_4493) ) ;
    buf_clk cell_2357 ( .C (CLK), .D (signal_4500), .Q (signal_4501) ) ;
    buf_clk cell_2363 ( .C (CLK), .D (signal_4506), .Q (signal_4507) ) ;
    buf_clk cell_2369 ( .C (CLK), .D (signal_4512), .Q (signal_4513) ) ;
    buf_clk cell_2377 ( .C (CLK), .D (signal_4520), .Q (signal_4521) ) ;
    buf_clk cell_2385 ( .C (CLK), .D (signal_4528), .Q (signal_4529) ) ;
    buf_clk cell_2393 ( .C (CLK), .D (signal_4536), .Q (signal_4537) ) ;
    buf_clk cell_2401 ( .C (CLK), .D (signal_4544), .Q (signal_4545) ) ;
    buf_clk cell_2409 ( .C (CLK), .D (signal_4552), .Q (signal_4553) ) ;
    buf_clk cell_2417 ( .C (CLK), .D (signal_4560), .Q (signal_4561) ) ;
    buf_clk cell_2425 ( .C (CLK), .D (signal_4568), .Q (signal_4569) ) ;
    buf_clk cell_2433 ( .C (CLK), .D (signal_4576), .Q (signal_4577) ) ;
    buf_clk cell_2441 ( .C (CLK), .D (signal_4584), .Q (signal_4585) ) ;
    buf_clk cell_2449 ( .C (CLK), .D (signal_4592), .Q (signal_4593) ) ;
    buf_clk cell_2457 ( .C (CLK), .D (signal_4600), .Q (signal_4601) ) ;
    buf_clk cell_2465 ( .C (CLK), .D (signal_4608), .Q (signal_4609) ) ;
    buf_clk cell_2473 ( .C (CLK), .D (signal_4616), .Q (signal_4617) ) ;
    buf_clk cell_2481 ( .C (CLK), .D (signal_4624), .Q (signal_4625) ) ;
    buf_clk cell_2489 ( .C (CLK), .D (signal_4632), .Q (signal_4633) ) ;
    buf_clk cell_2497 ( .C (CLK), .D (signal_4640), .Q (signal_4641) ) ;
    buf_clk cell_2505 ( .C (CLK), .D (signal_4648), .Q (signal_4649) ) ;
    buf_clk cell_2513 ( .C (CLK), .D (signal_4656), .Q (signal_4657) ) ;
    buf_clk cell_2521 ( .C (CLK), .D (signal_4664), .Q (signal_4665) ) ;
    buf_clk cell_2529 ( .C (CLK), .D (signal_4672), .Q (signal_4673) ) ;
    buf_clk cell_2537 ( .C (CLK), .D (signal_4680), .Q (signal_4681) ) ;
    buf_clk cell_2545 ( .C (CLK), .D (signal_4688), .Q (signal_4689) ) ;
    buf_clk cell_2553 ( .C (CLK), .D (signal_4696), .Q (signal_4697) ) ;
    buf_clk cell_2561 ( .C (CLK), .D (signal_4704), .Q (signal_4705) ) ;
    buf_clk cell_2569 ( .C (CLK), .D (signal_4712), .Q (signal_4713) ) ;
    buf_clk cell_2573 ( .C (CLK), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_2577 ( .C (CLK), .D (signal_4720), .Q (signal_4721) ) ;
    buf_clk cell_2581 ( .C (CLK), .D (signal_4724), .Q (signal_4725) ) ;
    buf_clk cell_2585 ( .C (CLK), .D (signal_4728), .Q (signal_4729) ) ;
    buf_clk cell_2593 ( .C (CLK), .D (signal_4736), .Q (signal_4737) ) ;
    buf_clk cell_2601 ( .C (CLK), .D (signal_4744), .Q (signal_4745) ) ;
    buf_clk cell_2609 ( .C (CLK), .D (signal_4752), .Q (signal_4753) ) ;
    buf_clk cell_2617 ( .C (CLK), .D (signal_4760), .Q (signal_4761) ) ;
    buf_clk cell_2621 ( .C (CLK), .D (signal_4764), .Q (signal_4765) ) ;
    buf_clk cell_2625 ( .C (CLK), .D (signal_4768), .Q (signal_4769) ) ;
    buf_clk cell_2631 ( .C (CLK), .D (signal_4774), .Q (signal_4775) ) ;
    buf_clk cell_2637 ( .C (CLK), .D (signal_4780), .Q (signal_4781) ) ;
    buf_clk cell_2645 ( .C (CLK), .D (signal_4788), .Q (signal_4789) ) ;
    buf_clk cell_2653 ( .C (CLK), .D (signal_4796), .Q (signal_4797) ) ;
    buf_clk cell_2661 ( .C (CLK), .D (signal_4804), .Q (signal_4805) ) ;
    buf_clk cell_2669 ( .C (CLK), .D (signal_4812), .Q (signal_4813) ) ;
    buf_clk cell_2675 ( .C (CLK), .D (signal_4818), .Q (signal_4819) ) ;
    buf_clk cell_2681 ( .C (CLK), .D (signal_4824), .Q (signal_4825) ) ;
    buf_clk cell_2685 ( .C (CLK), .D (signal_4828), .Q (signal_4829) ) ;
    buf_clk cell_2689 ( .C (CLK), .D (signal_4832), .Q (signal_4833) ) ;
    buf_clk cell_2697 ( .C (CLK), .D (signal_4840), .Q (signal_4841) ) ;
    buf_clk cell_2705 ( .C (CLK), .D (signal_4848), .Q (signal_4849) ) ;
    buf_clk cell_2713 ( .C (CLK), .D (signal_4856), .Q (signal_4857) ) ;
    buf_clk cell_2721 ( .C (CLK), .D (signal_4864), .Q (signal_4865) ) ;
    buf_clk cell_2729 ( .C (CLK), .D (signal_4872), .Q (signal_4873) ) ;
    buf_clk cell_2737 ( .C (CLK), .D (signal_4880), .Q (signal_4881) ) ;
    buf_clk cell_2745 ( .C (CLK), .D (signal_4888), .Q (signal_4889) ) ;
    buf_clk cell_2753 ( .C (CLK), .D (signal_4896), .Q (signal_4897) ) ;
    buf_clk cell_2761 ( .C (CLK), .D (signal_4904), .Q (signal_4905) ) ;
    buf_clk cell_2769 ( .C (CLK), .D (signal_4912), .Q (signal_4913) ) ;
    buf_clk cell_2777 ( .C (CLK), .D (signal_4920), .Q (signal_4921) ) ;
    buf_clk cell_2785 ( .C (CLK), .D (signal_4928), .Q (signal_4929) ) ;
    buf_clk cell_3011 ( .C (CLK), .D (signal_5154), .Q (signal_5155) ) ;
    buf_clk cell_3013 ( .C (CLK), .D (signal_5156), .Q (signal_5157) ) ;
    buf_clk cell_3019 ( .C (CLK), .D (signal_5162), .Q (signal_5163) ) ;
    buf_clk cell_3025 ( .C (CLK), .D (signal_5168), .Q (signal_5169) ) ;
    buf_clk cell_3027 ( .C (CLK), .D (signal_5170), .Q (signal_5171) ) ;
    buf_clk cell_3029 ( .C (CLK), .D (signal_5172), .Q (signal_5173) ) ;
    buf_clk cell_3031 ( .C (CLK), .D (signal_5174), .Q (signal_5175) ) ;
    buf_clk cell_3033 ( .C (CLK), .D (signal_5176), .Q (signal_5177) ) ;
    buf_clk cell_3035 ( .C (CLK), .D (signal_5178), .Q (signal_5179) ) ;
    buf_clk cell_3037 ( .C (CLK), .D (signal_5180), .Q (signal_5181) ) ;
    buf_clk cell_3039 ( .C (CLK), .D (signal_5182), .Q (signal_5183) ) ;
    buf_clk cell_3041 ( .C (CLK), .D (signal_5184), .Q (signal_5185) ) ;
    buf_clk cell_3043 ( .C (CLK), .D (signal_5186), .Q (signal_5187) ) ;
    buf_clk cell_3045 ( .C (CLK), .D (signal_5188), .Q (signal_5189) ) ;
    buf_clk cell_3047 ( .C (CLK), .D (signal_5190), .Q (signal_5191) ) ;
    buf_clk cell_3049 ( .C (CLK), .D (signal_5192), .Q (signal_5193) ) ;
    buf_clk cell_3051 ( .C (CLK), .D (signal_5194), .Q (signal_5195) ) ;
    buf_clk cell_3053 ( .C (CLK), .D (signal_5196), .Q (signal_5197) ) ;
    buf_clk cell_3061 ( .C (CLK), .D (signal_5204), .Q (signal_5205) ) ;
    buf_clk cell_3069 ( .C (CLK), .D (signal_5212), .Q (signal_5213) ) ;
    buf_clk cell_3071 ( .C (CLK), .D (signal_5214), .Q (signal_5215) ) ;
    buf_clk cell_3073 ( .C (CLK), .D (signal_5216), .Q (signal_5217) ) ;
    buf_clk cell_3075 ( .C (CLK), .D (signal_5218), .Q (signal_5219) ) ;
    buf_clk cell_3077 ( .C (CLK), .D (signal_5220), .Q (signal_5221) ) ;
    buf_clk cell_3079 ( .C (CLK), .D (signal_5222), .Q (signal_5223) ) ;
    buf_clk cell_3081 ( .C (CLK), .D (signal_5224), .Q (signal_5225) ) ;
    buf_clk cell_3083 ( .C (CLK), .D (signal_5226), .Q (signal_5227) ) ;
    buf_clk cell_3085 ( .C (CLK), .D (signal_5228), .Q (signal_5229) ) ;
    buf_clk cell_3089 ( .C (CLK), .D (signal_5232), .Q (signal_5233) ) ;
    buf_clk cell_3093 ( .C (CLK), .D (signal_5236), .Q (signal_5237) ) ;
    buf_clk cell_3095 ( .C (CLK), .D (signal_5238), .Q (signal_5239) ) ;
    buf_clk cell_3097 ( .C (CLK), .D (signal_5240), .Q (signal_5241) ) ;
    buf_clk cell_3099 ( .C (CLK), .D (signal_5242), .Q (signal_5243) ) ;
    buf_clk cell_3101 ( .C (CLK), .D (signal_5244), .Q (signal_5245) ) ;
    buf_clk cell_3103 ( .C (CLK), .D (signal_5246), .Q (signal_5247) ) ;
    buf_clk cell_3105 ( .C (CLK), .D (signal_5248), .Q (signal_5249) ) ;
    buf_clk cell_3107 ( .C (CLK), .D (signal_5250), .Q (signal_5251) ) ;
    buf_clk cell_3109 ( .C (CLK), .D (signal_5252), .Q (signal_5253) ) ;
    buf_clk cell_3111 ( .C (CLK), .D (signal_5254), .Q (signal_5255) ) ;
    buf_clk cell_3113 ( .C (CLK), .D (signal_5256), .Q (signal_5257) ) ;
    buf_clk cell_3115 ( .C (CLK), .D (signal_5258), .Q (signal_5259) ) ;
    buf_clk cell_3117 ( .C (CLK), .D (signal_5260), .Q (signal_5261) ) ;
    buf_clk cell_3119 ( .C (CLK), .D (signal_5262), .Q (signal_5263) ) ;
    buf_clk cell_3121 ( .C (CLK), .D (signal_5264), .Q (signal_5265) ) ;
    buf_clk cell_3123 ( .C (CLK), .D (signal_5266), .Q (signal_5267) ) ;
    buf_clk cell_3125 ( .C (CLK), .D (signal_5268), .Q (signal_5269) ) ;
    buf_clk cell_3127 ( .C (CLK), .D (signal_5270), .Q (signal_5271) ) ;
    buf_clk cell_3129 ( .C (CLK), .D (signal_5272), .Q (signal_5273) ) ;
    buf_clk cell_3199 ( .C (CLK), .D (signal_5342), .Q (signal_5343) ) ;
    buf_clk cell_3207 ( .C (CLK), .D (signal_5350), .Q (signal_5351) ) ;
    buf_clk cell_3231 ( .C (CLK), .D (signal_5374), .Q (signal_5375) ) ;
    buf_clk cell_3235 ( .C (CLK), .D (signal_5378), .Q (signal_5379) ) ;
    buf_clk cell_3299 ( .C (CLK), .D (signal_5442), .Q (signal_5443) ) ;
    buf_clk cell_3305 ( .C (CLK), .D (signal_5448), .Q (signal_5449) ) ;
    buf_clk cell_3321 ( .C (CLK), .D (signal_5464), .Q (signal_5465) ) ;
    buf_clk cell_3329 ( .C (CLK), .D (signal_5472), .Q (signal_5473) ) ;
    buf_clk cell_3339 ( .C (CLK), .D (signal_5482), .Q (signal_5483) ) ;
    buf_clk cell_3345 ( .C (CLK), .D (signal_5488), .Q (signal_5489) ) ;
    buf_clk cell_3357 ( .C (CLK), .D (signal_5500), .Q (signal_5501) ) ;
    buf_clk cell_3365 ( .C (CLK), .D (signal_5508), .Q (signal_5509) ) ;
    buf_clk cell_3453 ( .C (CLK), .D (signal_5596), .Q (signal_5597) ) ;
    buf_clk cell_3469 ( .C (CLK), .D (signal_5612), .Q (signal_5613) ) ;
    buf_clk cell_3493 ( .C (CLK), .D (signal_5636), .Q (signal_5637) ) ;
    buf_clk cell_3509 ( .C (CLK), .D (signal_5652), .Q (signal_5653) ) ;
    buf_clk cell_3533 ( .C (CLK), .D (signal_5676), .Q (signal_5677) ) ;
    buf_clk cell_3549 ( .C (CLK), .D (signal_5692), .Q (signal_5693) ) ;
    buf_clk cell_3565 ( .C (CLK), .D (signal_5708), .Q (signal_5709) ) ;
    buf_clk cell_3581 ( .C (CLK), .D (signal_5724), .Q (signal_5725) ) ;
    buf_clk cell_3641 ( .C (CLK), .D (signal_5784), .Q (signal_5785) ) ;
    buf_clk cell_3657 ( .C (CLK), .D (signal_5800), .Q (signal_5801) ) ;
    buf_clk cell_3673 ( .C (CLK), .D (signal_5816), .Q (signal_5817) ) ;
    buf_clk cell_3689 ( .C (CLK), .D (signal_5832), .Q (signal_5833) ) ;
    buf_clk cell_3705 ( .C (CLK), .D (signal_5848), .Q (signal_5849) ) ;
    buf_clk cell_3721 ( .C (CLK), .D (signal_5864), .Q (signal_5865) ) ;
    buf_clk cell_3737 ( .C (CLK), .D (signal_5880), .Q (signal_5881) ) ;
    buf_clk cell_3753 ( .C (CLK), .D (signal_5896), .Q (signal_5897) ) ;
    buf_clk cell_3769 ( .C (CLK), .D (signal_5912), .Q (signal_5913) ) ;
    buf_clk cell_3785 ( .C (CLK), .D (signal_5928), .Q (signal_5929) ) ;
    buf_clk cell_3893 ( .C (CLK), .D (signal_6036), .Q (signal_6037) ) ;
    buf_clk cell_3909 ( .C (CLK), .D (signal_6052), .Q (signal_6053) ) ;
    buf_clk cell_3925 ( .C (CLK), .D (signal_6068), .Q (signal_6069) ) ;
    buf_clk cell_3941 ( .C (CLK), .D (signal_6084), .Q (signal_6085) ) ;
    buf_clk cell_3957 ( .C (CLK), .D (signal_6100), .Q (signal_6101) ) ;
    buf_clk cell_3973 ( .C (CLK), .D (signal_6116), .Q (signal_6117) ) ;
    buf_clk cell_3989 ( .C (CLK), .D (signal_6132), .Q (signal_6133) ) ;
    buf_clk cell_4005 ( .C (CLK), .D (signal_6148), .Q (signal_6149) ) ;
    buf_clk cell_4021 ( .C (CLK), .D (signal_6164), .Q (signal_6165) ) ;
    buf_clk cell_4037 ( .C (CLK), .D (signal_6180), .Q (signal_6181) ) ;
    buf_clk cell_4053 ( .C (CLK), .D (signal_6196), .Q (signal_6197) ) ;
    buf_clk cell_4069 ( .C (CLK), .D (signal_6212), .Q (signal_6213) ) ;
    buf_clk cell_4085 ( .C (CLK), .D (signal_6228), .Q (signal_6229) ) ;
    buf_clk cell_4101 ( .C (CLK), .D (signal_6244), .Q (signal_6245) ) ;
    buf_clk cell_4111 ( .C (CLK), .D (signal_6254), .Q (signal_6255) ) ;
    buf_clk cell_4121 ( .C (CLK), .D (signal_6264), .Q (signal_6265) ) ;
    buf_clk cell_4159 ( .C (CLK), .D (signal_6302), .Q (signal_6303) ) ;
    buf_clk cell_4169 ( .C (CLK), .D (signal_6312), .Q (signal_6313) ) ;
    buf_clk cell_4185 ( .C (CLK), .D (signal_6328), .Q (signal_6329) ) ;
    buf_clk cell_4197 ( .C (CLK), .D (signal_6340), .Q (signal_6341) ) ;
    buf_clk cell_4209 ( .C (CLK), .D (signal_6352), .Q (signal_6353) ) ;
    buf_clk cell_4237 ( .C (CLK), .D (signal_6380), .Q (signal_6381) ) ;
    buf_clk cell_4249 ( .C (CLK), .D (signal_6392), .Q (signal_6393) ) ;
    buf_clk cell_4263 ( .C (CLK), .D (signal_6406), .Q (signal_6407) ) ;
    buf_clk cell_4277 ( .C (CLK), .D (signal_6420), .Q (signal_6421) ) ;
    buf_clk cell_4293 ( .C (CLK), .D (signal_6436), .Q (signal_6437) ) ;
    buf_clk cell_4309 ( .C (CLK), .D (signal_6452), .Q (signal_6453) ) ;
    buf_clk cell_4325 ( .C (CLK), .D (signal_6468), .Q (signal_6469) ) ;
    buf_clk cell_4341 ( .C (CLK), .D (signal_6484), .Q (signal_6485) ) ;
    buf_clk cell_4357 ( .C (CLK), .D (signal_6500), .Q (signal_6501) ) ;
    buf_clk cell_4373 ( .C (CLK), .D (signal_6516), .Q (signal_6517) ) ;
    buf_clk cell_4389 ( .C (CLK), .D (signal_6532), .Q (signal_6533) ) ;
    buf_clk cell_4405 ( .C (CLK), .D (signal_6548), .Q (signal_6549) ) ;
    buf_clk cell_4421 ( .C (CLK), .D (signal_6564), .Q (signal_6565) ) ;
    buf_clk cell_4437 ( .C (CLK), .D (signal_6580), .Q (signal_6581) ) ;
    buf_clk cell_4453 ( .C (CLK), .D (signal_6596), .Q (signal_6597) ) ;
    buf_clk cell_4469 ( .C (CLK), .D (signal_6612), .Q (signal_6613) ) ;
    buf_clk cell_4485 ( .C (CLK), .D (signal_6628), .Q (signal_6629) ) ;
    buf_clk cell_4501 ( .C (CLK), .D (signal_6644), .Q (signal_6645) ) ;
    buf_clk cell_4517 ( .C (CLK), .D (signal_6660), .Q (signal_6661) ) ;
    buf_clk cell_4533 ( .C (CLK), .D (signal_6676), .Q (signal_6677) ) ;
    buf_clk cell_4543 ( .C (CLK), .D (signal_6686), .Q (signal_6687) ) ;
    buf_clk cell_4553 ( .C (CLK), .D (signal_6696), .Q (signal_6697) ) ;
    buf_clk cell_4581 ( .C (CLK), .D (signal_6724), .Q (signal_6725) ) ;
    buf_clk cell_4593 ( .C (CLK), .D (signal_6736), .Q (signal_6737) ) ;
    buf_clk cell_4607 ( .C (CLK), .D (signal_6750), .Q (signal_6751) ) ;
    buf_clk cell_4621 ( .C (CLK), .D (signal_6764), .Q (signal_6765) ) ;
    buf_clk cell_4637 ( .C (CLK), .D (signal_6780), .Q (signal_6781) ) ;
    buf_clk cell_4653 ( .C (CLK), .D (signal_6796), .Q (signal_6797) ) ;
    buf_clk cell_4691 ( .C (CLK), .D (signal_6834), .Q (signal_6835) ) ;
    buf_clk cell_4701 ( .C (CLK), .D (signal_6844), .Q (signal_6845) ) ;
    buf_clk cell_4713 ( .C (CLK), .D (signal_6856), .Q (signal_6857) ) ;
    buf_clk cell_4725 ( .C (CLK), .D (signal_6868), .Q (signal_6869) ) ;
    buf_clk cell_4749 ( .C (CLK), .D (signal_6892), .Q (signal_6893) ) ;
    buf_clk cell_4765 ( .C (CLK), .D (signal_6908), .Q (signal_6909) ) ;
    buf_clk cell_4781 ( .C (CLK), .D (signal_6924), .Q (signal_6925) ) ;
    buf_clk cell_4797 ( .C (CLK), .D (signal_6940), .Q (signal_6941) ) ;
    buf_clk cell_4813 ( .C (CLK), .D (signal_6956), .Q (signal_6957) ) ;
    buf_clk cell_4829 ( .C (CLK), .D (signal_6972), .Q (signal_6973) ) ;
    buf_clk cell_4845 ( .C (CLK), .D (signal_6988), .Q (signal_6989) ) ;
    buf_clk cell_4861 ( .C (CLK), .D (signal_7004), .Q (signal_7005) ) ;
    buf_clk cell_4877 ( .C (CLK), .D (signal_7020), .Q (signal_7021) ) ;
    buf_clk cell_4893 ( .C (CLK), .D (signal_7036), .Q (signal_7037) ) ;
    buf_clk cell_4909 ( .C (CLK), .D (signal_7052), .Q (signal_7053) ) ;
    buf_clk cell_4925 ( .C (CLK), .D (signal_7068), .Q (signal_7069) ) ;
    buf_clk cell_4941 ( .C (CLK), .D (signal_7084), .Q (signal_7085) ) ;
    buf_clk cell_4957 ( .C (CLK), .D (signal_7100), .Q (signal_7101) ) ;
    buf_clk cell_4973 ( .C (CLK), .D (signal_7116), .Q (signal_7117) ) ;
    buf_clk cell_4989 ( .C (CLK), .D (signal_7132), .Q (signal_7133) ) ;
    buf_clk cell_5005 ( .C (CLK), .D (signal_7148), .Q (signal_7149) ) ;
    buf_clk cell_5021 ( .C (CLK), .D (signal_7164), .Q (signal_7165) ) ;
    buf_clk cell_5037 ( .C (CLK), .D (signal_7180), .Q (signal_7181) ) ;
    buf_clk cell_5053 ( .C (CLK), .D (signal_7196), .Q (signal_7197) ) ;
    buf_clk cell_5069 ( .C (CLK), .D (signal_7212), .Q (signal_7213) ) ;
    buf_clk cell_5085 ( .C (CLK), .D (signal_7228), .Q (signal_7229) ) ;
    buf_clk cell_5101 ( .C (CLK), .D (signal_7244), .Q (signal_7245) ) ;
    buf_clk cell_5117 ( .C (CLK), .D (signal_7260), .Q (signal_7261) ) ;
    buf_clk cell_5133 ( .C (CLK), .D (signal_7276), .Q (signal_7277) ) ;
    buf_clk cell_5149 ( .C (CLK), .D (signal_7292), .Q (signal_7293) ) ;
    buf_clk cell_5165 ( .C (CLK), .D (signal_7308), .Q (signal_7309) ) ;
    buf_clk cell_5181 ( .C (CLK), .D (signal_7324), .Q (signal_7325) ) ;
    buf_clk cell_5197 ( .C (CLK), .D (signal_7340), .Q (signal_7341) ) ;
    buf_clk cell_5213 ( .C (CLK), .D (signal_7356), .Q (signal_7357) ) ;
    buf_clk cell_5229 ( .C (CLK), .D (signal_7372), .Q (signal_7373) ) ;
    buf_clk cell_5245 ( .C (CLK), .D (signal_7388), .Q (signal_7389) ) ;
    buf_clk cell_5261 ( .C (CLK), .D (signal_7404), .Q (signal_7405) ) ;
    buf_clk cell_5277 ( .C (CLK), .D (signal_7420), .Q (signal_7421) ) ;
    buf_clk cell_5293 ( .C (CLK), .D (signal_7436), .Q (signal_7437) ) ;
    buf_clk cell_5309 ( .C (CLK), .D (signal_7452), .Q (signal_7453) ) ;
    buf_clk cell_5325 ( .C (CLK), .D (signal_7468), .Q (signal_7469) ) ;
    buf_clk cell_5341 ( .C (CLK), .D (signal_7484), .Q (signal_7485) ) ;
    buf_clk cell_5357 ( .C (CLK), .D (signal_7500), .Q (signal_7501) ) ;
    buf_clk cell_5373 ( .C (CLK), .D (signal_7516), .Q (signal_7517) ) ;
    buf_clk cell_5389 ( .C (CLK), .D (signal_7532), .Q (signal_7533) ) ;
    buf_clk cell_5405 ( .C (CLK), .D (signal_7548), .Q (signal_7549) ) ;
    buf_clk cell_5421 ( .C (CLK), .D (signal_7564), .Q (signal_7565) ) ;
    buf_clk cell_5437 ( .C (CLK), .D (signal_7580), .Q (signal_7581) ) ;
    buf_clk cell_5453 ( .C (CLK), .D (signal_7596), .Q (signal_7597) ) ;
    buf_clk cell_5469 ( .C (CLK), .D (signal_7612), .Q (signal_7613) ) ;
    buf_clk cell_5485 ( .C (CLK), .D (signal_7628), .Q (signal_7629) ) ;
    buf_clk cell_5501 ( .C (CLK), .D (signal_7644), .Q (signal_7645) ) ;
    buf_clk cell_5517 ( .C (CLK), .D (signal_7660), .Q (signal_7661) ) ;
    buf_clk cell_5533 ( .C (CLK), .D (signal_7676), .Q (signal_7677) ) ;
    buf_clk cell_5549 ( .C (CLK), .D (signal_7692), .Q (signal_7693) ) ;
    buf_clk cell_5565 ( .C (CLK), .D (signal_7708), .Q (signal_7709) ) ;
    buf_clk cell_5581 ( .C (CLK), .D (signal_7724), .Q (signal_7725) ) ;
    buf_clk cell_5597 ( .C (CLK), .D (signal_7740), .Q (signal_7741) ) ;
    buf_clk cell_5613 ( .C (CLK), .D (signal_7756), .Q (signal_7757) ) ;
    buf_clk cell_5629 ( .C (CLK), .D (signal_7772), .Q (signal_7773) ) ;
    buf_clk cell_5645 ( .C (CLK), .D (signal_7788), .Q (signal_7789) ) ;
    buf_clk cell_5661 ( .C (CLK), .D (signal_7804), .Q (signal_7805) ) ;
    buf_clk cell_5677 ( .C (CLK), .D (signal_7820), .Q (signal_7821) ) ;
    buf_clk cell_5693 ( .C (CLK), .D (signal_7836), .Q (signal_7837) ) ;
    buf_clk cell_5709 ( .C (CLK), .D (signal_7852), .Q (signal_7853) ) ;
    buf_clk cell_5725 ( .C (CLK), .D (signal_7868), .Q (signal_7869) ) ;
    buf_clk cell_5741 ( .C (CLK), .D (signal_7884), .Q (signal_7885) ) ;
    buf_clk cell_5757 ( .C (CLK), .D (signal_7900), .Q (signal_7901) ) ;
    buf_clk cell_5773 ( .C (CLK), .D (signal_7916), .Q (signal_7917) ) ;
    buf_clk cell_5789 ( .C (CLK), .D (signal_7932), .Q (signal_7933) ) ;
    buf_clk cell_5805 ( .C (CLK), .D (signal_7948), .Q (signal_7949) ) ;
    buf_clk cell_5821 ( .C (CLK), .D (signal_7964), .Q (signal_7965) ) ;
    buf_clk cell_5837 ( .C (CLK), .D (signal_7980), .Q (signal_7981) ) ;
    buf_clk cell_5853 ( .C (CLK), .D (signal_7996), .Q (signal_7997) ) ;
    buf_clk cell_5869 ( .C (CLK), .D (signal_8012), .Q (signal_8013) ) ;
    buf_clk cell_5885 ( .C (CLK), .D (signal_8028), .Q (signal_8029) ) ;
    buf_clk cell_5901 ( .C (CLK), .D (signal_8044), .Q (signal_8045) ) ;
    buf_clk cell_5917 ( .C (CLK), .D (signal_8060), .Q (signal_8061) ) ;
    buf_clk cell_5933 ( .C (CLK), .D (signal_8076), .Q (signal_8077) ) ;
    buf_clk cell_5949 ( .C (CLK), .D (signal_8092), .Q (signal_8093) ) ;
    buf_clk cell_5965 ( .C (CLK), .D (signal_8108), .Q (signal_8109) ) ;
    buf_clk cell_5981 ( .C (CLK), .D (signal_8124), .Q (signal_8125) ) ;
    buf_clk cell_5997 ( .C (CLK), .D (signal_8140), .Q (signal_8141) ) ;
    buf_clk cell_6013 ( .C (CLK), .D (signal_8156), .Q (signal_8157) ) ;
    buf_clk cell_6029 ( .C (CLK), .D (signal_8172), .Q (signal_8173) ) ;
    buf_clk cell_6045 ( .C (CLK), .D (signal_8188), .Q (signal_8189) ) ;
    buf_clk cell_6061 ( .C (CLK), .D (signal_8204), .Q (signal_8205) ) ;
    buf_clk cell_6077 ( .C (CLK), .D (signal_8220), .Q (signal_8221) ) ;
    buf_clk cell_6093 ( .C (CLK), .D (signal_8236), .Q (signal_8237) ) ;
    buf_clk cell_6109 ( .C (CLK), .D (signal_8252), .Q (signal_8253) ) ;
    buf_clk cell_6125 ( .C (CLK), .D (signal_8268), .Q (signal_8269) ) ;
    buf_clk cell_6141 ( .C (CLK), .D (signal_8284), .Q (signal_8285) ) ;
    buf_clk cell_6157 ( .C (CLK), .D (signal_8300), .Q (signal_8301) ) ;
    buf_clk cell_6173 ( .C (CLK), .D (signal_8316), .Q (signal_8317) ) ;
    buf_clk cell_6189 ( .C (CLK), .D (signal_8332), .Q (signal_8333) ) ;
    buf_clk cell_6205 ( .C (CLK), .D (signal_8348), .Q (signal_8349) ) ;
    buf_clk cell_6221 ( .C (CLK), .D (signal_8364), .Q (signal_8365) ) ;
    buf_clk cell_6237 ( .C (CLK), .D (signal_8380), .Q (signal_8381) ) ;
    buf_clk cell_6253 ( .C (CLK), .D (signal_8396), .Q (signal_8397) ) ;
    buf_clk cell_6269 ( .C (CLK), .D (signal_8412), .Q (signal_8413) ) ;
    buf_clk cell_6285 ( .C (CLK), .D (signal_8428), .Q (signal_8429) ) ;
    buf_clk cell_6301 ( .C (CLK), .D (signal_8444), .Q (signal_8445) ) ;
    buf_clk cell_6317 ( .C (CLK), .D (signal_8460), .Q (signal_8461) ) ;
    buf_clk cell_6333 ( .C (CLK), .D (signal_8476), .Q (signal_8477) ) ;
    buf_clk cell_6349 ( .C (CLK), .D (signal_8492), .Q (signal_8493) ) ;
    buf_clk cell_6365 ( .C (CLK), .D (signal_8508), .Q (signal_8509) ) ;
    buf_clk cell_6381 ( .C (CLK), .D (signal_8524), .Q (signal_8525) ) ;
    buf_clk cell_6397 ( .C (CLK), .D (signal_8540), .Q (signal_8541) ) ;
    buf_clk cell_7563 ( .C (CLK), .D (signal_9706), .Q (signal_9707) ) ;
    buf_clk cell_7571 ( .C (CLK), .D (signal_9714), .Q (signal_9715) ) ;
    buf_clk cell_7597 ( .C (CLK), .D (signal_9740), .Q (signal_9741) ) ;
    buf_clk cell_7613 ( .C (CLK), .D (signal_9756), .Q (signal_9757) ) ;
    buf_clk cell_7629 ( .C (CLK), .D (signal_9772), .Q (signal_9773) ) ;
    buf_clk cell_7645 ( .C (CLK), .D (signal_9788), .Q (signal_9789) ) ;
    buf_clk cell_7661 ( .C (CLK), .D (signal_9804), .Q (signal_9805) ) ;
    buf_clk cell_7677 ( .C (CLK), .D (signal_9820), .Q (signal_9821) ) ;
    buf_clk cell_7693 ( .C (CLK), .D (signal_9836), .Q (signal_9837) ) ;
    buf_clk cell_7709 ( .C (CLK), .D (signal_9852), .Q (signal_9853) ) ;
    buf_clk cell_7725 ( .C (CLK), .D (signal_9868), .Q (signal_9869) ) ;
    buf_clk cell_7741 ( .C (CLK), .D (signal_9884), .Q (signal_9885) ) ;
    buf_clk cell_7949 ( .C (CLK), .D (signal_10092), .Q (signal_10093) ) ;

    /* cells in depth 9 */
    buf_clk cell_3130 ( .C (CLK), .D (signal_5163), .Q (signal_5274) ) ;
    buf_clk cell_3132 ( .C (CLK), .D (signal_5169), .Q (signal_5276) ) ;
    buf_clk cell_3134 ( .C (CLK), .D (signal_898), .Q (signal_5278) ) ;
    buf_clk cell_3136 ( .C (CLK), .D (signal_2613), .Q (signal_5280) ) ;
    buf_clk cell_3138 ( .C (CLK), .D (signal_1660), .Q (signal_5282) ) ;
    buf_clk cell_3140 ( .C (CLK), .D (signal_2614), .Q (signal_5284) ) ;
    buf_clk cell_3142 ( .C (CLK), .D (signal_4841), .Q (signal_5286) ) ;
    buf_clk cell_3144 ( .C (CLK), .D (signal_4849), .Q (signal_5288) ) ;
    buf_clk cell_3146 ( .C (CLK), .D (signal_4717), .Q (signal_5290) ) ;
    buf_clk cell_3148 ( .C (CLK), .D (signal_4721), .Q (signal_5292) ) ;
    buf_clk cell_3150 ( .C (CLK), .D (signal_1672), .Q (signal_5294) ) ;
    buf_clk cell_3152 ( .C (CLK), .D (signal_2665), .Q (signal_5296) ) ;
    buf_clk cell_3154 ( .C (CLK), .D (signal_1676), .Q (signal_5298) ) ;
    buf_clk cell_3156 ( .C (CLK), .D (signal_2669), .Q (signal_5300) ) ;
    buf_clk cell_3158 ( .C (CLK), .D (signal_4507), .Q (signal_5302) ) ;
    buf_clk cell_3160 ( .C (CLK), .D (signal_4513), .Q (signal_5304) ) ;
    buf_clk cell_3162 ( .C (CLK), .D (signal_910), .Q (signal_5306) ) ;
    buf_clk cell_3164 ( .C (CLK), .D (signal_2674), .Q (signal_5308) ) ;
    buf_clk cell_3166 ( .C (CLK), .D (signal_1678), .Q (signal_5310) ) ;
    buf_clk cell_3168 ( .C (CLK), .D (signal_2678), .Q (signal_5312) ) ;
    buf_clk cell_3170 ( .C (CLK), .D (signal_4765), .Q (signal_5314) ) ;
    buf_clk cell_3172 ( .C (CLK), .D (signal_4769), .Q (signal_5316) ) ;
    buf_clk cell_3174 ( .C (CLK), .D (signal_1679), .Q (signal_5318) ) ;
    buf_clk cell_3176 ( .C (CLK), .D (signal_2682), .Q (signal_5320) ) ;
    buf_clk cell_3178 ( .C (CLK), .D (signal_1682), .Q (signal_5322) ) ;
    buf_clk cell_3180 ( .C (CLK), .D (signal_2685), .Q (signal_5324) ) ;
    buf_clk cell_3182 ( .C (CLK), .D (signal_1683), .Q (signal_5326) ) ;
    buf_clk cell_3184 ( .C (CLK), .D (signal_2686), .Q (signal_5328) ) ;
    buf_clk cell_3186 ( .C (CLK), .D (signal_1684), .Q (signal_5330) ) ;
    buf_clk cell_3188 ( .C (CLK), .D (signal_2687), .Q (signal_5332) ) ;
    buf_clk cell_3190 ( .C (CLK), .D (signal_4921), .Q (signal_5334) ) ;
    buf_clk cell_3192 ( .C (CLK), .D (signal_4929), .Q (signal_5336) ) ;
    buf_clk cell_3200 ( .C (CLK), .D (signal_5343), .Q (signal_5344) ) ;
    buf_clk cell_3208 ( .C (CLK), .D (signal_5351), .Q (signal_5352) ) ;
    buf_clk cell_3210 ( .C (CLK), .D (signal_4405), .Q (signal_5354) ) ;
    buf_clk cell_3212 ( .C (CLK), .D (signal_4413), .Q (signal_5356) ) ;
    buf_clk cell_3214 ( .C (CLK), .D (signal_5251), .Q (signal_5358) ) ;
    buf_clk cell_3216 ( .C (CLK), .D (signal_5253), .Q (signal_5360) ) ;
    buf_clk cell_3218 ( .C (CLK), .D (signal_4417), .Q (signal_5362) ) ;
    buf_clk cell_3220 ( .C (CLK), .D (signal_4421), .Q (signal_5364) ) ;
    buf_clk cell_3222 ( .C (CLK), .D (signal_1702), .Q (signal_5366) ) ;
    buf_clk cell_3224 ( .C (CLK), .D (signal_2625), .Q (signal_5368) ) ;
    buf_clk cell_3226 ( .C (CLK), .D (signal_1703), .Q (signal_5370) ) ;
    buf_clk cell_3228 ( .C (CLK), .D (signal_2626), .Q (signal_5372) ) ;
    buf_clk cell_3232 ( .C (CLK), .D (signal_5375), .Q (signal_5376) ) ;
    buf_clk cell_3236 ( .C (CLK), .D (signal_5379), .Q (signal_5380) ) ;
    buf_clk cell_3238 ( .C (CLK), .D (signal_4753), .Q (signal_5382) ) ;
    buf_clk cell_3240 ( .C (CLK), .D (signal_4761), .Q (signal_5384) ) ;
    buf_clk cell_3242 ( .C (CLK), .D (signal_899), .Q (signal_5386) ) ;
    buf_clk cell_3244 ( .C (CLK), .D (signal_2611), .Q (signal_5388) ) ;
    buf_clk cell_3246 ( .C (CLK), .D (signal_1709), .Q (signal_5390) ) ;
    buf_clk cell_3248 ( .C (CLK), .D (signal_2630), .Q (signal_5392) ) ;
    buf_clk cell_3250 ( .C (CLK), .D (signal_911), .Q (signal_5394) ) ;
    buf_clk cell_3252 ( .C (CLK), .D (signal_2676), .Q (signal_5396) ) ;
    buf_clk cell_3254 ( .C (CLK), .D (signal_1710), .Q (signal_5398) ) ;
    buf_clk cell_3256 ( .C (CLK), .D (signal_2710), .Q (signal_5400) ) ;
    buf_clk cell_3258 ( .C (CLK), .D (signal_1714), .Q (signal_5402) ) ;
    buf_clk cell_3260 ( .C (CLK), .D (signal_2716), .Q (signal_5404) ) ;
    buf_clk cell_3262 ( .C (CLK), .D (signal_1717), .Q (signal_5406) ) ;
    buf_clk cell_3264 ( .C (CLK), .D (signal_2719), .Q (signal_5408) ) ;
    buf_clk cell_3266 ( .C (CLK), .D (signal_1718), .Q (signal_5410) ) ;
    buf_clk cell_3268 ( .C (CLK), .D (signal_2720), .Q (signal_5412) ) ;
    buf_clk cell_3270 ( .C (CLK), .D (signal_1719), .Q (signal_5414) ) ;
    buf_clk cell_3272 ( .C (CLK), .D (signal_2721), .Q (signal_5416) ) ;
    buf_clk cell_3274 ( .C (CLK), .D (signal_4489), .Q (signal_5418) ) ;
    buf_clk cell_3278 ( .C (CLK), .D (signal_4493), .Q (signal_5422) ) ;
    buf_clk cell_3286 ( .C (CLK), .D (signal_5187), .Q (signal_5430) ) ;
    buf_clk cell_3290 ( .C (CLK), .D (signal_5189), .Q (signal_5434) ) ;
    buf_clk cell_3300 ( .C (CLK), .D (signal_5443), .Q (signal_5444) ) ;
    buf_clk cell_3306 ( .C (CLK), .D (signal_5449), .Q (signal_5450) ) ;
    buf_clk cell_3322 ( .C (CLK), .D (signal_5465), .Q (signal_5466) ) ;
    buf_clk cell_3330 ( .C (CLK), .D (signal_5473), .Q (signal_5474) ) ;
    buf_clk cell_3340 ( .C (CLK), .D (signal_5483), .Q (signal_5484) ) ;
    buf_clk cell_3346 ( .C (CLK), .D (signal_5489), .Q (signal_5490) ) ;
    buf_clk cell_3358 ( .C (CLK), .D (signal_5501), .Q (signal_5502) ) ;
    buf_clk cell_3366 ( .C (CLK), .D (signal_5509), .Q (signal_5510) ) ;
    buf_clk cell_3398 ( .C (CLK), .D (signal_4737), .Q (signal_5542) ) ;
    buf_clk cell_3402 ( .C (CLK), .D (signal_4745), .Q (signal_5546) ) ;
    buf_clk cell_3406 ( .C (CLK), .D (signal_4441), .Q (signal_5550) ) ;
    buf_clk cell_3410 ( .C (CLK), .D (signal_4445), .Q (signal_5554) ) ;
    buf_clk cell_3438 ( .C (CLK), .D (signal_4341), .Q (signal_5582) ) ;
    buf_clk cell_3454 ( .C (CLK), .D (signal_5597), .Q (signal_5598) ) ;
    buf_clk cell_3470 ( .C (CLK), .D (signal_5613), .Q (signal_5614) ) ;
    buf_clk cell_3478 ( .C (CLK), .D (signal_4501), .Q (signal_5622) ) ;
    buf_clk cell_3494 ( .C (CLK), .D (signal_5637), .Q (signal_5638) ) ;
    buf_clk cell_3510 ( .C (CLK), .D (signal_5653), .Q (signal_5654) ) ;
    buf_clk cell_3518 ( .C (CLK), .D (signal_4365), .Q (signal_5662) ) ;
    buf_clk cell_3534 ( .C (CLK), .D (signal_5677), .Q (signal_5678) ) ;
    buf_clk cell_3550 ( .C (CLK), .D (signal_5693), .Q (signal_5694) ) ;
    buf_clk cell_3566 ( .C (CLK), .D (signal_5709), .Q (signal_5710) ) ;
    buf_clk cell_3582 ( .C (CLK), .D (signal_5725), .Q (signal_5726) ) ;
    buf_clk cell_3642 ( .C (CLK), .D (signal_5785), .Q (signal_5786) ) ;
    buf_clk cell_3658 ( .C (CLK), .D (signal_5801), .Q (signal_5802) ) ;
    buf_clk cell_3674 ( .C (CLK), .D (signal_5817), .Q (signal_5818) ) ;
    buf_clk cell_3690 ( .C (CLK), .D (signal_5833), .Q (signal_5834) ) ;
    buf_clk cell_3706 ( .C (CLK), .D (signal_5849), .Q (signal_5850) ) ;
    buf_clk cell_3722 ( .C (CLK), .D (signal_5865), .Q (signal_5866) ) ;
    buf_clk cell_3738 ( .C (CLK), .D (signal_5881), .Q (signal_5882) ) ;
    buf_clk cell_3754 ( .C (CLK), .D (signal_5897), .Q (signal_5898) ) ;
    buf_clk cell_3770 ( .C (CLK), .D (signal_5913), .Q (signal_5914) ) ;
    buf_clk cell_3786 ( .C (CLK), .D (signal_5929), .Q (signal_5930) ) ;
    buf_clk cell_3802 ( .C (CLK), .D (signal_4789), .Q (signal_5946) ) ;
    buf_clk cell_3810 ( .C (CLK), .D (signal_4797), .Q (signal_5954) ) ;
    buf_clk cell_3830 ( .C (CLK), .D (signal_5155), .Q (signal_5974) ) ;
    buf_clk cell_3838 ( .C (CLK), .D (signal_5157), .Q (signal_5982) ) ;
    buf_clk cell_3846 ( .C (CLK), .D (signal_4805), .Q (signal_5990) ) ;
    buf_clk cell_3854 ( .C (CLK), .D (signal_4813), .Q (signal_5998) ) ;
    buf_clk cell_3870 ( .C (CLK), .D (signal_5205), .Q (signal_6014) ) ;
    buf_clk cell_3878 ( .C (CLK), .D (signal_5213), .Q (signal_6022) ) ;
    buf_clk cell_3894 ( .C (CLK), .D (signal_6037), .Q (signal_6038) ) ;
    buf_clk cell_3910 ( .C (CLK), .D (signal_6053), .Q (signal_6054) ) ;
    buf_clk cell_3926 ( .C (CLK), .D (signal_6069), .Q (signal_6070) ) ;
    buf_clk cell_3942 ( .C (CLK), .D (signal_6085), .Q (signal_6086) ) ;
    buf_clk cell_3958 ( .C (CLK), .D (signal_6101), .Q (signal_6102) ) ;
    buf_clk cell_3974 ( .C (CLK), .D (signal_6117), .Q (signal_6118) ) ;
    buf_clk cell_3990 ( .C (CLK), .D (signal_6133), .Q (signal_6134) ) ;
    buf_clk cell_4006 ( .C (CLK), .D (signal_6149), .Q (signal_6150) ) ;
    buf_clk cell_4022 ( .C (CLK), .D (signal_6165), .Q (signal_6166) ) ;
    buf_clk cell_4038 ( .C (CLK), .D (signal_6181), .Q (signal_6182) ) ;
    buf_clk cell_4054 ( .C (CLK), .D (signal_6197), .Q (signal_6198) ) ;
    buf_clk cell_4070 ( .C (CLK), .D (signal_6213), .Q (signal_6214) ) ;
    buf_clk cell_4086 ( .C (CLK), .D (signal_6229), .Q (signal_6230) ) ;
    buf_clk cell_4102 ( .C (CLK), .D (signal_6245), .Q (signal_6246) ) ;
    buf_clk cell_4112 ( .C (CLK), .D (signal_6255), .Q (signal_6256) ) ;
    buf_clk cell_4122 ( .C (CLK), .D (signal_6265), .Q (signal_6266) ) ;
    buf_clk cell_4142 ( .C (CLK), .D (signal_5171), .Q (signal_6286) ) ;
    buf_clk cell_4150 ( .C (CLK), .D (signal_5173), .Q (signal_6294) ) ;
    buf_clk cell_4160 ( .C (CLK), .D (signal_6303), .Q (signal_6304) ) ;
    buf_clk cell_4170 ( .C (CLK), .D (signal_6313), .Q (signal_6314) ) ;
    buf_clk cell_4186 ( .C (CLK), .D (signal_6329), .Q (signal_6330) ) ;
    buf_clk cell_4198 ( .C (CLK), .D (signal_6341), .Q (signal_6342) ) ;
    buf_clk cell_4210 ( .C (CLK), .D (signal_6353), .Q (signal_6354) ) ;
    buf_clk cell_4218 ( .C (CLK), .D (signal_4857), .Q (signal_6362) ) ;
    buf_clk cell_4226 ( .C (CLK), .D (signal_4865), .Q (signal_6370) ) ;
    buf_clk cell_4238 ( .C (CLK), .D (signal_6381), .Q (signal_6382) ) ;
    buf_clk cell_4250 ( .C (CLK), .D (signal_6393), .Q (signal_6394) ) ;
    buf_clk cell_4264 ( .C (CLK), .D (signal_6407), .Q (signal_6408) ) ;
    buf_clk cell_4278 ( .C (CLK), .D (signal_6421), .Q (signal_6422) ) ;
    buf_clk cell_4294 ( .C (CLK), .D (signal_6437), .Q (signal_6438) ) ;
    buf_clk cell_4310 ( .C (CLK), .D (signal_6453), .Q (signal_6454) ) ;
    buf_clk cell_4326 ( .C (CLK), .D (signal_6469), .Q (signal_6470) ) ;
    buf_clk cell_4342 ( .C (CLK), .D (signal_6485), .Q (signal_6486) ) ;
    buf_clk cell_4358 ( .C (CLK), .D (signal_6501), .Q (signal_6502) ) ;
    buf_clk cell_4374 ( .C (CLK), .D (signal_6517), .Q (signal_6518) ) ;
    buf_clk cell_4390 ( .C (CLK), .D (signal_6533), .Q (signal_6534) ) ;
    buf_clk cell_4406 ( .C (CLK), .D (signal_6549), .Q (signal_6550) ) ;
    buf_clk cell_4422 ( .C (CLK), .D (signal_6565), .Q (signal_6566) ) ;
    buf_clk cell_4438 ( .C (CLK), .D (signal_6581), .Q (signal_6582) ) ;
    buf_clk cell_4454 ( .C (CLK), .D (signal_6597), .Q (signal_6598) ) ;
    buf_clk cell_4470 ( .C (CLK), .D (signal_6613), .Q (signal_6614) ) ;
    buf_clk cell_4486 ( .C (CLK), .D (signal_6629), .Q (signal_6630) ) ;
    buf_clk cell_4502 ( .C (CLK), .D (signal_6645), .Q (signal_6646) ) ;
    buf_clk cell_4518 ( .C (CLK), .D (signal_6661), .Q (signal_6662) ) ;
    buf_clk cell_4534 ( .C (CLK), .D (signal_6677), .Q (signal_6678) ) ;
    buf_clk cell_4544 ( .C (CLK), .D (signal_6687), .Q (signal_6688) ) ;
    buf_clk cell_4554 ( .C (CLK), .D (signal_6697), .Q (signal_6698) ) ;
    buf_clk cell_4562 ( .C (CLK), .D (signal_4905), .Q (signal_6706) ) ;
    buf_clk cell_4570 ( .C (CLK), .D (signal_4913), .Q (signal_6714) ) ;
    buf_clk cell_4582 ( .C (CLK), .D (signal_6725), .Q (signal_6726) ) ;
    buf_clk cell_4594 ( .C (CLK), .D (signal_6737), .Q (signal_6738) ) ;
    buf_clk cell_4608 ( .C (CLK), .D (signal_6751), .Q (signal_6752) ) ;
    buf_clk cell_4622 ( .C (CLK), .D (signal_6765), .Q (signal_6766) ) ;
    buf_clk cell_4638 ( .C (CLK), .D (signal_6781), .Q (signal_6782) ) ;
    buf_clk cell_4654 ( .C (CLK), .D (signal_6797), .Q (signal_6798) ) ;
    buf_clk cell_4674 ( .C (CLK), .D (signal_5233), .Q (signal_6818) ) ;
    buf_clk cell_4682 ( .C (CLK), .D (signal_5237), .Q (signal_6826) ) ;
    buf_clk cell_4692 ( .C (CLK), .D (signal_6835), .Q (signal_6836) ) ;
    buf_clk cell_4702 ( .C (CLK), .D (signal_6845), .Q (signal_6846) ) ;
    buf_clk cell_4714 ( .C (CLK), .D (signal_6857), .Q (signal_6858) ) ;
    buf_clk cell_4726 ( .C (CLK), .D (signal_6869), .Q (signal_6870) ) ;
    buf_clk cell_4734 ( .C (CLK), .D (signal_4521), .Q (signal_6878) ) ;
    buf_clk cell_4750 ( .C (CLK), .D (signal_6893), .Q (signal_6894) ) ;
    buf_clk cell_4766 ( .C (CLK), .D (signal_6909), .Q (signal_6910) ) ;
    buf_clk cell_4782 ( .C (CLK), .D (signal_6925), .Q (signal_6926) ) ;
    buf_clk cell_4798 ( .C (CLK), .D (signal_6941), .Q (signal_6942) ) ;
    buf_clk cell_4814 ( .C (CLK), .D (signal_6957), .Q (signal_6958) ) ;
    buf_clk cell_4830 ( .C (CLK), .D (signal_6973), .Q (signal_6974) ) ;
    buf_clk cell_4846 ( .C (CLK), .D (signal_6989), .Q (signal_6990) ) ;
    buf_clk cell_4862 ( .C (CLK), .D (signal_7005), .Q (signal_7006) ) ;
    buf_clk cell_4878 ( .C (CLK), .D (signal_7021), .Q (signal_7022) ) ;
    buf_clk cell_4894 ( .C (CLK), .D (signal_7037), .Q (signal_7038) ) ;
    buf_clk cell_4910 ( .C (CLK), .D (signal_7053), .Q (signal_7054) ) ;
    buf_clk cell_4926 ( .C (CLK), .D (signal_7069), .Q (signal_7070) ) ;
    buf_clk cell_4942 ( .C (CLK), .D (signal_7085), .Q (signal_7086) ) ;
    buf_clk cell_4958 ( .C (CLK), .D (signal_7101), .Q (signal_7102) ) ;
    buf_clk cell_4974 ( .C (CLK), .D (signal_7117), .Q (signal_7118) ) ;
    buf_clk cell_4990 ( .C (CLK), .D (signal_7133), .Q (signal_7134) ) ;
    buf_clk cell_5006 ( .C (CLK), .D (signal_7149), .Q (signal_7150) ) ;
    buf_clk cell_5022 ( .C (CLK), .D (signal_7165), .Q (signal_7166) ) ;
    buf_clk cell_5038 ( .C (CLK), .D (signal_7181), .Q (signal_7182) ) ;
    buf_clk cell_5054 ( .C (CLK), .D (signal_7197), .Q (signal_7198) ) ;
    buf_clk cell_5070 ( .C (CLK), .D (signal_7213), .Q (signal_7214) ) ;
    buf_clk cell_5086 ( .C (CLK), .D (signal_7229), .Q (signal_7230) ) ;
    buf_clk cell_5102 ( .C (CLK), .D (signal_7245), .Q (signal_7246) ) ;
    buf_clk cell_5118 ( .C (CLK), .D (signal_7261), .Q (signal_7262) ) ;
    buf_clk cell_5134 ( .C (CLK), .D (signal_7277), .Q (signal_7278) ) ;
    buf_clk cell_5150 ( .C (CLK), .D (signal_7293), .Q (signal_7294) ) ;
    buf_clk cell_5166 ( .C (CLK), .D (signal_7309), .Q (signal_7310) ) ;
    buf_clk cell_5182 ( .C (CLK), .D (signal_7325), .Q (signal_7326) ) ;
    buf_clk cell_5198 ( .C (CLK), .D (signal_7341), .Q (signal_7342) ) ;
    buf_clk cell_5214 ( .C (CLK), .D (signal_7357), .Q (signal_7358) ) ;
    buf_clk cell_5230 ( .C (CLK), .D (signal_7373), .Q (signal_7374) ) ;
    buf_clk cell_5246 ( .C (CLK), .D (signal_7389), .Q (signal_7390) ) ;
    buf_clk cell_5262 ( .C (CLK), .D (signal_7405), .Q (signal_7406) ) ;
    buf_clk cell_5278 ( .C (CLK), .D (signal_7421), .Q (signal_7422) ) ;
    buf_clk cell_5294 ( .C (CLK), .D (signal_7437), .Q (signal_7438) ) ;
    buf_clk cell_5310 ( .C (CLK), .D (signal_7453), .Q (signal_7454) ) ;
    buf_clk cell_5326 ( .C (CLK), .D (signal_7469), .Q (signal_7470) ) ;
    buf_clk cell_5342 ( .C (CLK), .D (signal_7485), .Q (signal_7486) ) ;
    buf_clk cell_5358 ( .C (CLK), .D (signal_7501), .Q (signal_7502) ) ;
    buf_clk cell_5374 ( .C (CLK), .D (signal_7517), .Q (signal_7518) ) ;
    buf_clk cell_5390 ( .C (CLK), .D (signal_7533), .Q (signal_7534) ) ;
    buf_clk cell_5406 ( .C (CLK), .D (signal_7549), .Q (signal_7550) ) ;
    buf_clk cell_5422 ( .C (CLK), .D (signal_7565), .Q (signal_7566) ) ;
    buf_clk cell_5438 ( .C (CLK), .D (signal_7581), .Q (signal_7582) ) ;
    buf_clk cell_5454 ( .C (CLK), .D (signal_7597), .Q (signal_7598) ) ;
    buf_clk cell_5470 ( .C (CLK), .D (signal_7613), .Q (signal_7614) ) ;
    buf_clk cell_5486 ( .C (CLK), .D (signal_7629), .Q (signal_7630) ) ;
    buf_clk cell_5502 ( .C (CLK), .D (signal_7645), .Q (signal_7646) ) ;
    buf_clk cell_5518 ( .C (CLK), .D (signal_7661), .Q (signal_7662) ) ;
    buf_clk cell_5534 ( .C (CLK), .D (signal_7677), .Q (signal_7678) ) ;
    buf_clk cell_5550 ( .C (CLK), .D (signal_7693), .Q (signal_7694) ) ;
    buf_clk cell_5566 ( .C (CLK), .D (signal_7709), .Q (signal_7710) ) ;
    buf_clk cell_5582 ( .C (CLK), .D (signal_7725), .Q (signal_7726) ) ;
    buf_clk cell_5598 ( .C (CLK), .D (signal_7741), .Q (signal_7742) ) ;
    buf_clk cell_5614 ( .C (CLK), .D (signal_7757), .Q (signal_7758) ) ;
    buf_clk cell_5630 ( .C (CLK), .D (signal_7773), .Q (signal_7774) ) ;
    buf_clk cell_5646 ( .C (CLK), .D (signal_7789), .Q (signal_7790) ) ;
    buf_clk cell_5662 ( .C (CLK), .D (signal_7805), .Q (signal_7806) ) ;
    buf_clk cell_5678 ( .C (CLK), .D (signal_7821), .Q (signal_7822) ) ;
    buf_clk cell_5694 ( .C (CLK), .D (signal_7837), .Q (signal_7838) ) ;
    buf_clk cell_5710 ( .C (CLK), .D (signal_7853), .Q (signal_7854) ) ;
    buf_clk cell_5726 ( .C (CLK), .D (signal_7869), .Q (signal_7870) ) ;
    buf_clk cell_5742 ( .C (CLK), .D (signal_7885), .Q (signal_7886) ) ;
    buf_clk cell_5758 ( .C (CLK), .D (signal_7901), .Q (signal_7902) ) ;
    buf_clk cell_5774 ( .C (CLK), .D (signal_7917), .Q (signal_7918) ) ;
    buf_clk cell_5790 ( .C (CLK), .D (signal_7933), .Q (signal_7934) ) ;
    buf_clk cell_5806 ( .C (CLK), .D (signal_7949), .Q (signal_7950) ) ;
    buf_clk cell_5822 ( .C (CLK), .D (signal_7965), .Q (signal_7966) ) ;
    buf_clk cell_5838 ( .C (CLK), .D (signal_7981), .Q (signal_7982) ) ;
    buf_clk cell_5854 ( .C (CLK), .D (signal_7997), .Q (signal_7998) ) ;
    buf_clk cell_5870 ( .C (CLK), .D (signal_8013), .Q (signal_8014) ) ;
    buf_clk cell_5886 ( .C (CLK), .D (signal_8029), .Q (signal_8030) ) ;
    buf_clk cell_5902 ( .C (CLK), .D (signal_8045), .Q (signal_8046) ) ;
    buf_clk cell_5918 ( .C (CLK), .D (signal_8061), .Q (signal_8062) ) ;
    buf_clk cell_5934 ( .C (CLK), .D (signal_8077), .Q (signal_8078) ) ;
    buf_clk cell_5950 ( .C (CLK), .D (signal_8093), .Q (signal_8094) ) ;
    buf_clk cell_5966 ( .C (CLK), .D (signal_8109), .Q (signal_8110) ) ;
    buf_clk cell_5982 ( .C (CLK), .D (signal_8125), .Q (signal_8126) ) ;
    buf_clk cell_5998 ( .C (CLK), .D (signal_8141), .Q (signal_8142) ) ;
    buf_clk cell_6014 ( .C (CLK), .D (signal_8157), .Q (signal_8158) ) ;
    buf_clk cell_6030 ( .C (CLK), .D (signal_8173), .Q (signal_8174) ) ;
    buf_clk cell_6046 ( .C (CLK), .D (signal_8189), .Q (signal_8190) ) ;
    buf_clk cell_6062 ( .C (CLK), .D (signal_8205), .Q (signal_8206) ) ;
    buf_clk cell_6078 ( .C (CLK), .D (signal_8221), .Q (signal_8222) ) ;
    buf_clk cell_6094 ( .C (CLK), .D (signal_8237), .Q (signal_8238) ) ;
    buf_clk cell_6110 ( .C (CLK), .D (signal_8253), .Q (signal_8254) ) ;
    buf_clk cell_6126 ( .C (CLK), .D (signal_8269), .Q (signal_8270) ) ;
    buf_clk cell_6142 ( .C (CLK), .D (signal_8285), .Q (signal_8286) ) ;
    buf_clk cell_6158 ( .C (CLK), .D (signal_8301), .Q (signal_8302) ) ;
    buf_clk cell_6174 ( .C (CLK), .D (signal_8317), .Q (signal_8318) ) ;
    buf_clk cell_6190 ( .C (CLK), .D (signal_8333), .Q (signal_8334) ) ;
    buf_clk cell_6206 ( .C (CLK), .D (signal_8349), .Q (signal_8350) ) ;
    buf_clk cell_6222 ( .C (CLK), .D (signal_8365), .Q (signal_8366) ) ;
    buf_clk cell_6238 ( .C (CLK), .D (signal_8381), .Q (signal_8382) ) ;
    buf_clk cell_6254 ( .C (CLK), .D (signal_8397), .Q (signal_8398) ) ;
    buf_clk cell_6270 ( .C (CLK), .D (signal_8413), .Q (signal_8414) ) ;
    buf_clk cell_6286 ( .C (CLK), .D (signal_8429), .Q (signal_8430) ) ;
    buf_clk cell_6302 ( .C (CLK), .D (signal_8445), .Q (signal_8446) ) ;
    buf_clk cell_6318 ( .C (CLK), .D (signal_8461), .Q (signal_8462) ) ;
    buf_clk cell_6334 ( .C (CLK), .D (signal_8477), .Q (signal_8478) ) ;
    buf_clk cell_6350 ( .C (CLK), .D (signal_8493), .Q (signal_8494) ) ;
    buf_clk cell_6366 ( .C (CLK), .D (signal_8509), .Q (signal_8510) ) ;
    buf_clk cell_6382 ( .C (CLK), .D (signal_8525), .Q (signal_8526) ) ;
    buf_clk cell_6398 ( .C (CLK), .D (signal_8541), .Q (signal_8542) ) ;
    buf_clk cell_6406 ( .C (CLK), .D (signal_657), .Q (signal_8550) ) ;
    buf_clk cell_6414 ( .C (CLK), .D (signal_2958), .Q (signal_8558) ) ;
    buf_clk cell_6422 ( .C (CLK), .D (signal_1309), .Q (signal_8566) ) ;
    buf_clk cell_6430 ( .C (CLK), .D (signal_3041), .Q (signal_8574) ) ;
    buf_clk cell_6438 ( .C (CLK), .D (signal_658), .Q (signal_8582) ) ;
    buf_clk cell_6446 ( .C (CLK), .D (signal_2920), .Q (signal_8590) ) ;
    buf_clk cell_6454 ( .C (CLK), .D (signal_665), .Q (signal_8598) ) ;
    buf_clk cell_6462 ( .C (CLK), .D (signal_3001), .Q (signal_8606) ) ;
    buf_clk cell_6470 ( .C (CLK), .D (signal_668), .Q (signal_8614) ) ;
    buf_clk cell_6478 ( .C (CLK), .D (signal_2959), .Q (signal_8622) ) ;
    buf_clk cell_6486 ( .C (CLK), .D (signal_883), .Q (signal_8630) ) ;
    buf_clk cell_6494 ( .C (CLK), .D (signal_2610), .Q (signal_8638) ) ;
    buf_clk cell_6502 ( .C (CLK), .D (signal_881), .Q (signal_8646) ) ;
    buf_clk cell_6510 ( .C (CLK), .D (signal_2609), .Q (signal_8654) ) ;
    buf_clk cell_6518 ( .C (CLK), .D (signal_671), .Q (signal_8662) ) ;
    buf_clk cell_6526 ( .C (CLK), .D (signal_2742), .Q (signal_8670) ) ;
    buf_clk cell_6534 ( .C (CLK), .D (signal_681), .Q (signal_8678) ) ;
    buf_clk cell_6542 ( .C (CLK), .D (signal_2744), .Q (signal_8686) ) ;
    buf_clk cell_6550 ( .C (CLK), .D (signal_882), .Q (signal_8694) ) ;
    buf_clk cell_6558 ( .C (CLK), .D (signal_2622), .Q (signal_8702) ) ;
    buf_clk cell_6566 ( .C (CLK), .D (signal_684), .Q (signal_8710) ) ;
    buf_clk cell_6574 ( .C (CLK), .D (signal_2961), .Q (signal_8718) ) ;
    buf_clk cell_6582 ( .C (CLK), .D (signal_686), .Q (signal_8726) ) ;
    buf_clk cell_6590 ( .C (CLK), .D (signal_2745), .Q (signal_8734) ) ;
    buf_clk cell_6598 ( .C (CLK), .D (signal_922), .Q (signal_8742) ) ;
    buf_clk cell_6606 ( .C (CLK), .D (signal_2653), .Q (signal_8750) ) ;
    buf_clk cell_6614 ( .C (CLK), .D (signal_940), .Q (signal_8758) ) ;
    buf_clk cell_6622 ( .C (CLK), .D (signal_2734), .Q (signal_8766) ) ;
    buf_clk cell_6630 ( .C (CLK), .D (signal_677), .Q (signal_8774) ) ;
    buf_clk cell_6638 ( .C (CLK), .D (signal_2746), .Q (signal_8782) ) ;
    buf_clk cell_6646 ( .C (CLK), .D (signal_1324), .Q (signal_8790) ) ;
    buf_clk cell_6654 ( .C (CLK), .D (signal_2922), .Q (signal_8798) ) ;
    buf_clk cell_6662 ( .C (CLK), .D (signal_920), .Q (signal_8806) ) ;
    buf_clk cell_6670 ( .C (CLK), .D (signal_2737), .Q (signal_8814) ) ;
    buf_clk cell_6678 ( .C (CLK), .D (signal_692), .Q (signal_8822) ) ;
    buf_clk cell_6686 ( .C (CLK), .D (signal_2747), .Q (signal_8830) ) ;
    buf_clk cell_6694 ( .C (CLK), .D (signal_695), .Q (signal_8838) ) ;
    buf_clk cell_6702 ( .C (CLK), .D (signal_2923), .Q (signal_8846) ) ;
    buf_clk cell_6710 ( .C (CLK), .D (signal_1305), .Q (signal_8854) ) ;
    buf_clk cell_6718 ( .C (CLK), .D (signal_3045), .Q (signal_8862) ) ;
    buf_clk cell_6726 ( .C (CLK), .D (signal_696), .Q (signal_8870) ) ;
    buf_clk cell_6734 ( .C (CLK), .D (signal_2924), .Q (signal_8878) ) ;
    buf_clk cell_6742 ( .C (CLK), .D (signal_703), .Q (signal_8886) ) ;
    buf_clk cell_6750 ( .C (CLK), .D (signal_3006), .Q (signal_8894) ) ;
    buf_clk cell_6758 ( .C (CLK), .D (signal_706), .Q (signal_8902) ) ;
    buf_clk cell_6766 ( .C (CLK), .D (signal_2925), .Q (signal_8910) ) ;
    buf_clk cell_6774 ( .C (CLK), .D (signal_895), .Q (signal_8918) ) ;
    buf_clk cell_6782 ( .C (CLK), .D (signal_2672), .Q (signal_8926) ) ;
    buf_clk cell_6790 ( .C (CLK), .D (signal_893), .Q (signal_8934) ) ;
    buf_clk cell_6798 ( .C (CLK), .D (signal_2649), .Q (signal_8942) ) ;
    buf_clk cell_6806 ( .C (CLK), .D (signal_709), .Q (signal_8950) ) ;
    buf_clk cell_6814 ( .C (CLK), .D (signal_2817), .Q (signal_8958) ) ;
    buf_clk cell_6822 ( .C (CLK), .D (signal_719), .Q (signal_8966) ) ;
    buf_clk cell_6830 ( .C (CLK), .D (signal_2749), .Q (signal_8974) ) ;
    buf_clk cell_6838 ( .C (CLK), .D (signal_894), .Q (signal_8982) ) ;
    buf_clk cell_6846 ( .C (CLK), .D (signal_2671), .Q (signal_8990) ) ;
    buf_clk cell_6854 ( .C (CLK), .D (signal_722), .Q (signal_8998) ) ;
    buf_clk cell_6862 ( .C (CLK), .D (signal_2927), .Q (signal_9006) ) ;
    buf_clk cell_6870 ( .C (CLK), .D (signal_724), .Q (signal_9014) ) ;
    buf_clk cell_6878 ( .C (CLK), .D (signal_2750), .Q (signal_9022) ) ;
    buf_clk cell_6886 ( .C (CLK), .D (signal_918), .Q (signal_9030) ) ;
    buf_clk cell_6894 ( .C (CLK), .D (signal_2617), .Q (signal_9038) ) ;
    buf_clk cell_6902 ( .C (CLK), .D (signal_936), .Q (signal_9046) ) ;
    buf_clk cell_6910 ( .C (CLK), .D (signal_2735), .Q (signal_9054) ) ;
    buf_clk cell_6918 ( .C (CLK), .D (signal_715), .Q (signal_9062) ) ;
    buf_clk cell_6926 ( .C (CLK), .D (signal_2820), .Q (signal_9070) ) ;
    buf_clk cell_6934 ( .C (CLK), .D (signal_1320), .Q (signal_9078) ) ;
    buf_clk cell_6942 ( .C (CLK), .D (signal_2882), .Q (signal_9086) ) ;
    buf_clk cell_6950 ( .C (CLK), .D (signal_916), .Q (signal_9094) ) ;
    buf_clk cell_6958 ( .C (CLK), .D (signal_2635), .Q (signal_9102) ) ;
    buf_clk cell_6966 ( .C (CLK), .D (signal_730), .Q (signal_9110) ) ;
    buf_clk cell_6974 ( .C (CLK), .D (signal_2821), .Q (signal_9118) ) ;
    buf_clk cell_6982 ( .C (CLK), .D (signal_733), .Q (signal_9126) ) ;
    buf_clk cell_6990 ( .C (CLK), .D (signal_2930), .Q (signal_9134) ) ;
    buf_clk cell_6998 ( .C (CLK), .D (signal_1301), .Q (signal_9142) ) ;
    buf_clk cell_7006 ( .C (CLK), .D (signal_3010), .Q (signal_9150) ) ;
    buf_clk cell_7014 ( .C (CLK), .D (signal_734), .Q (signal_9158) ) ;
    buf_clk cell_7022 ( .C (CLK), .D (signal_2883), .Q (signal_9166) ) ;
    buf_clk cell_7030 ( .C (CLK), .D (signal_741), .Q (signal_9174) ) ;
    buf_clk cell_7038 ( .C (CLK), .D (signal_2969), .Q (signal_9182) ) ;
    buf_clk cell_7046 ( .C (CLK), .D (signal_744), .Q (signal_9190) ) ;
    buf_clk cell_7054 ( .C (CLK), .D (signal_2931), .Q (signal_9198) ) ;
    buf_clk cell_7062 ( .C (CLK), .D (signal_891), .Q (signal_9206) ) ;
    buf_clk cell_7070 ( .C (CLK), .D (signal_2679), .Q (signal_9214) ) ;
    buf_clk cell_7078 ( .C (CLK), .D (signal_889), .Q (signal_9222) ) ;
    buf_clk cell_7086 ( .C (CLK), .D (signal_2677), .Q (signal_9230) ) ;
    buf_clk cell_7094 ( .C (CLK), .D (signal_747), .Q (signal_9238) ) ;
    buf_clk cell_7102 ( .C (CLK), .D (signal_2823), .Q (signal_9246) ) ;
    buf_clk cell_7110 ( .C (CLK), .D (signal_757), .Q (signal_9254) ) ;
    buf_clk cell_7118 ( .C (CLK), .D (signal_2827), .Q (signal_9262) ) ;
    buf_clk cell_7126 ( .C (CLK), .D (signal_890), .Q (signal_9270) ) ;
    buf_clk cell_7134 ( .C (CLK), .D (signal_2675), .Q (signal_9278) ) ;
    buf_clk cell_7142 ( .C (CLK), .D (signal_760), .Q (signal_9286) ) ;
    buf_clk cell_7150 ( .C (CLK), .D (signal_2933), .Q (signal_9294) ) ;
    buf_clk cell_7158 ( .C (CLK), .D (signal_762), .Q (signal_9302) ) ;
    buf_clk cell_7166 ( .C (CLK), .D (signal_2828), .Q (signal_9310) ) ;
    buf_clk cell_7174 ( .C (CLK), .D (signal_914), .Q (signal_9318) ) ;
    buf_clk cell_7182 ( .C (CLK), .D (signal_2615), .Q (signal_9326) ) ;
    buf_clk cell_7190 ( .C (CLK), .D (signal_932), .Q (signal_9334) ) ;
    buf_clk cell_7198 ( .C (CLK), .D (signal_2633), .Q (signal_9342) ) ;
    buf_clk cell_7206 ( .C (CLK), .D (signal_753), .Q (signal_9350) ) ;
    buf_clk cell_7214 ( .C (CLK), .D (signal_2829), .Q (signal_9358) ) ;
    buf_clk cell_7222 ( .C (CLK), .D (signal_1316), .Q (signal_9366) ) ;
    buf_clk cell_7230 ( .C (CLK), .D (signal_2885), .Q (signal_9374) ) ;
    buf_clk cell_7238 ( .C (CLK), .D (signal_912), .Q (signal_9382) ) ;
    buf_clk cell_7246 ( .C (CLK), .D (signal_2636), .Q (signal_9390) ) ;
    buf_clk cell_7254 ( .C (CLK), .D (signal_768), .Q (signal_9398) ) ;
    buf_clk cell_7262 ( .C (CLK), .D (signal_2830), .Q (signal_9406) ) ;
    buf_clk cell_7270 ( .C (CLK), .D (signal_771), .Q (signal_9414) ) ;
    buf_clk cell_7278 ( .C (CLK), .D (signal_2975), .Q (signal_9422) ) ;
    buf_clk cell_7286 ( .C (CLK), .D (signal_1297), .Q (signal_9430) ) ;
    buf_clk cell_7294 ( .C (CLK), .D (signal_3014), .Q (signal_9438) ) ;
    buf_clk cell_7302 ( .C (CLK), .D (signal_772), .Q (signal_9446) ) ;
    buf_clk cell_7310 ( .C (CLK), .D (signal_2886), .Q (signal_9454) ) ;
    buf_clk cell_7318 ( .C (CLK), .D (signal_779), .Q (signal_9462) ) ;
    buf_clk cell_7326 ( .C (CLK), .D (signal_2976), .Q (signal_9470) ) ;
    buf_clk cell_7334 ( .C (CLK), .D (signal_782), .Q (signal_9478) ) ;
    buf_clk cell_7342 ( .C (CLK), .D (signal_2977), .Q (signal_9486) ) ;
    buf_clk cell_7350 ( .C (CLK), .D (signal_887), .Q (signal_9494) ) ;
    buf_clk cell_7358 ( .C (CLK), .D (signal_2616), .Q (signal_9502) ) ;
    buf_clk cell_7366 ( .C (CLK), .D (signal_885), .Q (signal_9510) ) ;
    buf_clk cell_7374 ( .C (CLK), .D (signal_2621), .Q (signal_9518) ) ;
    buf_clk cell_7382 ( .C (CLK), .D (signal_785), .Q (signal_9526) ) ;
    buf_clk cell_7390 ( .C (CLK), .D (signal_2754), .Q (signal_9534) ) ;
    buf_clk cell_7398 ( .C (CLK), .D (signal_795), .Q (signal_9542) ) ;
    buf_clk cell_7406 ( .C (CLK), .D (signal_2834), .Q (signal_9550) ) ;
    buf_clk cell_7414 ( .C (CLK), .D (signal_886), .Q (signal_9558) ) ;
    buf_clk cell_7422 ( .C (CLK), .D (signal_2627), .Q (signal_9566) ) ;
    buf_clk cell_7430 ( .C (CLK), .D (signal_798), .Q (signal_9574) ) ;
    buf_clk cell_7438 ( .C (CLK), .D (signal_2979), .Q (signal_9582) ) ;
    buf_clk cell_7446 ( .C (CLK), .D (signal_800), .Q (signal_9590) ) ;
    buf_clk cell_7454 ( .C (CLK), .D (signal_2835), .Q (signal_9598) ) ;
    buf_clk cell_7462 ( .C (CLK), .D (signal_926), .Q (signal_9606) ) ;
    buf_clk cell_7470 ( .C (CLK), .D (signal_2652), .Q (signal_9614) ) ;
    buf_clk cell_7478 ( .C (CLK), .D (signal_928), .Q (signal_9622) ) ;
    buf_clk cell_7486 ( .C (CLK), .D (signal_2634), .Q (signal_9630) ) ;
    buf_clk cell_7494 ( .C (CLK), .D (signal_791), .Q (signal_9638) ) ;
    buf_clk cell_7502 ( .C (CLK), .D (signal_2756), .Q (signal_9646) ) ;
    buf_clk cell_7510 ( .C (CLK), .D (signal_1312), .Q (signal_9654) ) ;
    buf_clk cell_7518 ( .C (CLK), .D (signal_2936), .Q (signal_9662) ) ;
    buf_clk cell_7526 ( .C (CLK), .D (signal_924), .Q (signal_9670) ) ;
    buf_clk cell_7534 ( .C (CLK), .D (signal_2736), .Q (signal_9678) ) ;
    buf_clk cell_7542 ( .C (CLK), .D (signal_806), .Q (signal_9686) ) ;
    buf_clk cell_7550 ( .C (CLK), .D (signal_2836), .Q (signal_9694) ) ;
    buf_clk cell_7564 ( .C (CLK), .D (signal_9707), .Q (signal_9708) ) ;
    buf_clk cell_7572 ( .C (CLK), .D (signal_9715), .Q (signal_9716) ) ;
    buf_clk cell_7598 ( .C (CLK), .D (signal_9741), .Q (signal_9742) ) ;
    buf_clk cell_7614 ( .C (CLK), .D (signal_9757), .Q (signal_9758) ) ;
    buf_clk cell_7630 ( .C (CLK), .D (signal_9773), .Q (signal_9774) ) ;
    buf_clk cell_7646 ( .C (CLK), .D (signal_9789), .Q (signal_9790) ) ;
    buf_clk cell_7662 ( .C (CLK), .D (signal_9805), .Q (signal_9806) ) ;
    buf_clk cell_7678 ( .C (CLK), .D (signal_9821), .Q (signal_9822) ) ;
    buf_clk cell_7694 ( .C (CLK), .D (signal_9837), .Q (signal_9838) ) ;
    buf_clk cell_7710 ( .C (CLK), .D (signal_9853), .Q (signal_9854) ) ;
    buf_clk cell_7726 ( .C (CLK), .D (signal_9869), .Q (signal_9870) ) ;
    buf_clk cell_7742 ( .C (CLK), .D (signal_9885), .Q (signal_9886) ) ;
    buf_clk cell_7750 ( .C (CLK), .D (signal_1198), .Q (signal_9894) ) ;
    buf_clk cell_7758 ( .C (CLK), .D (signal_3028), .Q (signal_9902) ) ;
    buf_clk cell_7766 ( .C (CLK), .D (signal_1196), .Q (signal_9910) ) ;
    buf_clk cell_7774 ( .C (CLK), .D (signal_2992), .Q (signal_9918) ) ;
    buf_clk cell_7782 ( .C (CLK), .D (signal_1194), .Q (signal_9926) ) ;
    buf_clk cell_7790 ( .C (CLK), .D (signal_3032), .Q (signal_9934) ) ;
    buf_clk cell_7798 ( .C (CLK), .D (signal_1192), .Q (signal_9942) ) ;
    buf_clk cell_7806 ( .C (CLK), .D (signal_2955), .Q (signal_9950) ) ;
    buf_clk cell_7814 ( .C (CLK), .D (signal_1190), .Q (signal_9958) ) ;
    buf_clk cell_7822 ( .C (CLK), .D (signal_2996), .Q (signal_9966) ) ;
    buf_clk cell_7830 ( .C (CLK), .D (signal_1188), .Q (signal_9974) ) ;
    buf_clk cell_7838 ( .C (CLK), .D (signal_2957), .Q (signal_9982) ) ;
    buf_clk cell_7846 ( .C (CLK), .D (signal_1186), .Q (signal_9990) ) ;
    buf_clk cell_7854 ( .C (CLK), .D (signal_2998), .Q (signal_9998) ) ;
    buf_clk cell_7862 ( .C (CLK), .D (signal_1184), .Q (signal_10006) ) ;
    buf_clk cell_7870 ( .C (CLK), .D (signal_3000), .Q (signal_10014) ) ;
    buf_clk cell_7878 ( .C (CLK), .D (signal_1181), .Q (signal_10022) ) ;
    buf_clk cell_7886 ( .C (CLK), .D (signal_3112), .Q (signal_10030) ) ;
    buf_clk cell_7894 ( .C (CLK), .D (signal_1177), .Q (signal_10038) ) ;
    buf_clk cell_7902 ( .C (CLK), .D (signal_3114), .Q (signal_10046) ) ;
    buf_clk cell_7910 ( .C (CLK), .D (signal_1173), .Q (signal_10054) ) ;
    buf_clk cell_7918 ( .C (CLK), .D (signal_3073), .Q (signal_10062) ) ;
    buf_clk cell_7926 ( .C (CLK), .D (signal_1169), .Q (signal_10070) ) ;
    buf_clk cell_7934 ( .C (CLK), .D (signal_3077), .Q (signal_10078) ) ;
    buf_clk cell_7950 ( .C (CLK), .D (signal_10093), .Q (signal_10094) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1576 ( .s ({signal_5157, signal_5155}), .b ({signal_2614, signal_1660}), .a ({signal_2613, signal_898}), .clk (CLK), .r (Fresh[448]), .c ({signal_2722, signal_1720}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1577 ( .s ({signal_5157, signal_5155}), .b ({signal_2613, signal_898}), .a ({signal_2614, signal_1660}), .clk (CLK), .r (Fresh[449]), .c ({signal_2723, signal_1721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1578 ( .s ({signal_5169, signal_5163}), .b ({signal_2614, signal_1660}), .a ({signal_2613, signal_898}), .clk (CLK), .r (Fresh[450]), .c ({signal_2724, signal_1722}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1579 ( .s ({signal_4849, signal_4841}), .b ({signal_2655, signal_1662}), .a ({signal_2654, signal_1661}), .clk (CLK), .r (Fresh[451]), .c ({signal_2757, signal_1723}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1580 ( .s ({signal_5173, signal_5171}), .b ({signal_5177, signal_5175}), .a ({signal_2656, signal_1663}), .clk (CLK), .r (Fresh[452]), .c ({signal_2758, signal_1724}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1581 ( .s ({signal_5173, signal_5171}), .b ({signal_2658, signal_1665}), .a ({signal_2657, signal_1664}), .clk (CLK), .r (Fresh[453]), .c ({signal_2759, signal_1725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1582 ( .s ({signal_5173, signal_5171}), .b ({signal_5181, signal_5179}), .a ({signal_2659, signal_1666}), .clk (CLK), .r (Fresh[454]), .c ({signal_2760, signal_1726}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1583 ( .s ({signal_5173, signal_5171}), .b ({signal_2661, signal_1668}), .a ({signal_2660, signal_1667}), .clk (CLK), .r (Fresh[455]), .c ({signal_2761, signal_1727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1584 ( .s ({signal_5173, signal_5171}), .b ({signal_5185, signal_5183}), .a ({signal_2662, signal_1669}), .clk (CLK), .r (Fresh[456]), .c ({signal_2762, signal_1728}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1585 ( .s ({signal_5173, signal_5171}), .b ({signal_2664, signal_1671}), .a ({signal_2663, signal_1670}), .clk (CLK), .r (Fresh[457]), .c ({signal_2763, signal_1729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1586 ( .s ({signal_5189, signal_5187}), .b ({signal_2667, signal_1674}), .a ({signal_2666, signal_1673}), .clk (CLK), .r (Fresh[458]), .c ({signal_2764, signal_1730}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1587 ( .s ({signal_4721, signal_4717}), .b ({signal_2668, signal_1675}), .a ({signal_5193, signal_5191}), .clk (CLK), .r (Fresh[459]), .c ({signal_2765, signal_1731}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1588 ( .s ({signal_5189, signal_5187}), .b ({signal_2666, signal_1673}), .a ({signal_2667, signal_1674}), .clk (CLK), .r (Fresh[460]), .c ({signal_2766, signal_1732}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1589 ( .s ({signal_4721, signal_4717}), .b ({signal_5197, signal_5195}), .a ({signal_2670, signal_1677}), .clk (CLK), .r (Fresh[461]), .c ({signal_2767, signal_1733}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1590 ( .s ({signal_5213, signal_5205}), .b ({signal_2678, signal_1678}), .a ({signal_2674, signal_910}), .clk (CLK), .r (Fresh[462]), .c ({signal_2768, signal_1734}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1591 ( .s ({signal_5213, signal_5205}), .b ({signal_2674, signal_910}), .a ({signal_2678, signal_1678}), .clk (CLK), .r (Fresh[463]), .c ({signal_2769, signal_1735}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1592 ( .s ({signal_4513, signal_4507}), .b ({signal_2678, signal_1678}), .a ({signal_2674, signal_910}), .clk (CLK), .r (Fresh[464]), .c ({signal_2770, signal_1736}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1593 ( .s ({signal_4833, signal_4829}), .b ({signal_5217, signal_5215}), .a ({signal_2683, signal_1680}), .clk (CLK), .r (Fresh[465]), .c ({signal_2771, signal_1737}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1594 ( .s ({signal_4833, signal_4829}), .b ({signal_5221, signal_5219}), .a ({signal_2684, signal_1681}), .clk (CLK), .r (Fresh[466]), .c ({signal_2772, signal_1738}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1595 ( .s ({signal_4833, signal_4829}), .b ({signal_5225, signal_5223}), .a ({signal_2684, signal_1681}), .clk (CLK), .r (Fresh[467]), .c ({signal_2773, signal_1739}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1596 ( .s ({signal_4833, signal_4829}), .b ({signal_5229, signal_5227}), .a ({signal_2683, signal_1680}), .clk (CLK), .r (Fresh[468]), .c ({signal_2774, signal_1740}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1597 ( .s ({signal_5237, signal_5233}), .b ({signal_5241, signal_5239}), .a ({signal_2689, signal_1685}), .clk (CLK), .r (Fresh[469]), .c ({signal_2775, signal_1741}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1598 ( .s ({signal_5237, signal_5233}), .b ({signal_2691, signal_1687}), .a ({signal_2690, signal_1686}), .clk (CLK), .r (Fresh[470]), .c ({signal_2776, signal_1742}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1599 ( .s ({signal_5237, signal_5233}), .b ({signal_5245, signal_5243}), .a ({signal_2692, signal_1688}), .clk (CLK), .r (Fresh[471]), .c ({signal_2777, signal_1743}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1600 ( .s ({signal_5237, signal_5233}), .b ({signal_2694, signal_1690}), .a ({signal_2693, signal_1689}), .clk (CLK), .r (Fresh[472]), .c ({signal_2778, signal_1744}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1601 ( .s ({signal_5249, signal_5247}), .b ({signal_2698, signal_1692}), .a ({signal_2697, signal_1691}), .clk (CLK), .r (Fresh[473]), .c ({signal_2779, signal_1745}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1602 ( .s ({signal_5249, signal_5247}), .b ({signal_2700, signal_1694}), .a ({signal_2699, signal_1693}), .clk (CLK), .r (Fresh[474]), .c ({signal_2780, signal_1746}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1603 ( .s ({signal_5169, signal_5163}), .b ({signal_2702, signal_1696}), .a ({signal_2701, signal_1695}), .clk (CLK), .r (Fresh[475]), .c ({signal_2781, signal_1747}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1604 ( .s ({signal_5169, signal_5163}), .b ({signal_2704, signal_1698}), .a ({signal_2703, signal_1697}), .clk (CLK), .r (Fresh[476]), .c ({signal_2782, signal_1748}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1605 ( .s ({signal_4413, signal_4405}), .b ({signal_2703, signal_1697}), .a ({signal_2701, signal_1695}), .clk (CLK), .r (Fresh[477]), .c ({signal_2783, signal_1749}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1606 ( .s ({signal_5169, signal_5163}), .b ({signal_2701, signal_1695}), .a ({signal_2702, signal_1696}), .clk (CLK), .r (Fresh[478]), .c ({signal_2784, signal_1750}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1607 ( .s ({signal_5169, signal_5163}), .b ({signal_2703, signal_1697}), .a ({signal_2704, signal_1698}), .clk (CLK), .r (Fresh[479]), .c ({signal_2785, signal_1751}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1608 ( .s ({signal_4413, signal_4405}), .b ({signal_2704, signal_1698}), .a ({signal_2702, signal_1696}), .clk (CLK), .r (Fresh[480]), .c ({signal_2786, signal_1752}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1609 ( .s ({signal_4437, signal_4429}), .b ({signal_2705, signal_1699}), .a ({signal_2675, signal_890}), .clk (CLK), .r (Fresh[481]), .c ({signal_2787, signal_1753}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1610 ( .s ({signal_4437, signal_4429}), .b ({signal_2675, signal_890}), .a ({signal_2705, signal_1699}), .clk (CLK), .r (Fresh[482]), .c ({signal_2788, signal_1754}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1611 ( .s ({signal_5253, signal_5251}), .b ({signal_5257, signal_5255}), .a ({signal_2623, signal_1700}), .clk (CLK), .r (Fresh[483]), .c ({signal_2725, signal_1755}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1612 ( .s ({signal_5253, signal_5251}), .b ({signal_5261, signal_5259}), .a ({signal_2624, signal_1701}), .clk (CLK), .r (Fresh[484]), .c ({signal_2726, signal_1756}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1613 ( .s ({signal_5253, signal_5251}), .b ({signal_2623, signal_1700}), .a ({signal_2624, signal_1701}), .clk (CLK), .r (Fresh[485]), .c ({signal_2727, signal_1757}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1614 ( .s ({signal_5253, signal_5251}), .b ({signal_2624, signal_1701}), .a ({signal_2623, signal_1700}), .clk (CLK), .r (Fresh[486]), .c ({signal_2728, signal_1758}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1615 ( .s ({signal_4453, signal_4449}), .b ({signal_2628, signal_1704}), .a ({signal_2627, signal_886}), .clk (CLK), .r (Fresh[487]), .c ({signal_2729, signal_1759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1616 ( .s ({signal_4453, signal_4449}), .b ({signal_2627, signal_886}), .a ({signal_2628, signal_1704}), .clk (CLK), .r (Fresh[488]), .c ({signal_2730, signal_1760}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1617 ( .s ({signal_4445, signal_4441}), .b ({signal_2707, signal_1706}), .a ({signal_2706, signal_1705}), .clk (CLK), .r (Fresh[489]), .c ({signal_2789, signal_1761}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1618 ( .s ({signal_4445, signal_4441}), .b ({signal_2708, signal_1707}), .a ({signal_5265, signal_5263}), .clk (CLK), .r (Fresh[490]), .c ({signal_2790, signal_1762}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1619 ( .s ({signal_4445, signal_4441}), .b ({signal_2706, signal_1705}), .a ({signal_2707, signal_1706}), .clk (CLK), .r (Fresh[491]), .c ({signal_2791, signal_1763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1620 ( .s ({signal_4445, signal_4441}), .b ({signal_2709, signal_1708}), .a ({signal_5269, signal_5267}), .clk (CLK), .r (Fresh[492]), .c ({signal_2792, signal_1764}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1621 ( .s ({signal_5157, signal_5155}), .b ({signal_2630, signal_1709}), .a ({signal_2611, signal_899}), .clk (CLK), .r (Fresh[493]), .c ({signal_2731, signal_1765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1622 ( .s ({signal_5157, signal_5155}), .b ({signal_2611, signal_899}), .a ({signal_2630, signal_1709}), .clk (CLK), .r (Fresh[494]), .c ({signal_2732, signal_1766}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1623 ( .s ({signal_5169, signal_5163}), .b ({signal_2630, signal_1709}), .a ({signal_2611, signal_899}), .clk (CLK), .r (Fresh[495]), .c ({signal_2733, signal_1767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1624 ( .s ({signal_5213, signal_5205}), .b ({signal_2710, signal_1710}), .a ({signal_2676, signal_911}), .clk (CLK), .r (Fresh[496]), .c ({signal_2793, signal_1768}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1625 ( .s ({signal_5213, signal_5205}), .b ({signal_2676, signal_911}), .a ({signal_2710, signal_1710}), .clk (CLK), .r (Fresh[497]), .c ({signal_2794, signal_1769}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1626 ( .s ({signal_4513, signal_4507}), .b ({signal_2710, signal_1710}), .a ({signal_2676, signal_911}), .clk (CLK), .r (Fresh[498]), .c ({signal_2795, signal_1770}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1627 ( .s ({signal_4849, signal_4841}), .b ({signal_2714, signal_1712}), .a ({signal_2713, signal_1711}), .clk (CLK), .r (Fresh[499]), .c ({signal_2796, signal_1771}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1628 ( .s ({signal_5173, signal_5171}), .b ({signal_2656, signal_1663}), .a ({signal_5185, signal_5183}), .clk (CLK), .r (Fresh[500]), .c ({signal_2797, signal_1772}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1629 ( .s ({signal_5173, signal_5171}), .b ({signal_2662, signal_1669}), .a ({signal_5177, signal_5175}), .clk (CLK), .r (Fresh[501]), .c ({signal_2798, signal_1773}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1630 ( .s ({signal_5173, signal_5171}), .b ({signal_2659, signal_1666}), .a ({signal_5273, signal_5271}), .clk (CLK), .r (Fresh[502]), .c ({signal_2799, signal_1774}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1631 ( .s ({signal_5173, signal_5171}), .b ({signal_2715, signal_1713}), .a ({signal_5181, signal_5179}), .clk (CLK), .r (Fresh[503]), .c ({signal_2800, signal_1775}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1632 ( .s ({signal_4833, signal_4829}), .b ({signal_2718, signal_1716}), .a ({signal_2717, signal_1715}), .clk (CLK), .r (Fresh[504]), .c ({signal_2801, signal_1776}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1633 ( .s ({signal_4833, signal_4829}), .b ({signal_2717, signal_1715}), .a ({signal_2718, signal_1716}), .clk (CLK), .r (Fresh[505]), .c ({signal_2802, signal_1777}) ) ;
    buf_clk cell_3131 ( .C (CLK), .D (signal_5274), .Q (signal_5275) ) ;
    buf_clk cell_3133 ( .C (CLK), .D (signal_5276), .Q (signal_5277) ) ;
    buf_clk cell_3135 ( .C (CLK), .D (signal_5278), .Q (signal_5279) ) ;
    buf_clk cell_3137 ( .C (CLK), .D (signal_5280), .Q (signal_5281) ) ;
    buf_clk cell_3139 ( .C (CLK), .D (signal_5282), .Q (signal_5283) ) ;
    buf_clk cell_3141 ( .C (CLK), .D (signal_5284), .Q (signal_5285) ) ;
    buf_clk cell_3143 ( .C (CLK), .D (signal_5286), .Q (signal_5287) ) ;
    buf_clk cell_3145 ( .C (CLK), .D (signal_5288), .Q (signal_5289) ) ;
    buf_clk cell_3147 ( .C (CLK), .D (signal_5290), .Q (signal_5291) ) ;
    buf_clk cell_3149 ( .C (CLK), .D (signal_5292), .Q (signal_5293) ) ;
    buf_clk cell_3151 ( .C (CLK), .D (signal_5294), .Q (signal_5295) ) ;
    buf_clk cell_3153 ( .C (CLK), .D (signal_5296), .Q (signal_5297) ) ;
    buf_clk cell_3155 ( .C (CLK), .D (signal_5298), .Q (signal_5299) ) ;
    buf_clk cell_3157 ( .C (CLK), .D (signal_5300), .Q (signal_5301) ) ;
    buf_clk cell_3159 ( .C (CLK), .D (signal_5302), .Q (signal_5303) ) ;
    buf_clk cell_3161 ( .C (CLK), .D (signal_5304), .Q (signal_5305) ) ;
    buf_clk cell_3163 ( .C (CLK), .D (signal_5306), .Q (signal_5307) ) ;
    buf_clk cell_3165 ( .C (CLK), .D (signal_5308), .Q (signal_5309) ) ;
    buf_clk cell_3167 ( .C (CLK), .D (signal_5310), .Q (signal_5311) ) ;
    buf_clk cell_3169 ( .C (CLK), .D (signal_5312), .Q (signal_5313) ) ;
    buf_clk cell_3171 ( .C (CLK), .D (signal_5314), .Q (signal_5315) ) ;
    buf_clk cell_3173 ( .C (CLK), .D (signal_5316), .Q (signal_5317) ) ;
    buf_clk cell_3175 ( .C (CLK), .D (signal_5318), .Q (signal_5319) ) ;
    buf_clk cell_3177 ( .C (CLK), .D (signal_5320), .Q (signal_5321) ) ;
    buf_clk cell_3179 ( .C (CLK), .D (signal_5322), .Q (signal_5323) ) ;
    buf_clk cell_3181 ( .C (CLK), .D (signal_5324), .Q (signal_5325) ) ;
    buf_clk cell_3183 ( .C (CLK), .D (signal_5326), .Q (signal_5327) ) ;
    buf_clk cell_3185 ( .C (CLK), .D (signal_5328), .Q (signal_5329) ) ;
    buf_clk cell_3187 ( .C (CLK), .D (signal_5330), .Q (signal_5331) ) ;
    buf_clk cell_3189 ( .C (CLK), .D (signal_5332), .Q (signal_5333) ) ;
    buf_clk cell_3191 ( .C (CLK), .D (signal_5334), .Q (signal_5335) ) ;
    buf_clk cell_3193 ( .C (CLK), .D (signal_5336), .Q (signal_5337) ) ;
    buf_clk cell_3201 ( .C (CLK), .D (signal_5344), .Q (signal_5345) ) ;
    buf_clk cell_3209 ( .C (CLK), .D (signal_5352), .Q (signal_5353) ) ;
    buf_clk cell_3211 ( .C (CLK), .D (signal_5354), .Q (signal_5355) ) ;
    buf_clk cell_3213 ( .C (CLK), .D (signal_5356), .Q (signal_5357) ) ;
    buf_clk cell_3215 ( .C (CLK), .D (signal_5358), .Q (signal_5359) ) ;
    buf_clk cell_3217 ( .C (CLK), .D (signal_5360), .Q (signal_5361) ) ;
    buf_clk cell_3219 ( .C (CLK), .D (signal_5362), .Q (signal_5363) ) ;
    buf_clk cell_3221 ( .C (CLK), .D (signal_5364), .Q (signal_5365) ) ;
    buf_clk cell_3223 ( .C (CLK), .D (signal_5366), .Q (signal_5367) ) ;
    buf_clk cell_3225 ( .C (CLK), .D (signal_5368), .Q (signal_5369) ) ;
    buf_clk cell_3227 ( .C (CLK), .D (signal_5370), .Q (signal_5371) ) ;
    buf_clk cell_3229 ( .C (CLK), .D (signal_5372), .Q (signal_5373) ) ;
    buf_clk cell_3233 ( .C (CLK), .D (signal_5376), .Q (signal_5377) ) ;
    buf_clk cell_3237 ( .C (CLK), .D (signal_5380), .Q (signal_5381) ) ;
    buf_clk cell_3239 ( .C (CLK), .D (signal_5382), .Q (signal_5383) ) ;
    buf_clk cell_3241 ( .C (CLK), .D (signal_5384), .Q (signal_5385) ) ;
    buf_clk cell_3243 ( .C (CLK), .D (signal_5386), .Q (signal_5387) ) ;
    buf_clk cell_3245 ( .C (CLK), .D (signal_5388), .Q (signal_5389) ) ;
    buf_clk cell_3247 ( .C (CLK), .D (signal_5390), .Q (signal_5391) ) ;
    buf_clk cell_3249 ( .C (CLK), .D (signal_5392), .Q (signal_5393) ) ;
    buf_clk cell_3251 ( .C (CLK), .D (signal_5394), .Q (signal_5395) ) ;
    buf_clk cell_3253 ( .C (CLK), .D (signal_5396), .Q (signal_5397) ) ;
    buf_clk cell_3255 ( .C (CLK), .D (signal_5398), .Q (signal_5399) ) ;
    buf_clk cell_3257 ( .C (CLK), .D (signal_5400), .Q (signal_5401) ) ;
    buf_clk cell_3259 ( .C (CLK), .D (signal_5402), .Q (signal_5403) ) ;
    buf_clk cell_3261 ( .C (CLK), .D (signal_5404), .Q (signal_5405) ) ;
    buf_clk cell_3263 ( .C (CLK), .D (signal_5406), .Q (signal_5407) ) ;
    buf_clk cell_3265 ( .C (CLK), .D (signal_5408), .Q (signal_5409) ) ;
    buf_clk cell_3267 ( .C (CLK), .D (signal_5410), .Q (signal_5411) ) ;
    buf_clk cell_3269 ( .C (CLK), .D (signal_5412), .Q (signal_5413) ) ;
    buf_clk cell_3271 ( .C (CLK), .D (signal_5414), .Q (signal_5415) ) ;
    buf_clk cell_3273 ( .C (CLK), .D (signal_5416), .Q (signal_5417) ) ;
    buf_clk cell_3275 ( .C (CLK), .D (signal_5418), .Q (signal_5419) ) ;
    buf_clk cell_3279 ( .C (CLK), .D (signal_5422), .Q (signal_5423) ) ;
    buf_clk cell_3287 ( .C (CLK), .D (signal_5430), .Q (signal_5431) ) ;
    buf_clk cell_3291 ( .C (CLK), .D (signal_5434), .Q (signal_5435) ) ;
    buf_clk cell_3301 ( .C (CLK), .D (signal_5444), .Q (signal_5445) ) ;
    buf_clk cell_3307 ( .C (CLK), .D (signal_5450), .Q (signal_5451) ) ;
    buf_clk cell_3323 ( .C (CLK), .D (signal_5466), .Q (signal_5467) ) ;
    buf_clk cell_3331 ( .C (CLK), .D (signal_5474), .Q (signal_5475) ) ;
    buf_clk cell_3341 ( .C (CLK), .D (signal_5484), .Q (signal_5485) ) ;
    buf_clk cell_3347 ( .C (CLK), .D (signal_5490), .Q (signal_5491) ) ;
    buf_clk cell_3359 ( .C (CLK), .D (signal_5502), .Q (signal_5503) ) ;
    buf_clk cell_3367 ( .C (CLK), .D (signal_5510), .Q (signal_5511) ) ;
    buf_clk cell_3399 ( .C (CLK), .D (signal_5542), .Q (signal_5543) ) ;
    buf_clk cell_3403 ( .C (CLK), .D (signal_5546), .Q (signal_5547) ) ;
    buf_clk cell_3407 ( .C (CLK), .D (signal_5550), .Q (signal_5551) ) ;
    buf_clk cell_3411 ( .C (CLK), .D (signal_5554), .Q (signal_5555) ) ;
    buf_clk cell_3439 ( .C (CLK), .D (signal_5582), .Q (signal_5583) ) ;
    buf_clk cell_3455 ( .C (CLK), .D (signal_5598), .Q (signal_5599) ) ;
    buf_clk cell_3471 ( .C (CLK), .D (signal_5614), .Q (signal_5615) ) ;
    buf_clk cell_3479 ( .C (CLK), .D (signal_5622), .Q (signal_5623) ) ;
    buf_clk cell_3495 ( .C (CLK), .D (signal_5638), .Q (signal_5639) ) ;
    buf_clk cell_3511 ( .C (CLK), .D (signal_5654), .Q (signal_5655) ) ;
    buf_clk cell_3519 ( .C (CLK), .D (signal_5662), .Q (signal_5663) ) ;
    buf_clk cell_3535 ( .C (CLK), .D (signal_5678), .Q (signal_5679) ) ;
    buf_clk cell_3551 ( .C (CLK), .D (signal_5694), .Q (signal_5695) ) ;
    buf_clk cell_3567 ( .C (CLK), .D (signal_5710), .Q (signal_5711) ) ;
    buf_clk cell_3583 ( .C (CLK), .D (signal_5726), .Q (signal_5727) ) ;
    buf_clk cell_3643 ( .C (CLK), .D (signal_5786), .Q (signal_5787) ) ;
    buf_clk cell_3659 ( .C (CLK), .D (signal_5802), .Q (signal_5803) ) ;
    buf_clk cell_3675 ( .C (CLK), .D (signal_5818), .Q (signal_5819) ) ;
    buf_clk cell_3691 ( .C (CLK), .D (signal_5834), .Q (signal_5835) ) ;
    buf_clk cell_3707 ( .C (CLK), .D (signal_5850), .Q (signal_5851) ) ;
    buf_clk cell_3723 ( .C (CLK), .D (signal_5866), .Q (signal_5867) ) ;
    buf_clk cell_3739 ( .C (CLK), .D (signal_5882), .Q (signal_5883) ) ;
    buf_clk cell_3755 ( .C (CLK), .D (signal_5898), .Q (signal_5899) ) ;
    buf_clk cell_3771 ( .C (CLK), .D (signal_5914), .Q (signal_5915) ) ;
    buf_clk cell_3787 ( .C (CLK), .D (signal_5930), .Q (signal_5931) ) ;
    buf_clk cell_3803 ( .C (CLK), .D (signal_5946), .Q (signal_5947) ) ;
    buf_clk cell_3811 ( .C (CLK), .D (signal_5954), .Q (signal_5955) ) ;
    buf_clk cell_3831 ( .C (CLK), .D (signal_5974), .Q (signal_5975) ) ;
    buf_clk cell_3839 ( .C (CLK), .D (signal_5982), .Q (signal_5983) ) ;
    buf_clk cell_3847 ( .C (CLK), .D (signal_5990), .Q (signal_5991) ) ;
    buf_clk cell_3855 ( .C (CLK), .D (signal_5998), .Q (signal_5999) ) ;
    buf_clk cell_3871 ( .C (CLK), .D (signal_6014), .Q (signal_6015) ) ;
    buf_clk cell_3879 ( .C (CLK), .D (signal_6022), .Q (signal_6023) ) ;
    buf_clk cell_3895 ( .C (CLK), .D (signal_6038), .Q (signal_6039) ) ;
    buf_clk cell_3911 ( .C (CLK), .D (signal_6054), .Q (signal_6055) ) ;
    buf_clk cell_3927 ( .C (CLK), .D (signal_6070), .Q (signal_6071) ) ;
    buf_clk cell_3943 ( .C (CLK), .D (signal_6086), .Q (signal_6087) ) ;
    buf_clk cell_3959 ( .C (CLK), .D (signal_6102), .Q (signal_6103) ) ;
    buf_clk cell_3975 ( .C (CLK), .D (signal_6118), .Q (signal_6119) ) ;
    buf_clk cell_3991 ( .C (CLK), .D (signal_6134), .Q (signal_6135) ) ;
    buf_clk cell_4007 ( .C (CLK), .D (signal_6150), .Q (signal_6151) ) ;
    buf_clk cell_4023 ( .C (CLK), .D (signal_6166), .Q (signal_6167) ) ;
    buf_clk cell_4039 ( .C (CLK), .D (signal_6182), .Q (signal_6183) ) ;
    buf_clk cell_4055 ( .C (CLK), .D (signal_6198), .Q (signal_6199) ) ;
    buf_clk cell_4071 ( .C (CLK), .D (signal_6214), .Q (signal_6215) ) ;
    buf_clk cell_4087 ( .C (CLK), .D (signal_6230), .Q (signal_6231) ) ;
    buf_clk cell_4103 ( .C (CLK), .D (signal_6246), .Q (signal_6247) ) ;
    buf_clk cell_4113 ( .C (CLK), .D (signal_6256), .Q (signal_6257) ) ;
    buf_clk cell_4123 ( .C (CLK), .D (signal_6266), .Q (signal_6267) ) ;
    buf_clk cell_4143 ( .C (CLK), .D (signal_6286), .Q (signal_6287) ) ;
    buf_clk cell_4151 ( .C (CLK), .D (signal_6294), .Q (signal_6295) ) ;
    buf_clk cell_4161 ( .C (CLK), .D (signal_6304), .Q (signal_6305) ) ;
    buf_clk cell_4171 ( .C (CLK), .D (signal_6314), .Q (signal_6315) ) ;
    buf_clk cell_4187 ( .C (CLK), .D (signal_6330), .Q (signal_6331) ) ;
    buf_clk cell_4199 ( .C (CLK), .D (signal_6342), .Q (signal_6343) ) ;
    buf_clk cell_4211 ( .C (CLK), .D (signal_6354), .Q (signal_6355) ) ;
    buf_clk cell_4219 ( .C (CLK), .D (signal_6362), .Q (signal_6363) ) ;
    buf_clk cell_4227 ( .C (CLK), .D (signal_6370), .Q (signal_6371) ) ;
    buf_clk cell_4239 ( .C (CLK), .D (signal_6382), .Q (signal_6383) ) ;
    buf_clk cell_4251 ( .C (CLK), .D (signal_6394), .Q (signal_6395) ) ;
    buf_clk cell_4265 ( .C (CLK), .D (signal_6408), .Q (signal_6409) ) ;
    buf_clk cell_4279 ( .C (CLK), .D (signal_6422), .Q (signal_6423) ) ;
    buf_clk cell_4295 ( .C (CLK), .D (signal_6438), .Q (signal_6439) ) ;
    buf_clk cell_4311 ( .C (CLK), .D (signal_6454), .Q (signal_6455) ) ;
    buf_clk cell_4327 ( .C (CLK), .D (signal_6470), .Q (signal_6471) ) ;
    buf_clk cell_4343 ( .C (CLK), .D (signal_6486), .Q (signal_6487) ) ;
    buf_clk cell_4359 ( .C (CLK), .D (signal_6502), .Q (signal_6503) ) ;
    buf_clk cell_4375 ( .C (CLK), .D (signal_6518), .Q (signal_6519) ) ;
    buf_clk cell_4391 ( .C (CLK), .D (signal_6534), .Q (signal_6535) ) ;
    buf_clk cell_4407 ( .C (CLK), .D (signal_6550), .Q (signal_6551) ) ;
    buf_clk cell_4423 ( .C (CLK), .D (signal_6566), .Q (signal_6567) ) ;
    buf_clk cell_4439 ( .C (CLK), .D (signal_6582), .Q (signal_6583) ) ;
    buf_clk cell_4455 ( .C (CLK), .D (signal_6598), .Q (signal_6599) ) ;
    buf_clk cell_4471 ( .C (CLK), .D (signal_6614), .Q (signal_6615) ) ;
    buf_clk cell_4487 ( .C (CLK), .D (signal_6630), .Q (signal_6631) ) ;
    buf_clk cell_4503 ( .C (CLK), .D (signal_6646), .Q (signal_6647) ) ;
    buf_clk cell_4519 ( .C (CLK), .D (signal_6662), .Q (signal_6663) ) ;
    buf_clk cell_4535 ( .C (CLK), .D (signal_6678), .Q (signal_6679) ) ;
    buf_clk cell_4545 ( .C (CLK), .D (signal_6688), .Q (signal_6689) ) ;
    buf_clk cell_4555 ( .C (CLK), .D (signal_6698), .Q (signal_6699) ) ;
    buf_clk cell_4563 ( .C (CLK), .D (signal_6706), .Q (signal_6707) ) ;
    buf_clk cell_4571 ( .C (CLK), .D (signal_6714), .Q (signal_6715) ) ;
    buf_clk cell_4583 ( .C (CLK), .D (signal_6726), .Q (signal_6727) ) ;
    buf_clk cell_4595 ( .C (CLK), .D (signal_6738), .Q (signal_6739) ) ;
    buf_clk cell_4609 ( .C (CLK), .D (signal_6752), .Q (signal_6753) ) ;
    buf_clk cell_4623 ( .C (CLK), .D (signal_6766), .Q (signal_6767) ) ;
    buf_clk cell_4639 ( .C (CLK), .D (signal_6782), .Q (signal_6783) ) ;
    buf_clk cell_4655 ( .C (CLK), .D (signal_6798), .Q (signal_6799) ) ;
    buf_clk cell_4675 ( .C (CLK), .D (signal_6818), .Q (signal_6819) ) ;
    buf_clk cell_4683 ( .C (CLK), .D (signal_6826), .Q (signal_6827) ) ;
    buf_clk cell_4693 ( .C (CLK), .D (signal_6836), .Q (signal_6837) ) ;
    buf_clk cell_4703 ( .C (CLK), .D (signal_6846), .Q (signal_6847) ) ;
    buf_clk cell_4715 ( .C (CLK), .D (signal_6858), .Q (signal_6859) ) ;
    buf_clk cell_4727 ( .C (CLK), .D (signal_6870), .Q (signal_6871) ) ;
    buf_clk cell_4735 ( .C (CLK), .D (signal_6878), .Q (signal_6879) ) ;
    buf_clk cell_4751 ( .C (CLK), .D (signal_6894), .Q (signal_6895) ) ;
    buf_clk cell_4767 ( .C (CLK), .D (signal_6910), .Q (signal_6911) ) ;
    buf_clk cell_4783 ( .C (CLK), .D (signal_6926), .Q (signal_6927) ) ;
    buf_clk cell_4799 ( .C (CLK), .D (signal_6942), .Q (signal_6943) ) ;
    buf_clk cell_4815 ( .C (CLK), .D (signal_6958), .Q (signal_6959) ) ;
    buf_clk cell_4831 ( .C (CLK), .D (signal_6974), .Q (signal_6975) ) ;
    buf_clk cell_4847 ( .C (CLK), .D (signal_6990), .Q (signal_6991) ) ;
    buf_clk cell_4863 ( .C (CLK), .D (signal_7006), .Q (signal_7007) ) ;
    buf_clk cell_4879 ( .C (CLK), .D (signal_7022), .Q (signal_7023) ) ;
    buf_clk cell_4895 ( .C (CLK), .D (signal_7038), .Q (signal_7039) ) ;
    buf_clk cell_4911 ( .C (CLK), .D (signal_7054), .Q (signal_7055) ) ;
    buf_clk cell_4927 ( .C (CLK), .D (signal_7070), .Q (signal_7071) ) ;
    buf_clk cell_4943 ( .C (CLK), .D (signal_7086), .Q (signal_7087) ) ;
    buf_clk cell_4959 ( .C (CLK), .D (signal_7102), .Q (signal_7103) ) ;
    buf_clk cell_4975 ( .C (CLK), .D (signal_7118), .Q (signal_7119) ) ;
    buf_clk cell_4991 ( .C (CLK), .D (signal_7134), .Q (signal_7135) ) ;
    buf_clk cell_5007 ( .C (CLK), .D (signal_7150), .Q (signal_7151) ) ;
    buf_clk cell_5023 ( .C (CLK), .D (signal_7166), .Q (signal_7167) ) ;
    buf_clk cell_5039 ( .C (CLK), .D (signal_7182), .Q (signal_7183) ) ;
    buf_clk cell_5055 ( .C (CLK), .D (signal_7198), .Q (signal_7199) ) ;
    buf_clk cell_5071 ( .C (CLK), .D (signal_7214), .Q (signal_7215) ) ;
    buf_clk cell_5087 ( .C (CLK), .D (signal_7230), .Q (signal_7231) ) ;
    buf_clk cell_5103 ( .C (CLK), .D (signal_7246), .Q (signal_7247) ) ;
    buf_clk cell_5119 ( .C (CLK), .D (signal_7262), .Q (signal_7263) ) ;
    buf_clk cell_5135 ( .C (CLK), .D (signal_7278), .Q (signal_7279) ) ;
    buf_clk cell_5151 ( .C (CLK), .D (signal_7294), .Q (signal_7295) ) ;
    buf_clk cell_5167 ( .C (CLK), .D (signal_7310), .Q (signal_7311) ) ;
    buf_clk cell_5183 ( .C (CLK), .D (signal_7326), .Q (signal_7327) ) ;
    buf_clk cell_5199 ( .C (CLK), .D (signal_7342), .Q (signal_7343) ) ;
    buf_clk cell_5215 ( .C (CLK), .D (signal_7358), .Q (signal_7359) ) ;
    buf_clk cell_5231 ( .C (CLK), .D (signal_7374), .Q (signal_7375) ) ;
    buf_clk cell_5247 ( .C (CLK), .D (signal_7390), .Q (signal_7391) ) ;
    buf_clk cell_5263 ( .C (CLK), .D (signal_7406), .Q (signal_7407) ) ;
    buf_clk cell_5279 ( .C (CLK), .D (signal_7422), .Q (signal_7423) ) ;
    buf_clk cell_5295 ( .C (CLK), .D (signal_7438), .Q (signal_7439) ) ;
    buf_clk cell_5311 ( .C (CLK), .D (signal_7454), .Q (signal_7455) ) ;
    buf_clk cell_5327 ( .C (CLK), .D (signal_7470), .Q (signal_7471) ) ;
    buf_clk cell_5343 ( .C (CLK), .D (signal_7486), .Q (signal_7487) ) ;
    buf_clk cell_5359 ( .C (CLK), .D (signal_7502), .Q (signal_7503) ) ;
    buf_clk cell_5375 ( .C (CLK), .D (signal_7518), .Q (signal_7519) ) ;
    buf_clk cell_5391 ( .C (CLK), .D (signal_7534), .Q (signal_7535) ) ;
    buf_clk cell_5407 ( .C (CLK), .D (signal_7550), .Q (signal_7551) ) ;
    buf_clk cell_5423 ( .C (CLK), .D (signal_7566), .Q (signal_7567) ) ;
    buf_clk cell_5439 ( .C (CLK), .D (signal_7582), .Q (signal_7583) ) ;
    buf_clk cell_5455 ( .C (CLK), .D (signal_7598), .Q (signal_7599) ) ;
    buf_clk cell_5471 ( .C (CLK), .D (signal_7614), .Q (signal_7615) ) ;
    buf_clk cell_5487 ( .C (CLK), .D (signal_7630), .Q (signal_7631) ) ;
    buf_clk cell_5503 ( .C (CLK), .D (signal_7646), .Q (signal_7647) ) ;
    buf_clk cell_5519 ( .C (CLK), .D (signal_7662), .Q (signal_7663) ) ;
    buf_clk cell_5535 ( .C (CLK), .D (signal_7678), .Q (signal_7679) ) ;
    buf_clk cell_5551 ( .C (CLK), .D (signal_7694), .Q (signal_7695) ) ;
    buf_clk cell_5567 ( .C (CLK), .D (signal_7710), .Q (signal_7711) ) ;
    buf_clk cell_5583 ( .C (CLK), .D (signal_7726), .Q (signal_7727) ) ;
    buf_clk cell_5599 ( .C (CLK), .D (signal_7742), .Q (signal_7743) ) ;
    buf_clk cell_5615 ( .C (CLK), .D (signal_7758), .Q (signal_7759) ) ;
    buf_clk cell_5631 ( .C (CLK), .D (signal_7774), .Q (signal_7775) ) ;
    buf_clk cell_5647 ( .C (CLK), .D (signal_7790), .Q (signal_7791) ) ;
    buf_clk cell_5663 ( .C (CLK), .D (signal_7806), .Q (signal_7807) ) ;
    buf_clk cell_5679 ( .C (CLK), .D (signal_7822), .Q (signal_7823) ) ;
    buf_clk cell_5695 ( .C (CLK), .D (signal_7838), .Q (signal_7839) ) ;
    buf_clk cell_5711 ( .C (CLK), .D (signal_7854), .Q (signal_7855) ) ;
    buf_clk cell_5727 ( .C (CLK), .D (signal_7870), .Q (signal_7871) ) ;
    buf_clk cell_5743 ( .C (CLK), .D (signal_7886), .Q (signal_7887) ) ;
    buf_clk cell_5759 ( .C (CLK), .D (signal_7902), .Q (signal_7903) ) ;
    buf_clk cell_5775 ( .C (CLK), .D (signal_7918), .Q (signal_7919) ) ;
    buf_clk cell_5791 ( .C (CLK), .D (signal_7934), .Q (signal_7935) ) ;
    buf_clk cell_5807 ( .C (CLK), .D (signal_7950), .Q (signal_7951) ) ;
    buf_clk cell_5823 ( .C (CLK), .D (signal_7966), .Q (signal_7967) ) ;
    buf_clk cell_5839 ( .C (CLK), .D (signal_7982), .Q (signal_7983) ) ;
    buf_clk cell_5855 ( .C (CLK), .D (signal_7998), .Q (signal_7999) ) ;
    buf_clk cell_5871 ( .C (CLK), .D (signal_8014), .Q (signal_8015) ) ;
    buf_clk cell_5887 ( .C (CLK), .D (signal_8030), .Q (signal_8031) ) ;
    buf_clk cell_5903 ( .C (CLK), .D (signal_8046), .Q (signal_8047) ) ;
    buf_clk cell_5919 ( .C (CLK), .D (signal_8062), .Q (signal_8063) ) ;
    buf_clk cell_5935 ( .C (CLK), .D (signal_8078), .Q (signal_8079) ) ;
    buf_clk cell_5951 ( .C (CLK), .D (signal_8094), .Q (signal_8095) ) ;
    buf_clk cell_5967 ( .C (CLK), .D (signal_8110), .Q (signal_8111) ) ;
    buf_clk cell_5983 ( .C (CLK), .D (signal_8126), .Q (signal_8127) ) ;
    buf_clk cell_5999 ( .C (CLK), .D (signal_8142), .Q (signal_8143) ) ;
    buf_clk cell_6015 ( .C (CLK), .D (signal_8158), .Q (signal_8159) ) ;
    buf_clk cell_6031 ( .C (CLK), .D (signal_8174), .Q (signal_8175) ) ;
    buf_clk cell_6047 ( .C (CLK), .D (signal_8190), .Q (signal_8191) ) ;
    buf_clk cell_6063 ( .C (CLK), .D (signal_8206), .Q (signal_8207) ) ;
    buf_clk cell_6079 ( .C (CLK), .D (signal_8222), .Q (signal_8223) ) ;
    buf_clk cell_6095 ( .C (CLK), .D (signal_8238), .Q (signal_8239) ) ;
    buf_clk cell_6111 ( .C (CLK), .D (signal_8254), .Q (signal_8255) ) ;
    buf_clk cell_6127 ( .C (CLK), .D (signal_8270), .Q (signal_8271) ) ;
    buf_clk cell_6143 ( .C (CLK), .D (signal_8286), .Q (signal_8287) ) ;
    buf_clk cell_6159 ( .C (CLK), .D (signal_8302), .Q (signal_8303) ) ;
    buf_clk cell_6175 ( .C (CLK), .D (signal_8318), .Q (signal_8319) ) ;
    buf_clk cell_6191 ( .C (CLK), .D (signal_8334), .Q (signal_8335) ) ;
    buf_clk cell_6207 ( .C (CLK), .D (signal_8350), .Q (signal_8351) ) ;
    buf_clk cell_6223 ( .C (CLK), .D (signal_8366), .Q (signal_8367) ) ;
    buf_clk cell_6239 ( .C (CLK), .D (signal_8382), .Q (signal_8383) ) ;
    buf_clk cell_6255 ( .C (CLK), .D (signal_8398), .Q (signal_8399) ) ;
    buf_clk cell_6271 ( .C (CLK), .D (signal_8414), .Q (signal_8415) ) ;
    buf_clk cell_6287 ( .C (CLK), .D (signal_8430), .Q (signal_8431) ) ;
    buf_clk cell_6303 ( .C (CLK), .D (signal_8446), .Q (signal_8447) ) ;
    buf_clk cell_6319 ( .C (CLK), .D (signal_8462), .Q (signal_8463) ) ;
    buf_clk cell_6335 ( .C (CLK), .D (signal_8478), .Q (signal_8479) ) ;
    buf_clk cell_6351 ( .C (CLK), .D (signal_8494), .Q (signal_8495) ) ;
    buf_clk cell_6367 ( .C (CLK), .D (signal_8510), .Q (signal_8511) ) ;
    buf_clk cell_6383 ( .C (CLK), .D (signal_8526), .Q (signal_8527) ) ;
    buf_clk cell_6399 ( .C (CLK), .D (signal_8542), .Q (signal_8543) ) ;
    buf_clk cell_6407 ( .C (CLK), .D (signal_8550), .Q (signal_8551) ) ;
    buf_clk cell_6415 ( .C (CLK), .D (signal_8558), .Q (signal_8559) ) ;
    buf_clk cell_6423 ( .C (CLK), .D (signal_8566), .Q (signal_8567) ) ;
    buf_clk cell_6431 ( .C (CLK), .D (signal_8574), .Q (signal_8575) ) ;
    buf_clk cell_6439 ( .C (CLK), .D (signal_8582), .Q (signal_8583) ) ;
    buf_clk cell_6447 ( .C (CLK), .D (signal_8590), .Q (signal_8591) ) ;
    buf_clk cell_6455 ( .C (CLK), .D (signal_8598), .Q (signal_8599) ) ;
    buf_clk cell_6463 ( .C (CLK), .D (signal_8606), .Q (signal_8607) ) ;
    buf_clk cell_6471 ( .C (CLK), .D (signal_8614), .Q (signal_8615) ) ;
    buf_clk cell_6479 ( .C (CLK), .D (signal_8622), .Q (signal_8623) ) ;
    buf_clk cell_6487 ( .C (CLK), .D (signal_8630), .Q (signal_8631) ) ;
    buf_clk cell_6495 ( .C (CLK), .D (signal_8638), .Q (signal_8639) ) ;
    buf_clk cell_6503 ( .C (CLK), .D (signal_8646), .Q (signal_8647) ) ;
    buf_clk cell_6511 ( .C (CLK), .D (signal_8654), .Q (signal_8655) ) ;
    buf_clk cell_6519 ( .C (CLK), .D (signal_8662), .Q (signal_8663) ) ;
    buf_clk cell_6527 ( .C (CLK), .D (signal_8670), .Q (signal_8671) ) ;
    buf_clk cell_6535 ( .C (CLK), .D (signal_8678), .Q (signal_8679) ) ;
    buf_clk cell_6543 ( .C (CLK), .D (signal_8686), .Q (signal_8687) ) ;
    buf_clk cell_6551 ( .C (CLK), .D (signal_8694), .Q (signal_8695) ) ;
    buf_clk cell_6559 ( .C (CLK), .D (signal_8702), .Q (signal_8703) ) ;
    buf_clk cell_6567 ( .C (CLK), .D (signal_8710), .Q (signal_8711) ) ;
    buf_clk cell_6575 ( .C (CLK), .D (signal_8718), .Q (signal_8719) ) ;
    buf_clk cell_6583 ( .C (CLK), .D (signal_8726), .Q (signal_8727) ) ;
    buf_clk cell_6591 ( .C (CLK), .D (signal_8734), .Q (signal_8735) ) ;
    buf_clk cell_6599 ( .C (CLK), .D (signal_8742), .Q (signal_8743) ) ;
    buf_clk cell_6607 ( .C (CLK), .D (signal_8750), .Q (signal_8751) ) ;
    buf_clk cell_6615 ( .C (CLK), .D (signal_8758), .Q (signal_8759) ) ;
    buf_clk cell_6623 ( .C (CLK), .D (signal_8766), .Q (signal_8767) ) ;
    buf_clk cell_6631 ( .C (CLK), .D (signal_8774), .Q (signal_8775) ) ;
    buf_clk cell_6639 ( .C (CLK), .D (signal_8782), .Q (signal_8783) ) ;
    buf_clk cell_6647 ( .C (CLK), .D (signal_8790), .Q (signal_8791) ) ;
    buf_clk cell_6655 ( .C (CLK), .D (signal_8798), .Q (signal_8799) ) ;
    buf_clk cell_6663 ( .C (CLK), .D (signal_8806), .Q (signal_8807) ) ;
    buf_clk cell_6671 ( .C (CLK), .D (signal_8814), .Q (signal_8815) ) ;
    buf_clk cell_6679 ( .C (CLK), .D (signal_8822), .Q (signal_8823) ) ;
    buf_clk cell_6687 ( .C (CLK), .D (signal_8830), .Q (signal_8831) ) ;
    buf_clk cell_6695 ( .C (CLK), .D (signal_8838), .Q (signal_8839) ) ;
    buf_clk cell_6703 ( .C (CLK), .D (signal_8846), .Q (signal_8847) ) ;
    buf_clk cell_6711 ( .C (CLK), .D (signal_8854), .Q (signal_8855) ) ;
    buf_clk cell_6719 ( .C (CLK), .D (signal_8862), .Q (signal_8863) ) ;
    buf_clk cell_6727 ( .C (CLK), .D (signal_8870), .Q (signal_8871) ) ;
    buf_clk cell_6735 ( .C (CLK), .D (signal_8878), .Q (signal_8879) ) ;
    buf_clk cell_6743 ( .C (CLK), .D (signal_8886), .Q (signal_8887) ) ;
    buf_clk cell_6751 ( .C (CLK), .D (signal_8894), .Q (signal_8895) ) ;
    buf_clk cell_6759 ( .C (CLK), .D (signal_8902), .Q (signal_8903) ) ;
    buf_clk cell_6767 ( .C (CLK), .D (signal_8910), .Q (signal_8911) ) ;
    buf_clk cell_6775 ( .C (CLK), .D (signal_8918), .Q (signal_8919) ) ;
    buf_clk cell_6783 ( .C (CLK), .D (signal_8926), .Q (signal_8927) ) ;
    buf_clk cell_6791 ( .C (CLK), .D (signal_8934), .Q (signal_8935) ) ;
    buf_clk cell_6799 ( .C (CLK), .D (signal_8942), .Q (signal_8943) ) ;
    buf_clk cell_6807 ( .C (CLK), .D (signal_8950), .Q (signal_8951) ) ;
    buf_clk cell_6815 ( .C (CLK), .D (signal_8958), .Q (signal_8959) ) ;
    buf_clk cell_6823 ( .C (CLK), .D (signal_8966), .Q (signal_8967) ) ;
    buf_clk cell_6831 ( .C (CLK), .D (signal_8974), .Q (signal_8975) ) ;
    buf_clk cell_6839 ( .C (CLK), .D (signal_8982), .Q (signal_8983) ) ;
    buf_clk cell_6847 ( .C (CLK), .D (signal_8990), .Q (signal_8991) ) ;
    buf_clk cell_6855 ( .C (CLK), .D (signal_8998), .Q (signal_8999) ) ;
    buf_clk cell_6863 ( .C (CLK), .D (signal_9006), .Q (signal_9007) ) ;
    buf_clk cell_6871 ( .C (CLK), .D (signal_9014), .Q (signal_9015) ) ;
    buf_clk cell_6879 ( .C (CLK), .D (signal_9022), .Q (signal_9023) ) ;
    buf_clk cell_6887 ( .C (CLK), .D (signal_9030), .Q (signal_9031) ) ;
    buf_clk cell_6895 ( .C (CLK), .D (signal_9038), .Q (signal_9039) ) ;
    buf_clk cell_6903 ( .C (CLK), .D (signal_9046), .Q (signal_9047) ) ;
    buf_clk cell_6911 ( .C (CLK), .D (signal_9054), .Q (signal_9055) ) ;
    buf_clk cell_6919 ( .C (CLK), .D (signal_9062), .Q (signal_9063) ) ;
    buf_clk cell_6927 ( .C (CLK), .D (signal_9070), .Q (signal_9071) ) ;
    buf_clk cell_6935 ( .C (CLK), .D (signal_9078), .Q (signal_9079) ) ;
    buf_clk cell_6943 ( .C (CLK), .D (signal_9086), .Q (signal_9087) ) ;
    buf_clk cell_6951 ( .C (CLK), .D (signal_9094), .Q (signal_9095) ) ;
    buf_clk cell_6959 ( .C (CLK), .D (signal_9102), .Q (signal_9103) ) ;
    buf_clk cell_6967 ( .C (CLK), .D (signal_9110), .Q (signal_9111) ) ;
    buf_clk cell_6975 ( .C (CLK), .D (signal_9118), .Q (signal_9119) ) ;
    buf_clk cell_6983 ( .C (CLK), .D (signal_9126), .Q (signal_9127) ) ;
    buf_clk cell_6991 ( .C (CLK), .D (signal_9134), .Q (signal_9135) ) ;
    buf_clk cell_6999 ( .C (CLK), .D (signal_9142), .Q (signal_9143) ) ;
    buf_clk cell_7007 ( .C (CLK), .D (signal_9150), .Q (signal_9151) ) ;
    buf_clk cell_7015 ( .C (CLK), .D (signal_9158), .Q (signal_9159) ) ;
    buf_clk cell_7023 ( .C (CLK), .D (signal_9166), .Q (signal_9167) ) ;
    buf_clk cell_7031 ( .C (CLK), .D (signal_9174), .Q (signal_9175) ) ;
    buf_clk cell_7039 ( .C (CLK), .D (signal_9182), .Q (signal_9183) ) ;
    buf_clk cell_7047 ( .C (CLK), .D (signal_9190), .Q (signal_9191) ) ;
    buf_clk cell_7055 ( .C (CLK), .D (signal_9198), .Q (signal_9199) ) ;
    buf_clk cell_7063 ( .C (CLK), .D (signal_9206), .Q (signal_9207) ) ;
    buf_clk cell_7071 ( .C (CLK), .D (signal_9214), .Q (signal_9215) ) ;
    buf_clk cell_7079 ( .C (CLK), .D (signal_9222), .Q (signal_9223) ) ;
    buf_clk cell_7087 ( .C (CLK), .D (signal_9230), .Q (signal_9231) ) ;
    buf_clk cell_7095 ( .C (CLK), .D (signal_9238), .Q (signal_9239) ) ;
    buf_clk cell_7103 ( .C (CLK), .D (signal_9246), .Q (signal_9247) ) ;
    buf_clk cell_7111 ( .C (CLK), .D (signal_9254), .Q (signal_9255) ) ;
    buf_clk cell_7119 ( .C (CLK), .D (signal_9262), .Q (signal_9263) ) ;
    buf_clk cell_7127 ( .C (CLK), .D (signal_9270), .Q (signal_9271) ) ;
    buf_clk cell_7135 ( .C (CLK), .D (signal_9278), .Q (signal_9279) ) ;
    buf_clk cell_7143 ( .C (CLK), .D (signal_9286), .Q (signal_9287) ) ;
    buf_clk cell_7151 ( .C (CLK), .D (signal_9294), .Q (signal_9295) ) ;
    buf_clk cell_7159 ( .C (CLK), .D (signal_9302), .Q (signal_9303) ) ;
    buf_clk cell_7167 ( .C (CLK), .D (signal_9310), .Q (signal_9311) ) ;
    buf_clk cell_7175 ( .C (CLK), .D (signal_9318), .Q (signal_9319) ) ;
    buf_clk cell_7183 ( .C (CLK), .D (signal_9326), .Q (signal_9327) ) ;
    buf_clk cell_7191 ( .C (CLK), .D (signal_9334), .Q (signal_9335) ) ;
    buf_clk cell_7199 ( .C (CLK), .D (signal_9342), .Q (signal_9343) ) ;
    buf_clk cell_7207 ( .C (CLK), .D (signal_9350), .Q (signal_9351) ) ;
    buf_clk cell_7215 ( .C (CLK), .D (signal_9358), .Q (signal_9359) ) ;
    buf_clk cell_7223 ( .C (CLK), .D (signal_9366), .Q (signal_9367) ) ;
    buf_clk cell_7231 ( .C (CLK), .D (signal_9374), .Q (signal_9375) ) ;
    buf_clk cell_7239 ( .C (CLK), .D (signal_9382), .Q (signal_9383) ) ;
    buf_clk cell_7247 ( .C (CLK), .D (signal_9390), .Q (signal_9391) ) ;
    buf_clk cell_7255 ( .C (CLK), .D (signal_9398), .Q (signal_9399) ) ;
    buf_clk cell_7263 ( .C (CLK), .D (signal_9406), .Q (signal_9407) ) ;
    buf_clk cell_7271 ( .C (CLK), .D (signal_9414), .Q (signal_9415) ) ;
    buf_clk cell_7279 ( .C (CLK), .D (signal_9422), .Q (signal_9423) ) ;
    buf_clk cell_7287 ( .C (CLK), .D (signal_9430), .Q (signal_9431) ) ;
    buf_clk cell_7295 ( .C (CLK), .D (signal_9438), .Q (signal_9439) ) ;
    buf_clk cell_7303 ( .C (CLK), .D (signal_9446), .Q (signal_9447) ) ;
    buf_clk cell_7311 ( .C (CLK), .D (signal_9454), .Q (signal_9455) ) ;
    buf_clk cell_7319 ( .C (CLK), .D (signal_9462), .Q (signal_9463) ) ;
    buf_clk cell_7327 ( .C (CLK), .D (signal_9470), .Q (signal_9471) ) ;
    buf_clk cell_7335 ( .C (CLK), .D (signal_9478), .Q (signal_9479) ) ;
    buf_clk cell_7343 ( .C (CLK), .D (signal_9486), .Q (signal_9487) ) ;
    buf_clk cell_7351 ( .C (CLK), .D (signal_9494), .Q (signal_9495) ) ;
    buf_clk cell_7359 ( .C (CLK), .D (signal_9502), .Q (signal_9503) ) ;
    buf_clk cell_7367 ( .C (CLK), .D (signal_9510), .Q (signal_9511) ) ;
    buf_clk cell_7375 ( .C (CLK), .D (signal_9518), .Q (signal_9519) ) ;
    buf_clk cell_7383 ( .C (CLK), .D (signal_9526), .Q (signal_9527) ) ;
    buf_clk cell_7391 ( .C (CLK), .D (signal_9534), .Q (signal_9535) ) ;
    buf_clk cell_7399 ( .C (CLK), .D (signal_9542), .Q (signal_9543) ) ;
    buf_clk cell_7407 ( .C (CLK), .D (signal_9550), .Q (signal_9551) ) ;
    buf_clk cell_7415 ( .C (CLK), .D (signal_9558), .Q (signal_9559) ) ;
    buf_clk cell_7423 ( .C (CLK), .D (signal_9566), .Q (signal_9567) ) ;
    buf_clk cell_7431 ( .C (CLK), .D (signal_9574), .Q (signal_9575) ) ;
    buf_clk cell_7439 ( .C (CLK), .D (signal_9582), .Q (signal_9583) ) ;
    buf_clk cell_7447 ( .C (CLK), .D (signal_9590), .Q (signal_9591) ) ;
    buf_clk cell_7455 ( .C (CLK), .D (signal_9598), .Q (signal_9599) ) ;
    buf_clk cell_7463 ( .C (CLK), .D (signal_9606), .Q (signal_9607) ) ;
    buf_clk cell_7471 ( .C (CLK), .D (signal_9614), .Q (signal_9615) ) ;
    buf_clk cell_7479 ( .C (CLK), .D (signal_9622), .Q (signal_9623) ) ;
    buf_clk cell_7487 ( .C (CLK), .D (signal_9630), .Q (signal_9631) ) ;
    buf_clk cell_7495 ( .C (CLK), .D (signal_9638), .Q (signal_9639) ) ;
    buf_clk cell_7503 ( .C (CLK), .D (signal_9646), .Q (signal_9647) ) ;
    buf_clk cell_7511 ( .C (CLK), .D (signal_9654), .Q (signal_9655) ) ;
    buf_clk cell_7519 ( .C (CLK), .D (signal_9662), .Q (signal_9663) ) ;
    buf_clk cell_7527 ( .C (CLK), .D (signal_9670), .Q (signal_9671) ) ;
    buf_clk cell_7535 ( .C (CLK), .D (signal_9678), .Q (signal_9679) ) ;
    buf_clk cell_7543 ( .C (CLK), .D (signal_9686), .Q (signal_9687) ) ;
    buf_clk cell_7551 ( .C (CLK), .D (signal_9694), .Q (signal_9695) ) ;
    buf_clk cell_7565 ( .C (CLK), .D (signal_9708), .Q (signal_9709) ) ;
    buf_clk cell_7573 ( .C (CLK), .D (signal_9716), .Q (signal_9717) ) ;
    buf_clk cell_7599 ( .C (CLK), .D (signal_9742), .Q (signal_9743) ) ;
    buf_clk cell_7615 ( .C (CLK), .D (signal_9758), .Q (signal_9759) ) ;
    buf_clk cell_7631 ( .C (CLK), .D (signal_9774), .Q (signal_9775) ) ;
    buf_clk cell_7647 ( .C (CLK), .D (signal_9790), .Q (signal_9791) ) ;
    buf_clk cell_7663 ( .C (CLK), .D (signal_9806), .Q (signal_9807) ) ;
    buf_clk cell_7679 ( .C (CLK), .D (signal_9822), .Q (signal_9823) ) ;
    buf_clk cell_7695 ( .C (CLK), .D (signal_9838), .Q (signal_9839) ) ;
    buf_clk cell_7711 ( .C (CLK), .D (signal_9854), .Q (signal_9855) ) ;
    buf_clk cell_7727 ( .C (CLK), .D (signal_9870), .Q (signal_9871) ) ;
    buf_clk cell_7743 ( .C (CLK), .D (signal_9886), .Q (signal_9887) ) ;
    buf_clk cell_7751 ( .C (CLK), .D (signal_9894), .Q (signal_9895) ) ;
    buf_clk cell_7759 ( .C (CLK), .D (signal_9902), .Q (signal_9903) ) ;
    buf_clk cell_7767 ( .C (CLK), .D (signal_9910), .Q (signal_9911) ) ;
    buf_clk cell_7775 ( .C (CLK), .D (signal_9918), .Q (signal_9919) ) ;
    buf_clk cell_7783 ( .C (CLK), .D (signal_9926), .Q (signal_9927) ) ;
    buf_clk cell_7791 ( .C (CLK), .D (signal_9934), .Q (signal_9935) ) ;
    buf_clk cell_7799 ( .C (CLK), .D (signal_9942), .Q (signal_9943) ) ;
    buf_clk cell_7807 ( .C (CLK), .D (signal_9950), .Q (signal_9951) ) ;
    buf_clk cell_7815 ( .C (CLK), .D (signal_9958), .Q (signal_9959) ) ;
    buf_clk cell_7823 ( .C (CLK), .D (signal_9966), .Q (signal_9967) ) ;
    buf_clk cell_7831 ( .C (CLK), .D (signal_9974), .Q (signal_9975) ) ;
    buf_clk cell_7839 ( .C (CLK), .D (signal_9982), .Q (signal_9983) ) ;
    buf_clk cell_7847 ( .C (CLK), .D (signal_9990), .Q (signal_9991) ) ;
    buf_clk cell_7855 ( .C (CLK), .D (signal_9998), .Q (signal_9999) ) ;
    buf_clk cell_7863 ( .C (CLK), .D (signal_10006), .Q (signal_10007) ) ;
    buf_clk cell_7871 ( .C (CLK), .D (signal_10014), .Q (signal_10015) ) ;
    buf_clk cell_7879 ( .C (CLK), .D (signal_10022), .Q (signal_10023) ) ;
    buf_clk cell_7887 ( .C (CLK), .D (signal_10030), .Q (signal_10031) ) ;
    buf_clk cell_7895 ( .C (CLK), .D (signal_10038), .Q (signal_10039) ) ;
    buf_clk cell_7903 ( .C (CLK), .D (signal_10046), .Q (signal_10047) ) ;
    buf_clk cell_7911 ( .C (CLK), .D (signal_10054), .Q (signal_10055) ) ;
    buf_clk cell_7919 ( .C (CLK), .D (signal_10062), .Q (signal_10063) ) ;
    buf_clk cell_7927 ( .C (CLK), .D (signal_10070), .Q (signal_10071) ) ;
    buf_clk cell_7935 ( .C (CLK), .D (signal_10078), .Q (signal_10079) ) ;
    buf_clk cell_7951 ( .C (CLK), .D (signal_10094), .Q (signal_10095) ) ;

    /* cells in depth 11 */
    buf_clk cell_3276 ( .C (CLK), .D (signal_5419), .Q (signal_5420) ) ;
    buf_clk cell_3280 ( .C (CLK), .D (signal_5423), .Q (signal_5424) ) ;
    buf_clk cell_3282 ( .C (CLK), .D (signal_1722), .Q (signal_5426) ) ;
    buf_clk cell_3284 ( .C (CLK), .D (signal_2724), .Q (signal_5428) ) ;
    buf_clk cell_3288 ( .C (CLK), .D (signal_5431), .Q (signal_5432) ) ;
    buf_clk cell_3292 ( .C (CLK), .D (signal_5435), .Q (signal_5436) ) ;
    buf_clk cell_3294 ( .C (CLK), .D (signal_1723), .Q (signal_5438) ) ;
    buf_clk cell_3296 ( .C (CLK), .D (signal_2757), .Q (signal_5440) ) ;
    buf_clk cell_3302 ( .C (CLK), .D (signal_5445), .Q (signal_5446) ) ;
    buf_clk cell_3308 ( .C (CLK), .D (signal_5451), .Q (signal_5452) ) ;
    buf_clk cell_3310 ( .C (CLK), .D (signal_1731), .Q (signal_5454) ) ;
    buf_clk cell_3312 ( .C (CLK), .D (signal_2765), .Q (signal_5456) ) ;
    buf_clk cell_3314 ( .C (CLK), .D (signal_1733), .Q (signal_5458) ) ;
    buf_clk cell_3316 ( .C (CLK), .D (signal_2767), .Q (signal_5460) ) ;
    buf_clk cell_3324 ( .C (CLK), .D (signal_5467), .Q (signal_5468) ) ;
    buf_clk cell_3332 ( .C (CLK), .D (signal_5475), .Q (signal_5476) ) ;
    buf_clk cell_3334 ( .C (CLK), .D (signal_1736), .Q (signal_5478) ) ;
    buf_clk cell_3336 ( .C (CLK), .D (signal_2770), .Q (signal_5480) ) ;
    buf_clk cell_3342 ( .C (CLK), .D (signal_5485), .Q (signal_5486) ) ;
    buf_clk cell_3348 ( .C (CLK), .D (signal_5491), .Q (signal_5492) ) ;
    buf_clk cell_3350 ( .C (CLK), .D (signal_5291), .Q (signal_5494) ) ;
    buf_clk cell_3352 ( .C (CLK), .D (signal_5293), .Q (signal_5496) ) ;
    buf_clk cell_3360 ( .C (CLK), .D (signal_5503), .Q (signal_5504) ) ;
    buf_clk cell_3368 ( .C (CLK), .D (signal_5511), .Q (signal_5512) ) ;
    buf_clk cell_3370 ( .C (CLK), .D (signal_1745), .Q (signal_5514) ) ;
    buf_clk cell_3372 ( .C (CLK), .D (signal_2779), .Q (signal_5516) ) ;
    buf_clk cell_3374 ( .C (CLK), .D (signal_1746), .Q (signal_5518) ) ;
    buf_clk cell_3376 ( .C (CLK), .D (signal_2780), .Q (signal_5520) ) ;
    buf_clk cell_3378 ( .C (CLK), .D (signal_1749), .Q (signal_5522) ) ;
    buf_clk cell_3380 ( .C (CLK), .D (signal_2783), .Q (signal_5524) ) ;
    buf_clk cell_3382 ( .C (CLK), .D (signal_1752), .Q (signal_5526) ) ;
    buf_clk cell_3384 ( .C (CLK), .D (signal_2786), .Q (signal_5528) ) ;
    buf_clk cell_3386 ( .C (CLK), .D (signal_5363), .Q (signal_5530) ) ;
    buf_clk cell_3388 ( .C (CLK), .D (signal_5365), .Q (signal_5532) ) ;
    buf_clk cell_3390 ( .C (CLK), .D (signal_1753), .Q (signal_5534) ) ;
    buf_clk cell_3392 ( .C (CLK), .D (signal_2787), .Q (signal_5536) ) ;
    buf_clk cell_3394 ( .C (CLK), .D (signal_1754), .Q (signal_5538) ) ;
    buf_clk cell_3396 ( .C (CLK), .D (signal_2788), .Q (signal_5540) ) ;
    buf_clk cell_3400 ( .C (CLK), .D (signal_5543), .Q (signal_5544) ) ;
    buf_clk cell_3404 ( .C (CLK), .D (signal_5547), .Q (signal_5548) ) ;
    buf_clk cell_3408 ( .C (CLK), .D (signal_5551), .Q (signal_5552) ) ;
    buf_clk cell_3412 ( .C (CLK), .D (signal_5555), .Q (signal_5556) ) ;
    buf_clk cell_3414 ( .C (CLK), .D (signal_1759), .Q (signal_5558) ) ;
    buf_clk cell_3416 ( .C (CLK), .D (signal_2729), .Q (signal_5560) ) ;
    buf_clk cell_3418 ( .C (CLK), .D (signal_1760), .Q (signal_5562) ) ;
    buf_clk cell_3420 ( .C (CLK), .D (signal_2730), .Q (signal_5564) ) ;
    buf_clk cell_3422 ( .C (CLK), .D (signal_5315), .Q (signal_5566) ) ;
    buf_clk cell_3424 ( .C (CLK), .D (signal_5317), .Q (signal_5568) ) ;
    buf_clk cell_3426 ( .C (CLK), .D (signal_1767), .Q (signal_5570) ) ;
    buf_clk cell_3428 ( .C (CLK), .D (signal_2733), .Q (signal_5572) ) ;
    buf_clk cell_3430 ( .C (CLK), .D (signal_1770), .Q (signal_5574) ) ;
    buf_clk cell_3432 ( .C (CLK), .D (signal_2795), .Q (signal_5576) ) ;
    buf_clk cell_3434 ( .C (CLK), .D (signal_1771), .Q (signal_5578) ) ;
    buf_clk cell_3436 ( .C (CLK), .D (signal_2796), .Q (signal_5580) ) ;
    buf_clk cell_3440 ( .C (CLK), .D (signal_5583), .Q (signal_5584) ) ;
    buf_clk cell_3456 ( .C (CLK), .D (signal_5599), .Q (signal_5600) ) ;
    buf_clk cell_3472 ( .C (CLK), .D (signal_5615), .Q (signal_5616) ) ;
    buf_clk cell_3480 ( .C (CLK), .D (signal_5623), .Q (signal_5624) ) ;
    buf_clk cell_3496 ( .C (CLK), .D (signal_5639), .Q (signal_5640) ) ;
    buf_clk cell_3512 ( .C (CLK), .D (signal_5655), .Q (signal_5656) ) ;
    buf_clk cell_3520 ( .C (CLK), .D (signal_5663), .Q (signal_5664) ) ;
    buf_clk cell_3536 ( .C (CLK), .D (signal_5679), .Q (signal_5680) ) ;
    buf_clk cell_3552 ( .C (CLK), .D (signal_5695), .Q (signal_5696) ) ;
    buf_clk cell_3568 ( .C (CLK), .D (signal_5711), .Q (signal_5712) ) ;
    buf_clk cell_3584 ( .C (CLK), .D (signal_5727), .Q (signal_5728) ) ;
    buf_clk cell_3598 ( .C (CLK), .D (signal_5359), .Q (signal_5742) ) ;
    buf_clk cell_3604 ( .C (CLK), .D (signal_5361), .Q (signal_5748) ) ;
    buf_clk cell_3610 ( .C (CLK), .D (signal_5383), .Q (signal_5754) ) ;
    buf_clk cell_3616 ( .C (CLK), .D (signal_5385), .Q (signal_5760) ) ;
    buf_clk cell_3622 ( .C (CLK), .D (signal_5377), .Q (signal_5766) ) ;
    buf_clk cell_3628 ( .C (CLK), .D (signal_5381), .Q (signal_5772) ) ;
    buf_clk cell_3644 ( .C (CLK), .D (signal_5787), .Q (signal_5788) ) ;
    buf_clk cell_3660 ( .C (CLK), .D (signal_5803), .Q (signal_5804) ) ;
    buf_clk cell_3676 ( .C (CLK), .D (signal_5819), .Q (signal_5820) ) ;
    buf_clk cell_3692 ( .C (CLK), .D (signal_5835), .Q (signal_5836) ) ;
    buf_clk cell_3708 ( .C (CLK), .D (signal_5851), .Q (signal_5852) ) ;
    buf_clk cell_3724 ( .C (CLK), .D (signal_5867), .Q (signal_5868) ) ;
    buf_clk cell_3740 ( .C (CLK), .D (signal_5883), .Q (signal_5884) ) ;
    buf_clk cell_3756 ( .C (CLK), .D (signal_5899), .Q (signal_5900) ) ;
    buf_clk cell_3772 ( .C (CLK), .D (signal_5915), .Q (signal_5916) ) ;
    buf_clk cell_3788 ( .C (CLK), .D (signal_5931), .Q (signal_5932) ) ;
    buf_clk cell_3804 ( .C (CLK), .D (signal_5947), .Q (signal_5948) ) ;
    buf_clk cell_3812 ( .C (CLK), .D (signal_5955), .Q (signal_5956) ) ;
    buf_clk cell_3818 ( .C (CLK), .D (signal_5275), .Q (signal_5962) ) ;
    buf_clk cell_3824 ( .C (CLK), .D (signal_5277), .Q (signal_5968) ) ;
    buf_clk cell_3832 ( .C (CLK), .D (signal_5975), .Q (signal_5976) ) ;
    buf_clk cell_3840 ( .C (CLK), .D (signal_5983), .Q (signal_5984) ) ;
    buf_clk cell_3848 ( .C (CLK), .D (signal_5991), .Q (signal_5992) ) ;
    buf_clk cell_3856 ( .C (CLK), .D (signal_5999), .Q (signal_6000) ) ;
    buf_clk cell_3872 ( .C (CLK), .D (signal_6015), .Q (signal_6016) ) ;
    buf_clk cell_3880 ( .C (CLK), .D (signal_6023), .Q (signal_6024) ) ;
    buf_clk cell_3896 ( .C (CLK), .D (signal_6039), .Q (signal_6040) ) ;
    buf_clk cell_3912 ( .C (CLK), .D (signal_6055), .Q (signal_6056) ) ;
    buf_clk cell_3928 ( .C (CLK), .D (signal_6071), .Q (signal_6072) ) ;
    buf_clk cell_3944 ( .C (CLK), .D (signal_6087), .Q (signal_6088) ) ;
    buf_clk cell_3960 ( .C (CLK), .D (signal_6103), .Q (signal_6104) ) ;
    buf_clk cell_3976 ( .C (CLK), .D (signal_6119), .Q (signal_6120) ) ;
    buf_clk cell_3992 ( .C (CLK), .D (signal_6135), .Q (signal_6136) ) ;
    buf_clk cell_4008 ( .C (CLK), .D (signal_6151), .Q (signal_6152) ) ;
    buf_clk cell_4024 ( .C (CLK), .D (signal_6167), .Q (signal_6168) ) ;
    buf_clk cell_4040 ( .C (CLK), .D (signal_6183), .Q (signal_6184) ) ;
    buf_clk cell_4056 ( .C (CLK), .D (signal_6199), .Q (signal_6200) ) ;
    buf_clk cell_4072 ( .C (CLK), .D (signal_6215), .Q (signal_6216) ) ;
    buf_clk cell_4088 ( .C (CLK), .D (signal_6231), .Q (signal_6232) ) ;
    buf_clk cell_4104 ( .C (CLK), .D (signal_6247), .Q (signal_6248) ) ;
    buf_clk cell_4114 ( .C (CLK), .D (signal_6257), .Q (signal_6258) ) ;
    buf_clk cell_4124 ( .C (CLK), .D (signal_6267), .Q (signal_6268) ) ;
    buf_clk cell_4130 ( .C (CLK), .D (signal_5287), .Q (signal_6274) ) ;
    buf_clk cell_4136 ( .C (CLK), .D (signal_5289), .Q (signal_6280) ) ;
    buf_clk cell_4144 ( .C (CLK), .D (signal_6287), .Q (signal_6288) ) ;
    buf_clk cell_4152 ( .C (CLK), .D (signal_6295), .Q (signal_6296) ) ;
    buf_clk cell_4162 ( .C (CLK), .D (signal_6305), .Q (signal_6306) ) ;
    buf_clk cell_4172 ( .C (CLK), .D (signal_6315), .Q (signal_6316) ) ;
    buf_clk cell_4188 ( .C (CLK), .D (signal_6331), .Q (signal_6332) ) ;
    buf_clk cell_4200 ( .C (CLK), .D (signal_6343), .Q (signal_6344) ) ;
    buf_clk cell_4212 ( .C (CLK), .D (signal_6355), .Q (signal_6356) ) ;
    buf_clk cell_4220 ( .C (CLK), .D (signal_6363), .Q (signal_6364) ) ;
    buf_clk cell_4228 ( .C (CLK), .D (signal_6371), .Q (signal_6372) ) ;
    buf_clk cell_4240 ( .C (CLK), .D (signal_6383), .Q (signal_6384) ) ;
    buf_clk cell_4252 ( .C (CLK), .D (signal_6395), .Q (signal_6396) ) ;
    buf_clk cell_4266 ( .C (CLK), .D (signal_6409), .Q (signal_6410) ) ;
    buf_clk cell_4280 ( .C (CLK), .D (signal_6423), .Q (signal_6424) ) ;
    buf_clk cell_4296 ( .C (CLK), .D (signal_6439), .Q (signal_6440) ) ;
    buf_clk cell_4312 ( .C (CLK), .D (signal_6455), .Q (signal_6456) ) ;
    buf_clk cell_4328 ( .C (CLK), .D (signal_6471), .Q (signal_6472) ) ;
    buf_clk cell_4344 ( .C (CLK), .D (signal_6487), .Q (signal_6488) ) ;
    buf_clk cell_4360 ( .C (CLK), .D (signal_6503), .Q (signal_6504) ) ;
    buf_clk cell_4376 ( .C (CLK), .D (signal_6519), .Q (signal_6520) ) ;
    buf_clk cell_4392 ( .C (CLK), .D (signal_6535), .Q (signal_6536) ) ;
    buf_clk cell_4408 ( .C (CLK), .D (signal_6551), .Q (signal_6552) ) ;
    buf_clk cell_4424 ( .C (CLK), .D (signal_6567), .Q (signal_6568) ) ;
    buf_clk cell_4440 ( .C (CLK), .D (signal_6583), .Q (signal_6584) ) ;
    buf_clk cell_4456 ( .C (CLK), .D (signal_6599), .Q (signal_6600) ) ;
    buf_clk cell_4472 ( .C (CLK), .D (signal_6615), .Q (signal_6616) ) ;
    buf_clk cell_4488 ( .C (CLK), .D (signal_6631), .Q (signal_6632) ) ;
    buf_clk cell_4504 ( .C (CLK), .D (signal_6647), .Q (signal_6648) ) ;
    buf_clk cell_4520 ( .C (CLK), .D (signal_6663), .Q (signal_6664) ) ;
    buf_clk cell_4536 ( .C (CLK), .D (signal_6679), .Q (signal_6680) ) ;
    buf_clk cell_4546 ( .C (CLK), .D (signal_6689), .Q (signal_6690) ) ;
    buf_clk cell_4556 ( .C (CLK), .D (signal_6699), .Q (signal_6700) ) ;
    buf_clk cell_4564 ( .C (CLK), .D (signal_6707), .Q (signal_6708) ) ;
    buf_clk cell_4572 ( .C (CLK), .D (signal_6715), .Q (signal_6716) ) ;
    buf_clk cell_4584 ( .C (CLK), .D (signal_6727), .Q (signal_6728) ) ;
    buf_clk cell_4596 ( .C (CLK), .D (signal_6739), .Q (signal_6740) ) ;
    buf_clk cell_4610 ( .C (CLK), .D (signal_6753), .Q (signal_6754) ) ;
    buf_clk cell_4624 ( .C (CLK), .D (signal_6767), .Q (signal_6768) ) ;
    buf_clk cell_4640 ( .C (CLK), .D (signal_6783), .Q (signal_6784) ) ;
    buf_clk cell_4656 ( .C (CLK), .D (signal_6799), .Q (signal_6800) ) ;
    buf_clk cell_4662 ( .C (CLK), .D (signal_5335), .Q (signal_6806) ) ;
    buf_clk cell_4668 ( .C (CLK), .D (signal_5337), .Q (signal_6812) ) ;
    buf_clk cell_4676 ( .C (CLK), .D (signal_6819), .Q (signal_6820) ) ;
    buf_clk cell_4684 ( .C (CLK), .D (signal_6827), .Q (signal_6828) ) ;
    buf_clk cell_4694 ( .C (CLK), .D (signal_6837), .Q (signal_6838) ) ;
    buf_clk cell_4704 ( .C (CLK), .D (signal_6847), .Q (signal_6848) ) ;
    buf_clk cell_4716 ( .C (CLK), .D (signal_6859), .Q (signal_6860) ) ;
    buf_clk cell_4728 ( .C (CLK), .D (signal_6871), .Q (signal_6872) ) ;
    buf_clk cell_4736 ( .C (CLK), .D (signal_6879), .Q (signal_6880) ) ;
    buf_clk cell_4752 ( .C (CLK), .D (signal_6895), .Q (signal_6896) ) ;
    buf_clk cell_4768 ( .C (CLK), .D (signal_6911), .Q (signal_6912) ) ;
    buf_clk cell_4784 ( .C (CLK), .D (signal_6927), .Q (signal_6928) ) ;
    buf_clk cell_4800 ( .C (CLK), .D (signal_6943), .Q (signal_6944) ) ;
    buf_clk cell_4816 ( .C (CLK), .D (signal_6959), .Q (signal_6960) ) ;
    buf_clk cell_4832 ( .C (CLK), .D (signal_6975), .Q (signal_6976) ) ;
    buf_clk cell_4848 ( .C (CLK), .D (signal_6991), .Q (signal_6992) ) ;
    buf_clk cell_4864 ( .C (CLK), .D (signal_7007), .Q (signal_7008) ) ;
    buf_clk cell_4880 ( .C (CLK), .D (signal_7023), .Q (signal_7024) ) ;
    buf_clk cell_4896 ( .C (CLK), .D (signal_7039), .Q (signal_7040) ) ;
    buf_clk cell_4912 ( .C (CLK), .D (signal_7055), .Q (signal_7056) ) ;
    buf_clk cell_4928 ( .C (CLK), .D (signal_7071), .Q (signal_7072) ) ;
    buf_clk cell_4944 ( .C (CLK), .D (signal_7087), .Q (signal_7088) ) ;
    buf_clk cell_4960 ( .C (CLK), .D (signal_7103), .Q (signal_7104) ) ;
    buf_clk cell_4976 ( .C (CLK), .D (signal_7119), .Q (signal_7120) ) ;
    buf_clk cell_4992 ( .C (CLK), .D (signal_7135), .Q (signal_7136) ) ;
    buf_clk cell_5008 ( .C (CLK), .D (signal_7151), .Q (signal_7152) ) ;
    buf_clk cell_5024 ( .C (CLK), .D (signal_7167), .Q (signal_7168) ) ;
    buf_clk cell_5040 ( .C (CLK), .D (signal_7183), .Q (signal_7184) ) ;
    buf_clk cell_5056 ( .C (CLK), .D (signal_7199), .Q (signal_7200) ) ;
    buf_clk cell_5072 ( .C (CLK), .D (signal_7215), .Q (signal_7216) ) ;
    buf_clk cell_5088 ( .C (CLK), .D (signal_7231), .Q (signal_7232) ) ;
    buf_clk cell_5104 ( .C (CLK), .D (signal_7247), .Q (signal_7248) ) ;
    buf_clk cell_5120 ( .C (CLK), .D (signal_7263), .Q (signal_7264) ) ;
    buf_clk cell_5136 ( .C (CLK), .D (signal_7279), .Q (signal_7280) ) ;
    buf_clk cell_5152 ( .C (CLK), .D (signal_7295), .Q (signal_7296) ) ;
    buf_clk cell_5168 ( .C (CLK), .D (signal_7311), .Q (signal_7312) ) ;
    buf_clk cell_5184 ( .C (CLK), .D (signal_7327), .Q (signal_7328) ) ;
    buf_clk cell_5200 ( .C (CLK), .D (signal_7343), .Q (signal_7344) ) ;
    buf_clk cell_5216 ( .C (CLK), .D (signal_7359), .Q (signal_7360) ) ;
    buf_clk cell_5232 ( .C (CLK), .D (signal_7375), .Q (signal_7376) ) ;
    buf_clk cell_5248 ( .C (CLK), .D (signal_7391), .Q (signal_7392) ) ;
    buf_clk cell_5264 ( .C (CLK), .D (signal_7407), .Q (signal_7408) ) ;
    buf_clk cell_5280 ( .C (CLK), .D (signal_7423), .Q (signal_7424) ) ;
    buf_clk cell_5296 ( .C (CLK), .D (signal_7439), .Q (signal_7440) ) ;
    buf_clk cell_5312 ( .C (CLK), .D (signal_7455), .Q (signal_7456) ) ;
    buf_clk cell_5328 ( .C (CLK), .D (signal_7471), .Q (signal_7472) ) ;
    buf_clk cell_5344 ( .C (CLK), .D (signal_7487), .Q (signal_7488) ) ;
    buf_clk cell_5360 ( .C (CLK), .D (signal_7503), .Q (signal_7504) ) ;
    buf_clk cell_5376 ( .C (CLK), .D (signal_7519), .Q (signal_7520) ) ;
    buf_clk cell_5392 ( .C (CLK), .D (signal_7535), .Q (signal_7536) ) ;
    buf_clk cell_5408 ( .C (CLK), .D (signal_7551), .Q (signal_7552) ) ;
    buf_clk cell_5424 ( .C (CLK), .D (signal_7567), .Q (signal_7568) ) ;
    buf_clk cell_5440 ( .C (CLK), .D (signal_7583), .Q (signal_7584) ) ;
    buf_clk cell_5456 ( .C (CLK), .D (signal_7599), .Q (signal_7600) ) ;
    buf_clk cell_5472 ( .C (CLK), .D (signal_7615), .Q (signal_7616) ) ;
    buf_clk cell_5488 ( .C (CLK), .D (signal_7631), .Q (signal_7632) ) ;
    buf_clk cell_5504 ( .C (CLK), .D (signal_7647), .Q (signal_7648) ) ;
    buf_clk cell_5520 ( .C (CLK), .D (signal_7663), .Q (signal_7664) ) ;
    buf_clk cell_5536 ( .C (CLK), .D (signal_7679), .Q (signal_7680) ) ;
    buf_clk cell_5552 ( .C (CLK), .D (signal_7695), .Q (signal_7696) ) ;
    buf_clk cell_5568 ( .C (CLK), .D (signal_7711), .Q (signal_7712) ) ;
    buf_clk cell_5584 ( .C (CLK), .D (signal_7727), .Q (signal_7728) ) ;
    buf_clk cell_5600 ( .C (CLK), .D (signal_7743), .Q (signal_7744) ) ;
    buf_clk cell_5616 ( .C (CLK), .D (signal_7759), .Q (signal_7760) ) ;
    buf_clk cell_5632 ( .C (CLK), .D (signal_7775), .Q (signal_7776) ) ;
    buf_clk cell_5648 ( .C (CLK), .D (signal_7791), .Q (signal_7792) ) ;
    buf_clk cell_5664 ( .C (CLK), .D (signal_7807), .Q (signal_7808) ) ;
    buf_clk cell_5680 ( .C (CLK), .D (signal_7823), .Q (signal_7824) ) ;
    buf_clk cell_5696 ( .C (CLK), .D (signal_7839), .Q (signal_7840) ) ;
    buf_clk cell_5712 ( .C (CLK), .D (signal_7855), .Q (signal_7856) ) ;
    buf_clk cell_5728 ( .C (CLK), .D (signal_7871), .Q (signal_7872) ) ;
    buf_clk cell_5744 ( .C (CLK), .D (signal_7887), .Q (signal_7888) ) ;
    buf_clk cell_5760 ( .C (CLK), .D (signal_7903), .Q (signal_7904) ) ;
    buf_clk cell_5776 ( .C (CLK), .D (signal_7919), .Q (signal_7920) ) ;
    buf_clk cell_5792 ( .C (CLK), .D (signal_7935), .Q (signal_7936) ) ;
    buf_clk cell_5808 ( .C (CLK), .D (signal_7951), .Q (signal_7952) ) ;
    buf_clk cell_5824 ( .C (CLK), .D (signal_7967), .Q (signal_7968) ) ;
    buf_clk cell_5840 ( .C (CLK), .D (signal_7983), .Q (signal_7984) ) ;
    buf_clk cell_5856 ( .C (CLK), .D (signal_7999), .Q (signal_8000) ) ;
    buf_clk cell_5872 ( .C (CLK), .D (signal_8015), .Q (signal_8016) ) ;
    buf_clk cell_5888 ( .C (CLK), .D (signal_8031), .Q (signal_8032) ) ;
    buf_clk cell_5904 ( .C (CLK), .D (signal_8047), .Q (signal_8048) ) ;
    buf_clk cell_5920 ( .C (CLK), .D (signal_8063), .Q (signal_8064) ) ;
    buf_clk cell_5936 ( .C (CLK), .D (signal_8079), .Q (signal_8080) ) ;
    buf_clk cell_5952 ( .C (CLK), .D (signal_8095), .Q (signal_8096) ) ;
    buf_clk cell_5968 ( .C (CLK), .D (signal_8111), .Q (signal_8112) ) ;
    buf_clk cell_5984 ( .C (CLK), .D (signal_8127), .Q (signal_8128) ) ;
    buf_clk cell_6000 ( .C (CLK), .D (signal_8143), .Q (signal_8144) ) ;
    buf_clk cell_6016 ( .C (CLK), .D (signal_8159), .Q (signal_8160) ) ;
    buf_clk cell_6032 ( .C (CLK), .D (signal_8175), .Q (signal_8176) ) ;
    buf_clk cell_6048 ( .C (CLK), .D (signal_8191), .Q (signal_8192) ) ;
    buf_clk cell_6064 ( .C (CLK), .D (signal_8207), .Q (signal_8208) ) ;
    buf_clk cell_6080 ( .C (CLK), .D (signal_8223), .Q (signal_8224) ) ;
    buf_clk cell_6096 ( .C (CLK), .D (signal_8239), .Q (signal_8240) ) ;
    buf_clk cell_6112 ( .C (CLK), .D (signal_8255), .Q (signal_8256) ) ;
    buf_clk cell_6128 ( .C (CLK), .D (signal_8271), .Q (signal_8272) ) ;
    buf_clk cell_6144 ( .C (CLK), .D (signal_8287), .Q (signal_8288) ) ;
    buf_clk cell_6160 ( .C (CLK), .D (signal_8303), .Q (signal_8304) ) ;
    buf_clk cell_6176 ( .C (CLK), .D (signal_8319), .Q (signal_8320) ) ;
    buf_clk cell_6192 ( .C (CLK), .D (signal_8335), .Q (signal_8336) ) ;
    buf_clk cell_6208 ( .C (CLK), .D (signal_8351), .Q (signal_8352) ) ;
    buf_clk cell_6224 ( .C (CLK), .D (signal_8367), .Q (signal_8368) ) ;
    buf_clk cell_6240 ( .C (CLK), .D (signal_8383), .Q (signal_8384) ) ;
    buf_clk cell_6256 ( .C (CLK), .D (signal_8399), .Q (signal_8400) ) ;
    buf_clk cell_6272 ( .C (CLK), .D (signal_8415), .Q (signal_8416) ) ;
    buf_clk cell_6288 ( .C (CLK), .D (signal_8431), .Q (signal_8432) ) ;
    buf_clk cell_6304 ( .C (CLK), .D (signal_8447), .Q (signal_8448) ) ;
    buf_clk cell_6320 ( .C (CLK), .D (signal_8463), .Q (signal_8464) ) ;
    buf_clk cell_6336 ( .C (CLK), .D (signal_8479), .Q (signal_8480) ) ;
    buf_clk cell_6352 ( .C (CLK), .D (signal_8495), .Q (signal_8496) ) ;
    buf_clk cell_6368 ( .C (CLK), .D (signal_8511), .Q (signal_8512) ) ;
    buf_clk cell_6384 ( .C (CLK), .D (signal_8527), .Q (signal_8528) ) ;
    buf_clk cell_6400 ( .C (CLK), .D (signal_8543), .Q (signal_8544) ) ;
    buf_clk cell_6408 ( .C (CLK), .D (signal_8551), .Q (signal_8552) ) ;
    buf_clk cell_6416 ( .C (CLK), .D (signal_8559), .Q (signal_8560) ) ;
    buf_clk cell_6424 ( .C (CLK), .D (signal_8567), .Q (signal_8568) ) ;
    buf_clk cell_6432 ( .C (CLK), .D (signal_8575), .Q (signal_8576) ) ;
    buf_clk cell_6440 ( .C (CLK), .D (signal_8583), .Q (signal_8584) ) ;
    buf_clk cell_6448 ( .C (CLK), .D (signal_8591), .Q (signal_8592) ) ;
    buf_clk cell_6456 ( .C (CLK), .D (signal_8599), .Q (signal_8600) ) ;
    buf_clk cell_6464 ( .C (CLK), .D (signal_8607), .Q (signal_8608) ) ;
    buf_clk cell_6472 ( .C (CLK), .D (signal_8615), .Q (signal_8616) ) ;
    buf_clk cell_6480 ( .C (CLK), .D (signal_8623), .Q (signal_8624) ) ;
    buf_clk cell_6488 ( .C (CLK), .D (signal_8631), .Q (signal_8632) ) ;
    buf_clk cell_6496 ( .C (CLK), .D (signal_8639), .Q (signal_8640) ) ;
    buf_clk cell_6504 ( .C (CLK), .D (signal_8647), .Q (signal_8648) ) ;
    buf_clk cell_6512 ( .C (CLK), .D (signal_8655), .Q (signal_8656) ) ;
    buf_clk cell_6520 ( .C (CLK), .D (signal_8663), .Q (signal_8664) ) ;
    buf_clk cell_6528 ( .C (CLK), .D (signal_8671), .Q (signal_8672) ) ;
    buf_clk cell_6536 ( .C (CLK), .D (signal_8679), .Q (signal_8680) ) ;
    buf_clk cell_6544 ( .C (CLK), .D (signal_8687), .Q (signal_8688) ) ;
    buf_clk cell_6552 ( .C (CLK), .D (signal_8695), .Q (signal_8696) ) ;
    buf_clk cell_6560 ( .C (CLK), .D (signal_8703), .Q (signal_8704) ) ;
    buf_clk cell_6568 ( .C (CLK), .D (signal_8711), .Q (signal_8712) ) ;
    buf_clk cell_6576 ( .C (CLK), .D (signal_8719), .Q (signal_8720) ) ;
    buf_clk cell_6584 ( .C (CLK), .D (signal_8727), .Q (signal_8728) ) ;
    buf_clk cell_6592 ( .C (CLK), .D (signal_8735), .Q (signal_8736) ) ;
    buf_clk cell_6600 ( .C (CLK), .D (signal_8743), .Q (signal_8744) ) ;
    buf_clk cell_6608 ( .C (CLK), .D (signal_8751), .Q (signal_8752) ) ;
    buf_clk cell_6616 ( .C (CLK), .D (signal_8759), .Q (signal_8760) ) ;
    buf_clk cell_6624 ( .C (CLK), .D (signal_8767), .Q (signal_8768) ) ;
    buf_clk cell_6632 ( .C (CLK), .D (signal_8775), .Q (signal_8776) ) ;
    buf_clk cell_6640 ( .C (CLK), .D (signal_8783), .Q (signal_8784) ) ;
    buf_clk cell_6648 ( .C (CLK), .D (signal_8791), .Q (signal_8792) ) ;
    buf_clk cell_6656 ( .C (CLK), .D (signal_8799), .Q (signal_8800) ) ;
    buf_clk cell_6664 ( .C (CLK), .D (signal_8807), .Q (signal_8808) ) ;
    buf_clk cell_6672 ( .C (CLK), .D (signal_8815), .Q (signal_8816) ) ;
    buf_clk cell_6680 ( .C (CLK), .D (signal_8823), .Q (signal_8824) ) ;
    buf_clk cell_6688 ( .C (CLK), .D (signal_8831), .Q (signal_8832) ) ;
    buf_clk cell_6696 ( .C (CLK), .D (signal_8839), .Q (signal_8840) ) ;
    buf_clk cell_6704 ( .C (CLK), .D (signal_8847), .Q (signal_8848) ) ;
    buf_clk cell_6712 ( .C (CLK), .D (signal_8855), .Q (signal_8856) ) ;
    buf_clk cell_6720 ( .C (CLK), .D (signal_8863), .Q (signal_8864) ) ;
    buf_clk cell_6728 ( .C (CLK), .D (signal_8871), .Q (signal_8872) ) ;
    buf_clk cell_6736 ( .C (CLK), .D (signal_8879), .Q (signal_8880) ) ;
    buf_clk cell_6744 ( .C (CLK), .D (signal_8887), .Q (signal_8888) ) ;
    buf_clk cell_6752 ( .C (CLK), .D (signal_8895), .Q (signal_8896) ) ;
    buf_clk cell_6760 ( .C (CLK), .D (signal_8903), .Q (signal_8904) ) ;
    buf_clk cell_6768 ( .C (CLK), .D (signal_8911), .Q (signal_8912) ) ;
    buf_clk cell_6776 ( .C (CLK), .D (signal_8919), .Q (signal_8920) ) ;
    buf_clk cell_6784 ( .C (CLK), .D (signal_8927), .Q (signal_8928) ) ;
    buf_clk cell_6792 ( .C (CLK), .D (signal_8935), .Q (signal_8936) ) ;
    buf_clk cell_6800 ( .C (CLK), .D (signal_8943), .Q (signal_8944) ) ;
    buf_clk cell_6808 ( .C (CLK), .D (signal_8951), .Q (signal_8952) ) ;
    buf_clk cell_6816 ( .C (CLK), .D (signal_8959), .Q (signal_8960) ) ;
    buf_clk cell_6824 ( .C (CLK), .D (signal_8967), .Q (signal_8968) ) ;
    buf_clk cell_6832 ( .C (CLK), .D (signal_8975), .Q (signal_8976) ) ;
    buf_clk cell_6840 ( .C (CLK), .D (signal_8983), .Q (signal_8984) ) ;
    buf_clk cell_6848 ( .C (CLK), .D (signal_8991), .Q (signal_8992) ) ;
    buf_clk cell_6856 ( .C (CLK), .D (signal_8999), .Q (signal_9000) ) ;
    buf_clk cell_6864 ( .C (CLK), .D (signal_9007), .Q (signal_9008) ) ;
    buf_clk cell_6872 ( .C (CLK), .D (signal_9015), .Q (signal_9016) ) ;
    buf_clk cell_6880 ( .C (CLK), .D (signal_9023), .Q (signal_9024) ) ;
    buf_clk cell_6888 ( .C (CLK), .D (signal_9031), .Q (signal_9032) ) ;
    buf_clk cell_6896 ( .C (CLK), .D (signal_9039), .Q (signal_9040) ) ;
    buf_clk cell_6904 ( .C (CLK), .D (signal_9047), .Q (signal_9048) ) ;
    buf_clk cell_6912 ( .C (CLK), .D (signal_9055), .Q (signal_9056) ) ;
    buf_clk cell_6920 ( .C (CLK), .D (signal_9063), .Q (signal_9064) ) ;
    buf_clk cell_6928 ( .C (CLK), .D (signal_9071), .Q (signal_9072) ) ;
    buf_clk cell_6936 ( .C (CLK), .D (signal_9079), .Q (signal_9080) ) ;
    buf_clk cell_6944 ( .C (CLK), .D (signal_9087), .Q (signal_9088) ) ;
    buf_clk cell_6952 ( .C (CLK), .D (signal_9095), .Q (signal_9096) ) ;
    buf_clk cell_6960 ( .C (CLK), .D (signal_9103), .Q (signal_9104) ) ;
    buf_clk cell_6968 ( .C (CLK), .D (signal_9111), .Q (signal_9112) ) ;
    buf_clk cell_6976 ( .C (CLK), .D (signal_9119), .Q (signal_9120) ) ;
    buf_clk cell_6984 ( .C (CLK), .D (signal_9127), .Q (signal_9128) ) ;
    buf_clk cell_6992 ( .C (CLK), .D (signal_9135), .Q (signal_9136) ) ;
    buf_clk cell_7000 ( .C (CLK), .D (signal_9143), .Q (signal_9144) ) ;
    buf_clk cell_7008 ( .C (CLK), .D (signal_9151), .Q (signal_9152) ) ;
    buf_clk cell_7016 ( .C (CLK), .D (signal_9159), .Q (signal_9160) ) ;
    buf_clk cell_7024 ( .C (CLK), .D (signal_9167), .Q (signal_9168) ) ;
    buf_clk cell_7032 ( .C (CLK), .D (signal_9175), .Q (signal_9176) ) ;
    buf_clk cell_7040 ( .C (CLK), .D (signal_9183), .Q (signal_9184) ) ;
    buf_clk cell_7048 ( .C (CLK), .D (signal_9191), .Q (signal_9192) ) ;
    buf_clk cell_7056 ( .C (CLK), .D (signal_9199), .Q (signal_9200) ) ;
    buf_clk cell_7064 ( .C (CLK), .D (signal_9207), .Q (signal_9208) ) ;
    buf_clk cell_7072 ( .C (CLK), .D (signal_9215), .Q (signal_9216) ) ;
    buf_clk cell_7080 ( .C (CLK), .D (signal_9223), .Q (signal_9224) ) ;
    buf_clk cell_7088 ( .C (CLK), .D (signal_9231), .Q (signal_9232) ) ;
    buf_clk cell_7096 ( .C (CLK), .D (signal_9239), .Q (signal_9240) ) ;
    buf_clk cell_7104 ( .C (CLK), .D (signal_9247), .Q (signal_9248) ) ;
    buf_clk cell_7112 ( .C (CLK), .D (signal_9255), .Q (signal_9256) ) ;
    buf_clk cell_7120 ( .C (CLK), .D (signal_9263), .Q (signal_9264) ) ;
    buf_clk cell_7128 ( .C (CLK), .D (signal_9271), .Q (signal_9272) ) ;
    buf_clk cell_7136 ( .C (CLK), .D (signal_9279), .Q (signal_9280) ) ;
    buf_clk cell_7144 ( .C (CLK), .D (signal_9287), .Q (signal_9288) ) ;
    buf_clk cell_7152 ( .C (CLK), .D (signal_9295), .Q (signal_9296) ) ;
    buf_clk cell_7160 ( .C (CLK), .D (signal_9303), .Q (signal_9304) ) ;
    buf_clk cell_7168 ( .C (CLK), .D (signal_9311), .Q (signal_9312) ) ;
    buf_clk cell_7176 ( .C (CLK), .D (signal_9319), .Q (signal_9320) ) ;
    buf_clk cell_7184 ( .C (CLK), .D (signal_9327), .Q (signal_9328) ) ;
    buf_clk cell_7192 ( .C (CLK), .D (signal_9335), .Q (signal_9336) ) ;
    buf_clk cell_7200 ( .C (CLK), .D (signal_9343), .Q (signal_9344) ) ;
    buf_clk cell_7208 ( .C (CLK), .D (signal_9351), .Q (signal_9352) ) ;
    buf_clk cell_7216 ( .C (CLK), .D (signal_9359), .Q (signal_9360) ) ;
    buf_clk cell_7224 ( .C (CLK), .D (signal_9367), .Q (signal_9368) ) ;
    buf_clk cell_7232 ( .C (CLK), .D (signal_9375), .Q (signal_9376) ) ;
    buf_clk cell_7240 ( .C (CLK), .D (signal_9383), .Q (signal_9384) ) ;
    buf_clk cell_7248 ( .C (CLK), .D (signal_9391), .Q (signal_9392) ) ;
    buf_clk cell_7256 ( .C (CLK), .D (signal_9399), .Q (signal_9400) ) ;
    buf_clk cell_7264 ( .C (CLK), .D (signal_9407), .Q (signal_9408) ) ;
    buf_clk cell_7272 ( .C (CLK), .D (signal_9415), .Q (signal_9416) ) ;
    buf_clk cell_7280 ( .C (CLK), .D (signal_9423), .Q (signal_9424) ) ;
    buf_clk cell_7288 ( .C (CLK), .D (signal_9431), .Q (signal_9432) ) ;
    buf_clk cell_7296 ( .C (CLK), .D (signal_9439), .Q (signal_9440) ) ;
    buf_clk cell_7304 ( .C (CLK), .D (signal_9447), .Q (signal_9448) ) ;
    buf_clk cell_7312 ( .C (CLK), .D (signal_9455), .Q (signal_9456) ) ;
    buf_clk cell_7320 ( .C (CLK), .D (signal_9463), .Q (signal_9464) ) ;
    buf_clk cell_7328 ( .C (CLK), .D (signal_9471), .Q (signal_9472) ) ;
    buf_clk cell_7336 ( .C (CLK), .D (signal_9479), .Q (signal_9480) ) ;
    buf_clk cell_7344 ( .C (CLK), .D (signal_9487), .Q (signal_9488) ) ;
    buf_clk cell_7352 ( .C (CLK), .D (signal_9495), .Q (signal_9496) ) ;
    buf_clk cell_7360 ( .C (CLK), .D (signal_9503), .Q (signal_9504) ) ;
    buf_clk cell_7368 ( .C (CLK), .D (signal_9511), .Q (signal_9512) ) ;
    buf_clk cell_7376 ( .C (CLK), .D (signal_9519), .Q (signal_9520) ) ;
    buf_clk cell_7384 ( .C (CLK), .D (signal_9527), .Q (signal_9528) ) ;
    buf_clk cell_7392 ( .C (CLK), .D (signal_9535), .Q (signal_9536) ) ;
    buf_clk cell_7400 ( .C (CLK), .D (signal_9543), .Q (signal_9544) ) ;
    buf_clk cell_7408 ( .C (CLK), .D (signal_9551), .Q (signal_9552) ) ;
    buf_clk cell_7416 ( .C (CLK), .D (signal_9559), .Q (signal_9560) ) ;
    buf_clk cell_7424 ( .C (CLK), .D (signal_9567), .Q (signal_9568) ) ;
    buf_clk cell_7432 ( .C (CLK), .D (signal_9575), .Q (signal_9576) ) ;
    buf_clk cell_7440 ( .C (CLK), .D (signal_9583), .Q (signal_9584) ) ;
    buf_clk cell_7448 ( .C (CLK), .D (signal_9591), .Q (signal_9592) ) ;
    buf_clk cell_7456 ( .C (CLK), .D (signal_9599), .Q (signal_9600) ) ;
    buf_clk cell_7464 ( .C (CLK), .D (signal_9607), .Q (signal_9608) ) ;
    buf_clk cell_7472 ( .C (CLK), .D (signal_9615), .Q (signal_9616) ) ;
    buf_clk cell_7480 ( .C (CLK), .D (signal_9623), .Q (signal_9624) ) ;
    buf_clk cell_7488 ( .C (CLK), .D (signal_9631), .Q (signal_9632) ) ;
    buf_clk cell_7496 ( .C (CLK), .D (signal_9639), .Q (signal_9640) ) ;
    buf_clk cell_7504 ( .C (CLK), .D (signal_9647), .Q (signal_9648) ) ;
    buf_clk cell_7512 ( .C (CLK), .D (signal_9655), .Q (signal_9656) ) ;
    buf_clk cell_7520 ( .C (CLK), .D (signal_9663), .Q (signal_9664) ) ;
    buf_clk cell_7528 ( .C (CLK), .D (signal_9671), .Q (signal_9672) ) ;
    buf_clk cell_7536 ( .C (CLK), .D (signal_9679), .Q (signal_9680) ) ;
    buf_clk cell_7544 ( .C (CLK), .D (signal_9687), .Q (signal_9688) ) ;
    buf_clk cell_7552 ( .C (CLK), .D (signal_9695), .Q (signal_9696) ) ;
    buf_clk cell_7566 ( .C (CLK), .D (signal_9709), .Q (signal_9710) ) ;
    buf_clk cell_7574 ( .C (CLK), .D (signal_9717), .Q (signal_9718) ) ;
    buf_clk cell_7578 ( .C (CLK), .D (signal_5355), .Q (signal_9722) ) ;
    buf_clk cell_7582 ( .C (CLK), .D (signal_5357), .Q (signal_9726) ) ;
    buf_clk cell_7600 ( .C (CLK), .D (signal_9743), .Q (signal_9744) ) ;
    buf_clk cell_7616 ( .C (CLK), .D (signal_9759), .Q (signal_9760) ) ;
    buf_clk cell_7632 ( .C (CLK), .D (signal_9775), .Q (signal_9776) ) ;
    buf_clk cell_7648 ( .C (CLK), .D (signal_9791), .Q (signal_9792) ) ;
    buf_clk cell_7664 ( .C (CLK), .D (signal_9807), .Q (signal_9808) ) ;
    buf_clk cell_7680 ( .C (CLK), .D (signal_9823), .Q (signal_9824) ) ;
    buf_clk cell_7696 ( .C (CLK), .D (signal_9839), .Q (signal_9840) ) ;
    buf_clk cell_7712 ( .C (CLK), .D (signal_9855), .Q (signal_9856) ) ;
    buf_clk cell_7728 ( .C (CLK), .D (signal_9871), .Q (signal_9872) ) ;
    buf_clk cell_7744 ( .C (CLK), .D (signal_9887), .Q (signal_9888) ) ;
    buf_clk cell_7752 ( .C (CLK), .D (signal_9895), .Q (signal_9896) ) ;
    buf_clk cell_7760 ( .C (CLK), .D (signal_9903), .Q (signal_9904) ) ;
    buf_clk cell_7768 ( .C (CLK), .D (signal_9911), .Q (signal_9912) ) ;
    buf_clk cell_7776 ( .C (CLK), .D (signal_9919), .Q (signal_9920) ) ;
    buf_clk cell_7784 ( .C (CLK), .D (signal_9927), .Q (signal_9928) ) ;
    buf_clk cell_7792 ( .C (CLK), .D (signal_9935), .Q (signal_9936) ) ;
    buf_clk cell_7800 ( .C (CLK), .D (signal_9943), .Q (signal_9944) ) ;
    buf_clk cell_7808 ( .C (CLK), .D (signal_9951), .Q (signal_9952) ) ;
    buf_clk cell_7816 ( .C (CLK), .D (signal_9959), .Q (signal_9960) ) ;
    buf_clk cell_7824 ( .C (CLK), .D (signal_9967), .Q (signal_9968) ) ;
    buf_clk cell_7832 ( .C (CLK), .D (signal_9975), .Q (signal_9976) ) ;
    buf_clk cell_7840 ( .C (CLK), .D (signal_9983), .Q (signal_9984) ) ;
    buf_clk cell_7848 ( .C (CLK), .D (signal_9991), .Q (signal_9992) ) ;
    buf_clk cell_7856 ( .C (CLK), .D (signal_9999), .Q (signal_10000) ) ;
    buf_clk cell_7864 ( .C (CLK), .D (signal_10007), .Q (signal_10008) ) ;
    buf_clk cell_7872 ( .C (CLK), .D (signal_10015), .Q (signal_10016) ) ;
    buf_clk cell_7880 ( .C (CLK), .D (signal_10023), .Q (signal_10024) ) ;
    buf_clk cell_7888 ( .C (CLK), .D (signal_10031), .Q (signal_10032) ) ;
    buf_clk cell_7896 ( .C (CLK), .D (signal_10039), .Q (signal_10040) ) ;
    buf_clk cell_7904 ( .C (CLK), .D (signal_10047), .Q (signal_10048) ) ;
    buf_clk cell_7912 ( .C (CLK), .D (signal_10055), .Q (signal_10056) ) ;
    buf_clk cell_7920 ( .C (CLK), .D (signal_10063), .Q (signal_10064) ) ;
    buf_clk cell_7928 ( .C (CLK), .D (signal_10071), .Q (signal_10072) ) ;
    buf_clk cell_7936 ( .C (CLK), .D (signal_10079), .Q (signal_10080) ) ;
    buf_clk cell_7952 ( .C (CLK), .D (signal_10095), .Q (signal_10096) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1634 ( .s ({signal_5277, signal_5275}), .b ({signal_2723, signal_1721}), .a ({signal_2722, signal_1720}), .clk (CLK), .r (Fresh[506]), .c ({signal_2803, signal_1778}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1635 ( .s ({signal_5277, signal_5275}), .b ({signal_2723, signal_1721}), .a ({signal_5281, signal_5279}), .clk (CLK), .r (Fresh[507]), .c ({signal_2804, signal_1779}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1636 ( .s ({signal_5277, signal_5275}), .b ({signal_2722, signal_1720}), .a ({signal_5285, signal_5283}), .clk (CLK), .r (Fresh[508]), .c ({signal_2805, signal_1780}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1637 ( .s ({signal_5289, signal_5287}), .b ({signal_2759, signal_1725}), .a ({signal_2758, signal_1724}), .clk (CLK), .r (Fresh[509]), .c ({signal_2838, signal_1781}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1638 ( .s ({signal_5289, signal_5287}), .b ({signal_2761, signal_1727}), .a ({signal_2760, signal_1726}), .clk (CLK), .r (Fresh[510]), .c ({signal_2839, signal_1782}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1639 ( .s ({signal_5289, signal_5287}), .b ({signal_2763, signal_1729}), .a ({signal_2762, signal_1728}), .clk (CLK), .r (Fresh[511]), .c ({signal_2840, signal_1783}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1640 ( .s ({signal_5293, signal_5291}), .b ({signal_2764, signal_1730}), .a ({signal_5297, signal_5295}), .clk (CLK), .r (Fresh[512]), .c ({signal_2841, signal_1784}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1641 ( .s ({signal_5293, signal_5291}), .b ({signal_5301, signal_5299}), .a ({signal_2766, signal_1732}), .clk (CLK), .r (Fresh[513]), .c ({signal_2842, signal_1785}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1642 ( .s ({signal_5305, signal_5303}), .b ({signal_5309, signal_5307}), .a ({signal_2768, signal_1734}), .clk (CLK), .r (Fresh[514]), .c ({signal_2843, signal_1786}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1643 ( .s ({signal_5305, signal_5303}), .b ({signal_5313, signal_5311}), .a ({signal_2769, signal_1735}), .clk (CLK), .r (Fresh[515]), .c ({signal_2844, signal_1787}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1644 ( .s ({signal_5305, signal_5303}), .b ({signal_2768, signal_1734}), .a ({signal_2769, signal_1735}), .clk (CLK), .r (Fresh[516]), .c ({signal_2845, signal_1788}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1645 ( .s ({signal_5317, signal_5315}), .b ({signal_2771, signal_1737}), .a ({signal_5321, signal_5319}), .clk (CLK), .r (Fresh[517]), .c ({signal_2846, signal_1789}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1646 ( .s ({signal_5317, signal_5315}), .b ({signal_5325, signal_5323}), .a ({signal_2772, signal_1738}), .clk (CLK), .r (Fresh[518]), .c ({signal_2847, signal_1790}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1647 ( .s ({signal_5317, signal_5315}), .b ({signal_2773, signal_1739}), .a ({signal_5329, signal_5327}), .clk (CLK), .r (Fresh[519]), .c ({signal_2848, signal_1791}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1648 ( .s ({signal_5317, signal_5315}), .b ({signal_5333, signal_5331}), .a ({signal_2774, signal_1740}), .clk (CLK), .r (Fresh[520]), .c ({signal_2849, signal_1792}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1649 ( .s ({signal_5337, signal_5335}), .b ({signal_2776, signal_1742}), .a ({signal_2775, signal_1741}), .clk (CLK), .r (Fresh[521]), .c ({signal_2850, signal_1793}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1650 ( .s ({signal_5337, signal_5335}), .b ({signal_2778, signal_1744}), .a ({signal_2777, signal_1743}), .clk (CLK), .r (Fresh[522]), .c ({signal_2851, signal_1794}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1651 ( .s ({signal_5353, signal_5345}), .b ({signal_2780, signal_1746}), .a ({signal_2779, signal_1745}), .clk (CLK), .r (Fresh[523]), .c ({signal_2852, signal_1795}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1652 ( .s ({signal_5353, signal_5345}), .b ({signal_2779, signal_1745}), .a ({signal_2780, signal_1746}), .clk (CLK), .r (Fresh[524]), .c ({signal_2853, signal_1796}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1653 ( .s ({signal_5357, signal_5355}), .b ({signal_2782, signal_1748}), .a ({signal_2781, signal_1747}), .clk (CLK), .r (Fresh[525]), .c ({signal_2854, signal_1797}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1654 ( .s ({signal_5357, signal_5355}), .b ({signal_2785, signal_1751}), .a ({signal_2784, signal_1750}), .clk (CLK), .r (Fresh[526]), .c ({signal_2855, signal_1798}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1655 ( .s ({signal_5361, signal_5359}), .b ({signal_2787, signal_1753}), .a ({signal_2788, signal_1754}), .clk (CLK), .r (Fresh[527]), .c ({signal_2856, signal_1799}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1656 ( .s ({signal_5361, signal_5359}), .b ({signal_2788, signal_1754}), .a ({signal_2787, signal_1753}), .clk (CLK), .r (Fresh[528]), .c ({signal_2857, signal_1800}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1657 ( .s ({signal_5365, signal_5363}), .b ({signal_2726, signal_1756}), .a ({signal_2725, signal_1755}), .clk (CLK), .r (Fresh[529]), .c ({signal_2806, signal_1801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1658 ( .s ({signal_5365, signal_5363}), .b ({signal_2727, signal_1757}), .a ({signal_5369, signal_5367}), .clk (CLK), .r (Fresh[530]), .c ({signal_2807, signal_1802}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1659 ( .s ({signal_5365, signal_5363}), .b ({signal_2725, signal_1755}), .a ({signal_2726, signal_1756}), .clk (CLK), .r (Fresh[531]), .c ({signal_2808, signal_1803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1660 ( .s ({signal_5365, signal_5363}), .b ({signal_2728, signal_1758}), .a ({signal_5373, signal_5371}), .clk (CLK), .r (Fresh[532]), .c ({signal_2809, signal_1804}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1661 ( .s ({signal_5381, signal_5377}), .b ({signal_2729, signal_1759}), .a ({signal_2730, signal_1760}), .clk (CLK), .r (Fresh[533]), .c ({signal_2810, signal_1805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1662 ( .s ({signal_5381, signal_5377}), .b ({signal_2730, signal_1760}), .a ({signal_2729, signal_1759}), .clk (CLK), .r (Fresh[534]), .c ({signal_2811, signal_1806}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1663 ( .s ({signal_5385, signal_5383}), .b ({signal_2790, signal_1762}), .a ({signal_2789, signal_1761}), .clk (CLK), .r (Fresh[535]), .c ({signal_2858, signal_1807}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1664 ( .s ({signal_5385, signal_5383}), .b ({signal_2792, signal_1764}), .a ({signal_2791, signal_1763}), .clk (CLK), .r (Fresh[536]), .c ({signal_2859, signal_1808}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1665 ( .s ({signal_5277, signal_5275}), .b ({signal_2732, signal_1766}), .a ({signal_2731, signal_1765}), .clk (CLK), .r (Fresh[537]), .c ({signal_2812, signal_1809}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1666 ( .s ({signal_5277, signal_5275}), .b ({signal_2732, signal_1766}), .a ({signal_5389, signal_5387}), .clk (CLK), .r (Fresh[538]), .c ({signal_2813, signal_1810}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1667 ( .s ({signal_5277, signal_5275}), .b ({signal_2731, signal_1765}), .a ({signal_5393, signal_5391}), .clk (CLK), .r (Fresh[539]), .c ({signal_2814, signal_1811}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1668 ( .s ({signal_5305, signal_5303}), .b ({signal_5397, signal_5395}), .a ({signal_2793, signal_1768}), .clk (CLK), .r (Fresh[540]), .c ({signal_2860, signal_1812}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1669 ( .s ({signal_5305, signal_5303}), .b ({signal_5401, signal_5399}), .a ({signal_2794, signal_1769}), .clk (CLK), .r (Fresh[541]), .c ({signal_2861, signal_1813}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1670 ( .s ({signal_5305, signal_5303}), .b ({signal_2793, signal_1768}), .a ({signal_2794, signal_1769}), .clk (CLK), .r (Fresh[542]), .c ({signal_2862, signal_1814}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1671 ( .s ({signal_5289, signal_5287}), .b ({signal_2798, signal_1773}), .a ({signal_2797, signal_1772}), .clk (CLK), .r (Fresh[543]), .c ({signal_2863, signal_1815}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1672 ( .s ({signal_5289, signal_5287}), .b ({signal_2800, signal_1775}), .a ({signal_2799, signal_1774}), .clk (CLK), .r (Fresh[544]), .c ({signal_2864, signal_1816}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1673 ( .s ({signal_5289, signal_5287}), .b ({signal_2797, signal_1772}), .a ({signal_2798, signal_1773}), .clk (CLK), .r (Fresh[545]), .c ({signal_2865, signal_1817}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1674 ( .s ({signal_5317, signal_5315}), .b ({signal_2801, signal_1776}), .a ({signal_5405, signal_5403}), .clk (CLK), .r (Fresh[546]), .c ({signal_2866, signal_1818}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1675 ( .s ({signal_5317, signal_5315}), .b ({signal_5409, signal_5407}), .a ({signal_2802, signal_1777}), .clk (CLK), .r (Fresh[547]), .c ({signal_2867, signal_1819}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1676 ( .s ({signal_5317, signal_5315}), .b ({signal_2802, signal_1777}), .a ({signal_5413, signal_5411}), .clk (CLK), .r (Fresh[548]), .c ({signal_2868, signal_1820}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1677 ( .s ({signal_5317, signal_5315}), .b ({signal_5417, signal_5415}), .a ({signal_2801, signal_1776}), .clk (CLK), .r (Fresh[549]), .c ({signal_2869, signal_1821}) ) ;
    buf_clk cell_3277 ( .C (CLK), .D (signal_5420), .Q (signal_5421) ) ;
    buf_clk cell_3281 ( .C (CLK), .D (signal_5424), .Q (signal_5425) ) ;
    buf_clk cell_3283 ( .C (CLK), .D (signal_5426), .Q (signal_5427) ) ;
    buf_clk cell_3285 ( .C (CLK), .D (signal_5428), .Q (signal_5429) ) ;
    buf_clk cell_3289 ( .C (CLK), .D (signal_5432), .Q (signal_5433) ) ;
    buf_clk cell_3293 ( .C (CLK), .D (signal_5436), .Q (signal_5437) ) ;
    buf_clk cell_3295 ( .C (CLK), .D (signal_5438), .Q (signal_5439) ) ;
    buf_clk cell_3297 ( .C (CLK), .D (signal_5440), .Q (signal_5441) ) ;
    buf_clk cell_3303 ( .C (CLK), .D (signal_5446), .Q (signal_5447) ) ;
    buf_clk cell_3309 ( .C (CLK), .D (signal_5452), .Q (signal_5453) ) ;
    buf_clk cell_3311 ( .C (CLK), .D (signal_5454), .Q (signal_5455) ) ;
    buf_clk cell_3313 ( .C (CLK), .D (signal_5456), .Q (signal_5457) ) ;
    buf_clk cell_3315 ( .C (CLK), .D (signal_5458), .Q (signal_5459) ) ;
    buf_clk cell_3317 ( .C (CLK), .D (signal_5460), .Q (signal_5461) ) ;
    buf_clk cell_3325 ( .C (CLK), .D (signal_5468), .Q (signal_5469) ) ;
    buf_clk cell_3333 ( .C (CLK), .D (signal_5476), .Q (signal_5477) ) ;
    buf_clk cell_3335 ( .C (CLK), .D (signal_5478), .Q (signal_5479) ) ;
    buf_clk cell_3337 ( .C (CLK), .D (signal_5480), .Q (signal_5481) ) ;
    buf_clk cell_3343 ( .C (CLK), .D (signal_5486), .Q (signal_5487) ) ;
    buf_clk cell_3349 ( .C (CLK), .D (signal_5492), .Q (signal_5493) ) ;
    buf_clk cell_3351 ( .C (CLK), .D (signal_5494), .Q (signal_5495) ) ;
    buf_clk cell_3353 ( .C (CLK), .D (signal_5496), .Q (signal_5497) ) ;
    buf_clk cell_3361 ( .C (CLK), .D (signal_5504), .Q (signal_5505) ) ;
    buf_clk cell_3369 ( .C (CLK), .D (signal_5512), .Q (signal_5513) ) ;
    buf_clk cell_3371 ( .C (CLK), .D (signal_5514), .Q (signal_5515) ) ;
    buf_clk cell_3373 ( .C (CLK), .D (signal_5516), .Q (signal_5517) ) ;
    buf_clk cell_3375 ( .C (CLK), .D (signal_5518), .Q (signal_5519) ) ;
    buf_clk cell_3377 ( .C (CLK), .D (signal_5520), .Q (signal_5521) ) ;
    buf_clk cell_3379 ( .C (CLK), .D (signal_5522), .Q (signal_5523) ) ;
    buf_clk cell_3381 ( .C (CLK), .D (signal_5524), .Q (signal_5525) ) ;
    buf_clk cell_3383 ( .C (CLK), .D (signal_5526), .Q (signal_5527) ) ;
    buf_clk cell_3385 ( .C (CLK), .D (signal_5528), .Q (signal_5529) ) ;
    buf_clk cell_3387 ( .C (CLK), .D (signal_5530), .Q (signal_5531) ) ;
    buf_clk cell_3389 ( .C (CLK), .D (signal_5532), .Q (signal_5533) ) ;
    buf_clk cell_3391 ( .C (CLK), .D (signal_5534), .Q (signal_5535) ) ;
    buf_clk cell_3393 ( .C (CLK), .D (signal_5536), .Q (signal_5537) ) ;
    buf_clk cell_3395 ( .C (CLK), .D (signal_5538), .Q (signal_5539) ) ;
    buf_clk cell_3397 ( .C (CLK), .D (signal_5540), .Q (signal_5541) ) ;
    buf_clk cell_3401 ( .C (CLK), .D (signal_5544), .Q (signal_5545) ) ;
    buf_clk cell_3405 ( .C (CLK), .D (signal_5548), .Q (signal_5549) ) ;
    buf_clk cell_3409 ( .C (CLK), .D (signal_5552), .Q (signal_5553) ) ;
    buf_clk cell_3413 ( .C (CLK), .D (signal_5556), .Q (signal_5557) ) ;
    buf_clk cell_3415 ( .C (CLK), .D (signal_5558), .Q (signal_5559) ) ;
    buf_clk cell_3417 ( .C (CLK), .D (signal_5560), .Q (signal_5561) ) ;
    buf_clk cell_3419 ( .C (CLK), .D (signal_5562), .Q (signal_5563) ) ;
    buf_clk cell_3421 ( .C (CLK), .D (signal_5564), .Q (signal_5565) ) ;
    buf_clk cell_3423 ( .C (CLK), .D (signal_5566), .Q (signal_5567) ) ;
    buf_clk cell_3425 ( .C (CLK), .D (signal_5568), .Q (signal_5569) ) ;
    buf_clk cell_3427 ( .C (CLK), .D (signal_5570), .Q (signal_5571) ) ;
    buf_clk cell_3429 ( .C (CLK), .D (signal_5572), .Q (signal_5573) ) ;
    buf_clk cell_3431 ( .C (CLK), .D (signal_5574), .Q (signal_5575) ) ;
    buf_clk cell_3433 ( .C (CLK), .D (signal_5576), .Q (signal_5577) ) ;
    buf_clk cell_3435 ( .C (CLK), .D (signal_5578), .Q (signal_5579) ) ;
    buf_clk cell_3437 ( .C (CLK), .D (signal_5580), .Q (signal_5581) ) ;
    buf_clk cell_3441 ( .C (CLK), .D (signal_5584), .Q (signal_5585) ) ;
    buf_clk cell_3457 ( .C (CLK), .D (signal_5600), .Q (signal_5601) ) ;
    buf_clk cell_3473 ( .C (CLK), .D (signal_5616), .Q (signal_5617) ) ;
    buf_clk cell_3481 ( .C (CLK), .D (signal_5624), .Q (signal_5625) ) ;
    buf_clk cell_3497 ( .C (CLK), .D (signal_5640), .Q (signal_5641) ) ;
    buf_clk cell_3513 ( .C (CLK), .D (signal_5656), .Q (signal_5657) ) ;
    buf_clk cell_3521 ( .C (CLK), .D (signal_5664), .Q (signal_5665) ) ;
    buf_clk cell_3537 ( .C (CLK), .D (signal_5680), .Q (signal_5681) ) ;
    buf_clk cell_3553 ( .C (CLK), .D (signal_5696), .Q (signal_5697) ) ;
    buf_clk cell_3569 ( .C (CLK), .D (signal_5712), .Q (signal_5713) ) ;
    buf_clk cell_3585 ( .C (CLK), .D (signal_5728), .Q (signal_5729) ) ;
    buf_clk cell_3599 ( .C (CLK), .D (signal_5742), .Q (signal_5743) ) ;
    buf_clk cell_3605 ( .C (CLK), .D (signal_5748), .Q (signal_5749) ) ;
    buf_clk cell_3611 ( .C (CLK), .D (signal_5754), .Q (signal_5755) ) ;
    buf_clk cell_3617 ( .C (CLK), .D (signal_5760), .Q (signal_5761) ) ;
    buf_clk cell_3623 ( .C (CLK), .D (signal_5766), .Q (signal_5767) ) ;
    buf_clk cell_3629 ( .C (CLK), .D (signal_5772), .Q (signal_5773) ) ;
    buf_clk cell_3645 ( .C (CLK), .D (signal_5788), .Q (signal_5789) ) ;
    buf_clk cell_3661 ( .C (CLK), .D (signal_5804), .Q (signal_5805) ) ;
    buf_clk cell_3677 ( .C (CLK), .D (signal_5820), .Q (signal_5821) ) ;
    buf_clk cell_3693 ( .C (CLK), .D (signal_5836), .Q (signal_5837) ) ;
    buf_clk cell_3709 ( .C (CLK), .D (signal_5852), .Q (signal_5853) ) ;
    buf_clk cell_3725 ( .C (CLK), .D (signal_5868), .Q (signal_5869) ) ;
    buf_clk cell_3741 ( .C (CLK), .D (signal_5884), .Q (signal_5885) ) ;
    buf_clk cell_3757 ( .C (CLK), .D (signal_5900), .Q (signal_5901) ) ;
    buf_clk cell_3773 ( .C (CLK), .D (signal_5916), .Q (signal_5917) ) ;
    buf_clk cell_3789 ( .C (CLK), .D (signal_5932), .Q (signal_5933) ) ;
    buf_clk cell_3805 ( .C (CLK), .D (signal_5948), .Q (signal_5949) ) ;
    buf_clk cell_3813 ( .C (CLK), .D (signal_5956), .Q (signal_5957) ) ;
    buf_clk cell_3819 ( .C (CLK), .D (signal_5962), .Q (signal_5963) ) ;
    buf_clk cell_3825 ( .C (CLK), .D (signal_5968), .Q (signal_5969) ) ;
    buf_clk cell_3833 ( .C (CLK), .D (signal_5976), .Q (signal_5977) ) ;
    buf_clk cell_3841 ( .C (CLK), .D (signal_5984), .Q (signal_5985) ) ;
    buf_clk cell_3849 ( .C (CLK), .D (signal_5992), .Q (signal_5993) ) ;
    buf_clk cell_3857 ( .C (CLK), .D (signal_6000), .Q (signal_6001) ) ;
    buf_clk cell_3873 ( .C (CLK), .D (signal_6016), .Q (signal_6017) ) ;
    buf_clk cell_3881 ( .C (CLK), .D (signal_6024), .Q (signal_6025) ) ;
    buf_clk cell_3897 ( .C (CLK), .D (signal_6040), .Q (signal_6041) ) ;
    buf_clk cell_3913 ( .C (CLK), .D (signal_6056), .Q (signal_6057) ) ;
    buf_clk cell_3929 ( .C (CLK), .D (signal_6072), .Q (signal_6073) ) ;
    buf_clk cell_3945 ( .C (CLK), .D (signal_6088), .Q (signal_6089) ) ;
    buf_clk cell_3961 ( .C (CLK), .D (signal_6104), .Q (signal_6105) ) ;
    buf_clk cell_3977 ( .C (CLK), .D (signal_6120), .Q (signal_6121) ) ;
    buf_clk cell_3993 ( .C (CLK), .D (signal_6136), .Q (signal_6137) ) ;
    buf_clk cell_4009 ( .C (CLK), .D (signal_6152), .Q (signal_6153) ) ;
    buf_clk cell_4025 ( .C (CLK), .D (signal_6168), .Q (signal_6169) ) ;
    buf_clk cell_4041 ( .C (CLK), .D (signal_6184), .Q (signal_6185) ) ;
    buf_clk cell_4057 ( .C (CLK), .D (signal_6200), .Q (signal_6201) ) ;
    buf_clk cell_4073 ( .C (CLK), .D (signal_6216), .Q (signal_6217) ) ;
    buf_clk cell_4089 ( .C (CLK), .D (signal_6232), .Q (signal_6233) ) ;
    buf_clk cell_4105 ( .C (CLK), .D (signal_6248), .Q (signal_6249) ) ;
    buf_clk cell_4115 ( .C (CLK), .D (signal_6258), .Q (signal_6259) ) ;
    buf_clk cell_4125 ( .C (CLK), .D (signal_6268), .Q (signal_6269) ) ;
    buf_clk cell_4131 ( .C (CLK), .D (signal_6274), .Q (signal_6275) ) ;
    buf_clk cell_4137 ( .C (CLK), .D (signal_6280), .Q (signal_6281) ) ;
    buf_clk cell_4145 ( .C (CLK), .D (signal_6288), .Q (signal_6289) ) ;
    buf_clk cell_4153 ( .C (CLK), .D (signal_6296), .Q (signal_6297) ) ;
    buf_clk cell_4163 ( .C (CLK), .D (signal_6306), .Q (signal_6307) ) ;
    buf_clk cell_4173 ( .C (CLK), .D (signal_6316), .Q (signal_6317) ) ;
    buf_clk cell_4189 ( .C (CLK), .D (signal_6332), .Q (signal_6333) ) ;
    buf_clk cell_4201 ( .C (CLK), .D (signal_6344), .Q (signal_6345) ) ;
    buf_clk cell_4213 ( .C (CLK), .D (signal_6356), .Q (signal_6357) ) ;
    buf_clk cell_4221 ( .C (CLK), .D (signal_6364), .Q (signal_6365) ) ;
    buf_clk cell_4229 ( .C (CLK), .D (signal_6372), .Q (signal_6373) ) ;
    buf_clk cell_4241 ( .C (CLK), .D (signal_6384), .Q (signal_6385) ) ;
    buf_clk cell_4253 ( .C (CLK), .D (signal_6396), .Q (signal_6397) ) ;
    buf_clk cell_4267 ( .C (CLK), .D (signal_6410), .Q (signal_6411) ) ;
    buf_clk cell_4281 ( .C (CLK), .D (signal_6424), .Q (signal_6425) ) ;
    buf_clk cell_4297 ( .C (CLK), .D (signal_6440), .Q (signal_6441) ) ;
    buf_clk cell_4313 ( .C (CLK), .D (signal_6456), .Q (signal_6457) ) ;
    buf_clk cell_4329 ( .C (CLK), .D (signal_6472), .Q (signal_6473) ) ;
    buf_clk cell_4345 ( .C (CLK), .D (signal_6488), .Q (signal_6489) ) ;
    buf_clk cell_4361 ( .C (CLK), .D (signal_6504), .Q (signal_6505) ) ;
    buf_clk cell_4377 ( .C (CLK), .D (signal_6520), .Q (signal_6521) ) ;
    buf_clk cell_4393 ( .C (CLK), .D (signal_6536), .Q (signal_6537) ) ;
    buf_clk cell_4409 ( .C (CLK), .D (signal_6552), .Q (signal_6553) ) ;
    buf_clk cell_4425 ( .C (CLK), .D (signal_6568), .Q (signal_6569) ) ;
    buf_clk cell_4441 ( .C (CLK), .D (signal_6584), .Q (signal_6585) ) ;
    buf_clk cell_4457 ( .C (CLK), .D (signal_6600), .Q (signal_6601) ) ;
    buf_clk cell_4473 ( .C (CLK), .D (signal_6616), .Q (signal_6617) ) ;
    buf_clk cell_4489 ( .C (CLK), .D (signal_6632), .Q (signal_6633) ) ;
    buf_clk cell_4505 ( .C (CLK), .D (signal_6648), .Q (signal_6649) ) ;
    buf_clk cell_4521 ( .C (CLK), .D (signal_6664), .Q (signal_6665) ) ;
    buf_clk cell_4537 ( .C (CLK), .D (signal_6680), .Q (signal_6681) ) ;
    buf_clk cell_4547 ( .C (CLK), .D (signal_6690), .Q (signal_6691) ) ;
    buf_clk cell_4557 ( .C (CLK), .D (signal_6700), .Q (signal_6701) ) ;
    buf_clk cell_4565 ( .C (CLK), .D (signal_6708), .Q (signal_6709) ) ;
    buf_clk cell_4573 ( .C (CLK), .D (signal_6716), .Q (signal_6717) ) ;
    buf_clk cell_4585 ( .C (CLK), .D (signal_6728), .Q (signal_6729) ) ;
    buf_clk cell_4597 ( .C (CLK), .D (signal_6740), .Q (signal_6741) ) ;
    buf_clk cell_4611 ( .C (CLK), .D (signal_6754), .Q (signal_6755) ) ;
    buf_clk cell_4625 ( .C (CLK), .D (signal_6768), .Q (signal_6769) ) ;
    buf_clk cell_4641 ( .C (CLK), .D (signal_6784), .Q (signal_6785) ) ;
    buf_clk cell_4657 ( .C (CLK), .D (signal_6800), .Q (signal_6801) ) ;
    buf_clk cell_4663 ( .C (CLK), .D (signal_6806), .Q (signal_6807) ) ;
    buf_clk cell_4669 ( .C (CLK), .D (signal_6812), .Q (signal_6813) ) ;
    buf_clk cell_4677 ( .C (CLK), .D (signal_6820), .Q (signal_6821) ) ;
    buf_clk cell_4685 ( .C (CLK), .D (signal_6828), .Q (signal_6829) ) ;
    buf_clk cell_4695 ( .C (CLK), .D (signal_6838), .Q (signal_6839) ) ;
    buf_clk cell_4705 ( .C (CLK), .D (signal_6848), .Q (signal_6849) ) ;
    buf_clk cell_4717 ( .C (CLK), .D (signal_6860), .Q (signal_6861) ) ;
    buf_clk cell_4729 ( .C (CLK), .D (signal_6872), .Q (signal_6873) ) ;
    buf_clk cell_4737 ( .C (CLK), .D (signal_6880), .Q (signal_6881) ) ;
    buf_clk cell_4753 ( .C (CLK), .D (signal_6896), .Q (signal_6897) ) ;
    buf_clk cell_4769 ( .C (CLK), .D (signal_6912), .Q (signal_6913) ) ;
    buf_clk cell_4785 ( .C (CLK), .D (signal_6928), .Q (signal_6929) ) ;
    buf_clk cell_4801 ( .C (CLK), .D (signal_6944), .Q (signal_6945) ) ;
    buf_clk cell_4817 ( .C (CLK), .D (signal_6960), .Q (signal_6961) ) ;
    buf_clk cell_4833 ( .C (CLK), .D (signal_6976), .Q (signal_6977) ) ;
    buf_clk cell_4849 ( .C (CLK), .D (signal_6992), .Q (signal_6993) ) ;
    buf_clk cell_4865 ( .C (CLK), .D (signal_7008), .Q (signal_7009) ) ;
    buf_clk cell_4881 ( .C (CLK), .D (signal_7024), .Q (signal_7025) ) ;
    buf_clk cell_4897 ( .C (CLK), .D (signal_7040), .Q (signal_7041) ) ;
    buf_clk cell_4913 ( .C (CLK), .D (signal_7056), .Q (signal_7057) ) ;
    buf_clk cell_4929 ( .C (CLK), .D (signal_7072), .Q (signal_7073) ) ;
    buf_clk cell_4945 ( .C (CLK), .D (signal_7088), .Q (signal_7089) ) ;
    buf_clk cell_4961 ( .C (CLK), .D (signal_7104), .Q (signal_7105) ) ;
    buf_clk cell_4977 ( .C (CLK), .D (signal_7120), .Q (signal_7121) ) ;
    buf_clk cell_4993 ( .C (CLK), .D (signal_7136), .Q (signal_7137) ) ;
    buf_clk cell_5009 ( .C (CLK), .D (signal_7152), .Q (signal_7153) ) ;
    buf_clk cell_5025 ( .C (CLK), .D (signal_7168), .Q (signal_7169) ) ;
    buf_clk cell_5041 ( .C (CLK), .D (signal_7184), .Q (signal_7185) ) ;
    buf_clk cell_5057 ( .C (CLK), .D (signal_7200), .Q (signal_7201) ) ;
    buf_clk cell_5073 ( .C (CLK), .D (signal_7216), .Q (signal_7217) ) ;
    buf_clk cell_5089 ( .C (CLK), .D (signal_7232), .Q (signal_7233) ) ;
    buf_clk cell_5105 ( .C (CLK), .D (signal_7248), .Q (signal_7249) ) ;
    buf_clk cell_5121 ( .C (CLK), .D (signal_7264), .Q (signal_7265) ) ;
    buf_clk cell_5137 ( .C (CLK), .D (signal_7280), .Q (signal_7281) ) ;
    buf_clk cell_5153 ( .C (CLK), .D (signal_7296), .Q (signal_7297) ) ;
    buf_clk cell_5169 ( .C (CLK), .D (signal_7312), .Q (signal_7313) ) ;
    buf_clk cell_5185 ( .C (CLK), .D (signal_7328), .Q (signal_7329) ) ;
    buf_clk cell_5201 ( .C (CLK), .D (signal_7344), .Q (signal_7345) ) ;
    buf_clk cell_5217 ( .C (CLK), .D (signal_7360), .Q (signal_7361) ) ;
    buf_clk cell_5233 ( .C (CLK), .D (signal_7376), .Q (signal_7377) ) ;
    buf_clk cell_5249 ( .C (CLK), .D (signal_7392), .Q (signal_7393) ) ;
    buf_clk cell_5265 ( .C (CLK), .D (signal_7408), .Q (signal_7409) ) ;
    buf_clk cell_5281 ( .C (CLK), .D (signal_7424), .Q (signal_7425) ) ;
    buf_clk cell_5297 ( .C (CLK), .D (signal_7440), .Q (signal_7441) ) ;
    buf_clk cell_5313 ( .C (CLK), .D (signal_7456), .Q (signal_7457) ) ;
    buf_clk cell_5329 ( .C (CLK), .D (signal_7472), .Q (signal_7473) ) ;
    buf_clk cell_5345 ( .C (CLK), .D (signal_7488), .Q (signal_7489) ) ;
    buf_clk cell_5361 ( .C (CLK), .D (signal_7504), .Q (signal_7505) ) ;
    buf_clk cell_5377 ( .C (CLK), .D (signal_7520), .Q (signal_7521) ) ;
    buf_clk cell_5393 ( .C (CLK), .D (signal_7536), .Q (signal_7537) ) ;
    buf_clk cell_5409 ( .C (CLK), .D (signal_7552), .Q (signal_7553) ) ;
    buf_clk cell_5425 ( .C (CLK), .D (signal_7568), .Q (signal_7569) ) ;
    buf_clk cell_5441 ( .C (CLK), .D (signal_7584), .Q (signal_7585) ) ;
    buf_clk cell_5457 ( .C (CLK), .D (signal_7600), .Q (signal_7601) ) ;
    buf_clk cell_5473 ( .C (CLK), .D (signal_7616), .Q (signal_7617) ) ;
    buf_clk cell_5489 ( .C (CLK), .D (signal_7632), .Q (signal_7633) ) ;
    buf_clk cell_5505 ( .C (CLK), .D (signal_7648), .Q (signal_7649) ) ;
    buf_clk cell_5521 ( .C (CLK), .D (signal_7664), .Q (signal_7665) ) ;
    buf_clk cell_5537 ( .C (CLK), .D (signal_7680), .Q (signal_7681) ) ;
    buf_clk cell_5553 ( .C (CLK), .D (signal_7696), .Q (signal_7697) ) ;
    buf_clk cell_5569 ( .C (CLK), .D (signal_7712), .Q (signal_7713) ) ;
    buf_clk cell_5585 ( .C (CLK), .D (signal_7728), .Q (signal_7729) ) ;
    buf_clk cell_5601 ( .C (CLK), .D (signal_7744), .Q (signal_7745) ) ;
    buf_clk cell_5617 ( .C (CLK), .D (signal_7760), .Q (signal_7761) ) ;
    buf_clk cell_5633 ( .C (CLK), .D (signal_7776), .Q (signal_7777) ) ;
    buf_clk cell_5649 ( .C (CLK), .D (signal_7792), .Q (signal_7793) ) ;
    buf_clk cell_5665 ( .C (CLK), .D (signal_7808), .Q (signal_7809) ) ;
    buf_clk cell_5681 ( .C (CLK), .D (signal_7824), .Q (signal_7825) ) ;
    buf_clk cell_5697 ( .C (CLK), .D (signal_7840), .Q (signal_7841) ) ;
    buf_clk cell_5713 ( .C (CLK), .D (signal_7856), .Q (signal_7857) ) ;
    buf_clk cell_5729 ( .C (CLK), .D (signal_7872), .Q (signal_7873) ) ;
    buf_clk cell_5745 ( .C (CLK), .D (signal_7888), .Q (signal_7889) ) ;
    buf_clk cell_5761 ( .C (CLK), .D (signal_7904), .Q (signal_7905) ) ;
    buf_clk cell_5777 ( .C (CLK), .D (signal_7920), .Q (signal_7921) ) ;
    buf_clk cell_5793 ( .C (CLK), .D (signal_7936), .Q (signal_7937) ) ;
    buf_clk cell_5809 ( .C (CLK), .D (signal_7952), .Q (signal_7953) ) ;
    buf_clk cell_5825 ( .C (CLK), .D (signal_7968), .Q (signal_7969) ) ;
    buf_clk cell_5841 ( .C (CLK), .D (signal_7984), .Q (signal_7985) ) ;
    buf_clk cell_5857 ( .C (CLK), .D (signal_8000), .Q (signal_8001) ) ;
    buf_clk cell_5873 ( .C (CLK), .D (signal_8016), .Q (signal_8017) ) ;
    buf_clk cell_5889 ( .C (CLK), .D (signal_8032), .Q (signal_8033) ) ;
    buf_clk cell_5905 ( .C (CLK), .D (signal_8048), .Q (signal_8049) ) ;
    buf_clk cell_5921 ( .C (CLK), .D (signal_8064), .Q (signal_8065) ) ;
    buf_clk cell_5937 ( .C (CLK), .D (signal_8080), .Q (signal_8081) ) ;
    buf_clk cell_5953 ( .C (CLK), .D (signal_8096), .Q (signal_8097) ) ;
    buf_clk cell_5969 ( .C (CLK), .D (signal_8112), .Q (signal_8113) ) ;
    buf_clk cell_5985 ( .C (CLK), .D (signal_8128), .Q (signal_8129) ) ;
    buf_clk cell_6001 ( .C (CLK), .D (signal_8144), .Q (signal_8145) ) ;
    buf_clk cell_6017 ( .C (CLK), .D (signal_8160), .Q (signal_8161) ) ;
    buf_clk cell_6033 ( .C (CLK), .D (signal_8176), .Q (signal_8177) ) ;
    buf_clk cell_6049 ( .C (CLK), .D (signal_8192), .Q (signal_8193) ) ;
    buf_clk cell_6065 ( .C (CLK), .D (signal_8208), .Q (signal_8209) ) ;
    buf_clk cell_6081 ( .C (CLK), .D (signal_8224), .Q (signal_8225) ) ;
    buf_clk cell_6097 ( .C (CLK), .D (signal_8240), .Q (signal_8241) ) ;
    buf_clk cell_6113 ( .C (CLK), .D (signal_8256), .Q (signal_8257) ) ;
    buf_clk cell_6129 ( .C (CLK), .D (signal_8272), .Q (signal_8273) ) ;
    buf_clk cell_6145 ( .C (CLK), .D (signal_8288), .Q (signal_8289) ) ;
    buf_clk cell_6161 ( .C (CLK), .D (signal_8304), .Q (signal_8305) ) ;
    buf_clk cell_6177 ( .C (CLK), .D (signal_8320), .Q (signal_8321) ) ;
    buf_clk cell_6193 ( .C (CLK), .D (signal_8336), .Q (signal_8337) ) ;
    buf_clk cell_6209 ( .C (CLK), .D (signal_8352), .Q (signal_8353) ) ;
    buf_clk cell_6225 ( .C (CLK), .D (signal_8368), .Q (signal_8369) ) ;
    buf_clk cell_6241 ( .C (CLK), .D (signal_8384), .Q (signal_8385) ) ;
    buf_clk cell_6257 ( .C (CLK), .D (signal_8400), .Q (signal_8401) ) ;
    buf_clk cell_6273 ( .C (CLK), .D (signal_8416), .Q (signal_8417) ) ;
    buf_clk cell_6289 ( .C (CLK), .D (signal_8432), .Q (signal_8433) ) ;
    buf_clk cell_6305 ( .C (CLK), .D (signal_8448), .Q (signal_8449) ) ;
    buf_clk cell_6321 ( .C (CLK), .D (signal_8464), .Q (signal_8465) ) ;
    buf_clk cell_6337 ( .C (CLK), .D (signal_8480), .Q (signal_8481) ) ;
    buf_clk cell_6353 ( .C (CLK), .D (signal_8496), .Q (signal_8497) ) ;
    buf_clk cell_6369 ( .C (CLK), .D (signal_8512), .Q (signal_8513) ) ;
    buf_clk cell_6385 ( .C (CLK), .D (signal_8528), .Q (signal_8529) ) ;
    buf_clk cell_6401 ( .C (CLK), .D (signal_8544), .Q (signal_8545) ) ;
    buf_clk cell_6409 ( .C (CLK), .D (signal_8552), .Q (signal_8553) ) ;
    buf_clk cell_6417 ( .C (CLK), .D (signal_8560), .Q (signal_8561) ) ;
    buf_clk cell_6425 ( .C (CLK), .D (signal_8568), .Q (signal_8569) ) ;
    buf_clk cell_6433 ( .C (CLK), .D (signal_8576), .Q (signal_8577) ) ;
    buf_clk cell_6441 ( .C (CLK), .D (signal_8584), .Q (signal_8585) ) ;
    buf_clk cell_6449 ( .C (CLK), .D (signal_8592), .Q (signal_8593) ) ;
    buf_clk cell_6457 ( .C (CLK), .D (signal_8600), .Q (signal_8601) ) ;
    buf_clk cell_6465 ( .C (CLK), .D (signal_8608), .Q (signal_8609) ) ;
    buf_clk cell_6473 ( .C (CLK), .D (signal_8616), .Q (signal_8617) ) ;
    buf_clk cell_6481 ( .C (CLK), .D (signal_8624), .Q (signal_8625) ) ;
    buf_clk cell_6489 ( .C (CLK), .D (signal_8632), .Q (signal_8633) ) ;
    buf_clk cell_6497 ( .C (CLK), .D (signal_8640), .Q (signal_8641) ) ;
    buf_clk cell_6505 ( .C (CLK), .D (signal_8648), .Q (signal_8649) ) ;
    buf_clk cell_6513 ( .C (CLK), .D (signal_8656), .Q (signal_8657) ) ;
    buf_clk cell_6521 ( .C (CLK), .D (signal_8664), .Q (signal_8665) ) ;
    buf_clk cell_6529 ( .C (CLK), .D (signal_8672), .Q (signal_8673) ) ;
    buf_clk cell_6537 ( .C (CLK), .D (signal_8680), .Q (signal_8681) ) ;
    buf_clk cell_6545 ( .C (CLK), .D (signal_8688), .Q (signal_8689) ) ;
    buf_clk cell_6553 ( .C (CLK), .D (signal_8696), .Q (signal_8697) ) ;
    buf_clk cell_6561 ( .C (CLK), .D (signal_8704), .Q (signal_8705) ) ;
    buf_clk cell_6569 ( .C (CLK), .D (signal_8712), .Q (signal_8713) ) ;
    buf_clk cell_6577 ( .C (CLK), .D (signal_8720), .Q (signal_8721) ) ;
    buf_clk cell_6585 ( .C (CLK), .D (signal_8728), .Q (signal_8729) ) ;
    buf_clk cell_6593 ( .C (CLK), .D (signal_8736), .Q (signal_8737) ) ;
    buf_clk cell_6601 ( .C (CLK), .D (signal_8744), .Q (signal_8745) ) ;
    buf_clk cell_6609 ( .C (CLK), .D (signal_8752), .Q (signal_8753) ) ;
    buf_clk cell_6617 ( .C (CLK), .D (signal_8760), .Q (signal_8761) ) ;
    buf_clk cell_6625 ( .C (CLK), .D (signal_8768), .Q (signal_8769) ) ;
    buf_clk cell_6633 ( .C (CLK), .D (signal_8776), .Q (signal_8777) ) ;
    buf_clk cell_6641 ( .C (CLK), .D (signal_8784), .Q (signal_8785) ) ;
    buf_clk cell_6649 ( .C (CLK), .D (signal_8792), .Q (signal_8793) ) ;
    buf_clk cell_6657 ( .C (CLK), .D (signal_8800), .Q (signal_8801) ) ;
    buf_clk cell_6665 ( .C (CLK), .D (signal_8808), .Q (signal_8809) ) ;
    buf_clk cell_6673 ( .C (CLK), .D (signal_8816), .Q (signal_8817) ) ;
    buf_clk cell_6681 ( .C (CLK), .D (signal_8824), .Q (signal_8825) ) ;
    buf_clk cell_6689 ( .C (CLK), .D (signal_8832), .Q (signal_8833) ) ;
    buf_clk cell_6697 ( .C (CLK), .D (signal_8840), .Q (signal_8841) ) ;
    buf_clk cell_6705 ( .C (CLK), .D (signal_8848), .Q (signal_8849) ) ;
    buf_clk cell_6713 ( .C (CLK), .D (signal_8856), .Q (signal_8857) ) ;
    buf_clk cell_6721 ( .C (CLK), .D (signal_8864), .Q (signal_8865) ) ;
    buf_clk cell_6729 ( .C (CLK), .D (signal_8872), .Q (signal_8873) ) ;
    buf_clk cell_6737 ( .C (CLK), .D (signal_8880), .Q (signal_8881) ) ;
    buf_clk cell_6745 ( .C (CLK), .D (signal_8888), .Q (signal_8889) ) ;
    buf_clk cell_6753 ( .C (CLK), .D (signal_8896), .Q (signal_8897) ) ;
    buf_clk cell_6761 ( .C (CLK), .D (signal_8904), .Q (signal_8905) ) ;
    buf_clk cell_6769 ( .C (CLK), .D (signal_8912), .Q (signal_8913) ) ;
    buf_clk cell_6777 ( .C (CLK), .D (signal_8920), .Q (signal_8921) ) ;
    buf_clk cell_6785 ( .C (CLK), .D (signal_8928), .Q (signal_8929) ) ;
    buf_clk cell_6793 ( .C (CLK), .D (signal_8936), .Q (signal_8937) ) ;
    buf_clk cell_6801 ( .C (CLK), .D (signal_8944), .Q (signal_8945) ) ;
    buf_clk cell_6809 ( .C (CLK), .D (signal_8952), .Q (signal_8953) ) ;
    buf_clk cell_6817 ( .C (CLK), .D (signal_8960), .Q (signal_8961) ) ;
    buf_clk cell_6825 ( .C (CLK), .D (signal_8968), .Q (signal_8969) ) ;
    buf_clk cell_6833 ( .C (CLK), .D (signal_8976), .Q (signal_8977) ) ;
    buf_clk cell_6841 ( .C (CLK), .D (signal_8984), .Q (signal_8985) ) ;
    buf_clk cell_6849 ( .C (CLK), .D (signal_8992), .Q (signal_8993) ) ;
    buf_clk cell_6857 ( .C (CLK), .D (signal_9000), .Q (signal_9001) ) ;
    buf_clk cell_6865 ( .C (CLK), .D (signal_9008), .Q (signal_9009) ) ;
    buf_clk cell_6873 ( .C (CLK), .D (signal_9016), .Q (signal_9017) ) ;
    buf_clk cell_6881 ( .C (CLK), .D (signal_9024), .Q (signal_9025) ) ;
    buf_clk cell_6889 ( .C (CLK), .D (signal_9032), .Q (signal_9033) ) ;
    buf_clk cell_6897 ( .C (CLK), .D (signal_9040), .Q (signal_9041) ) ;
    buf_clk cell_6905 ( .C (CLK), .D (signal_9048), .Q (signal_9049) ) ;
    buf_clk cell_6913 ( .C (CLK), .D (signal_9056), .Q (signal_9057) ) ;
    buf_clk cell_6921 ( .C (CLK), .D (signal_9064), .Q (signal_9065) ) ;
    buf_clk cell_6929 ( .C (CLK), .D (signal_9072), .Q (signal_9073) ) ;
    buf_clk cell_6937 ( .C (CLK), .D (signal_9080), .Q (signal_9081) ) ;
    buf_clk cell_6945 ( .C (CLK), .D (signal_9088), .Q (signal_9089) ) ;
    buf_clk cell_6953 ( .C (CLK), .D (signal_9096), .Q (signal_9097) ) ;
    buf_clk cell_6961 ( .C (CLK), .D (signal_9104), .Q (signal_9105) ) ;
    buf_clk cell_6969 ( .C (CLK), .D (signal_9112), .Q (signal_9113) ) ;
    buf_clk cell_6977 ( .C (CLK), .D (signal_9120), .Q (signal_9121) ) ;
    buf_clk cell_6985 ( .C (CLK), .D (signal_9128), .Q (signal_9129) ) ;
    buf_clk cell_6993 ( .C (CLK), .D (signal_9136), .Q (signal_9137) ) ;
    buf_clk cell_7001 ( .C (CLK), .D (signal_9144), .Q (signal_9145) ) ;
    buf_clk cell_7009 ( .C (CLK), .D (signal_9152), .Q (signal_9153) ) ;
    buf_clk cell_7017 ( .C (CLK), .D (signal_9160), .Q (signal_9161) ) ;
    buf_clk cell_7025 ( .C (CLK), .D (signal_9168), .Q (signal_9169) ) ;
    buf_clk cell_7033 ( .C (CLK), .D (signal_9176), .Q (signal_9177) ) ;
    buf_clk cell_7041 ( .C (CLK), .D (signal_9184), .Q (signal_9185) ) ;
    buf_clk cell_7049 ( .C (CLK), .D (signal_9192), .Q (signal_9193) ) ;
    buf_clk cell_7057 ( .C (CLK), .D (signal_9200), .Q (signal_9201) ) ;
    buf_clk cell_7065 ( .C (CLK), .D (signal_9208), .Q (signal_9209) ) ;
    buf_clk cell_7073 ( .C (CLK), .D (signal_9216), .Q (signal_9217) ) ;
    buf_clk cell_7081 ( .C (CLK), .D (signal_9224), .Q (signal_9225) ) ;
    buf_clk cell_7089 ( .C (CLK), .D (signal_9232), .Q (signal_9233) ) ;
    buf_clk cell_7097 ( .C (CLK), .D (signal_9240), .Q (signal_9241) ) ;
    buf_clk cell_7105 ( .C (CLK), .D (signal_9248), .Q (signal_9249) ) ;
    buf_clk cell_7113 ( .C (CLK), .D (signal_9256), .Q (signal_9257) ) ;
    buf_clk cell_7121 ( .C (CLK), .D (signal_9264), .Q (signal_9265) ) ;
    buf_clk cell_7129 ( .C (CLK), .D (signal_9272), .Q (signal_9273) ) ;
    buf_clk cell_7137 ( .C (CLK), .D (signal_9280), .Q (signal_9281) ) ;
    buf_clk cell_7145 ( .C (CLK), .D (signal_9288), .Q (signal_9289) ) ;
    buf_clk cell_7153 ( .C (CLK), .D (signal_9296), .Q (signal_9297) ) ;
    buf_clk cell_7161 ( .C (CLK), .D (signal_9304), .Q (signal_9305) ) ;
    buf_clk cell_7169 ( .C (CLK), .D (signal_9312), .Q (signal_9313) ) ;
    buf_clk cell_7177 ( .C (CLK), .D (signal_9320), .Q (signal_9321) ) ;
    buf_clk cell_7185 ( .C (CLK), .D (signal_9328), .Q (signal_9329) ) ;
    buf_clk cell_7193 ( .C (CLK), .D (signal_9336), .Q (signal_9337) ) ;
    buf_clk cell_7201 ( .C (CLK), .D (signal_9344), .Q (signal_9345) ) ;
    buf_clk cell_7209 ( .C (CLK), .D (signal_9352), .Q (signal_9353) ) ;
    buf_clk cell_7217 ( .C (CLK), .D (signal_9360), .Q (signal_9361) ) ;
    buf_clk cell_7225 ( .C (CLK), .D (signal_9368), .Q (signal_9369) ) ;
    buf_clk cell_7233 ( .C (CLK), .D (signal_9376), .Q (signal_9377) ) ;
    buf_clk cell_7241 ( .C (CLK), .D (signal_9384), .Q (signal_9385) ) ;
    buf_clk cell_7249 ( .C (CLK), .D (signal_9392), .Q (signal_9393) ) ;
    buf_clk cell_7257 ( .C (CLK), .D (signal_9400), .Q (signal_9401) ) ;
    buf_clk cell_7265 ( .C (CLK), .D (signal_9408), .Q (signal_9409) ) ;
    buf_clk cell_7273 ( .C (CLK), .D (signal_9416), .Q (signal_9417) ) ;
    buf_clk cell_7281 ( .C (CLK), .D (signal_9424), .Q (signal_9425) ) ;
    buf_clk cell_7289 ( .C (CLK), .D (signal_9432), .Q (signal_9433) ) ;
    buf_clk cell_7297 ( .C (CLK), .D (signal_9440), .Q (signal_9441) ) ;
    buf_clk cell_7305 ( .C (CLK), .D (signal_9448), .Q (signal_9449) ) ;
    buf_clk cell_7313 ( .C (CLK), .D (signal_9456), .Q (signal_9457) ) ;
    buf_clk cell_7321 ( .C (CLK), .D (signal_9464), .Q (signal_9465) ) ;
    buf_clk cell_7329 ( .C (CLK), .D (signal_9472), .Q (signal_9473) ) ;
    buf_clk cell_7337 ( .C (CLK), .D (signal_9480), .Q (signal_9481) ) ;
    buf_clk cell_7345 ( .C (CLK), .D (signal_9488), .Q (signal_9489) ) ;
    buf_clk cell_7353 ( .C (CLK), .D (signal_9496), .Q (signal_9497) ) ;
    buf_clk cell_7361 ( .C (CLK), .D (signal_9504), .Q (signal_9505) ) ;
    buf_clk cell_7369 ( .C (CLK), .D (signal_9512), .Q (signal_9513) ) ;
    buf_clk cell_7377 ( .C (CLK), .D (signal_9520), .Q (signal_9521) ) ;
    buf_clk cell_7385 ( .C (CLK), .D (signal_9528), .Q (signal_9529) ) ;
    buf_clk cell_7393 ( .C (CLK), .D (signal_9536), .Q (signal_9537) ) ;
    buf_clk cell_7401 ( .C (CLK), .D (signal_9544), .Q (signal_9545) ) ;
    buf_clk cell_7409 ( .C (CLK), .D (signal_9552), .Q (signal_9553) ) ;
    buf_clk cell_7417 ( .C (CLK), .D (signal_9560), .Q (signal_9561) ) ;
    buf_clk cell_7425 ( .C (CLK), .D (signal_9568), .Q (signal_9569) ) ;
    buf_clk cell_7433 ( .C (CLK), .D (signal_9576), .Q (signal_9577) ) ;
    buf_clk cell_7441 ( .C (CLK), .D (signal_9584), .Q (signal_9585) ) ;
    buf_clk cell_7449 ( .C (CLK), .D (signal_9592), .Q (signal_9593) ) ;
    buf_clk cell_7457 ( .C (CLK), .D (signal_9600), .Q (signal_9601) ) ;
    buf_clk cell_7465 ( .C (CLK), .D (signal_9608), .Q (signal_9609) ) ;
    buf_clk cell_7473 ( .C (CLK), .D (signal_9616), .Q (signal_9617) ) ;
    buf_clk cell_7481 ( .C (CLK), .D (signal_9624), .Q (signal_9625) ) ;
    buf_clk cell_7489 ( .C (CLK), .D (signal_9632), .Q (signal_9633) ) ;
    buf_clk cell_7497 ( .C (CLK), .D (signal_9640), .Q (signal_9641) ) ;
    buf_clk cell_7505 ( .C (CLK), .D (signal_9648), .Q (signal_9649) ) ;
    buf_clk cell_7513 ( .C (CLK), .D (signal_9656), .Q (signal_9657) ) ;
    buf_clk cell_7521 ( .C (CLK), .D (signal_9664), .Q (signal_9665) ) ;
    buf_clk cell_7529 ( .C (CLK), .D (signal_9672), .Q (signal_9673) ) ;
    buf_clk cell_7537 ( .C (CLK), .D (signal_9680), .Q (signal_9681) ) ;
    buf_clk cell_7545 ( .C (CLK), .D (signal_9688), .Q (signal_9689) ) ;
    buf_clk cell_7553 ( .C (CLK), .D (signal_9696), .Q (signal_9697) ) ;
    buf_clk cell_7567 ( .C (CLK), .D (signal_9710), .Q (signal_9711) ) ;
    buf_clk cell_7575 ( .C (CLK), .D (signal_9718), .Q (signal_9719) ) ;
    buf_clk cell_7579 ( .C (CLK), .D (signal_9722), .Q (signal_9723) ) ;
    buf_clk cell_7583 ( .C (CLK), .D (signal_9726), .Q (signal_9727) ) ;
    buf_clk cell_7601 ( .C (CLK), .D (signal_9744), .Q (signal_9745) ) ;
    buf_clk cell_7617 ( .C (CLK), .D (signal_9760), .Q (signal_9761) ) ;
    buf_clk cell_7633 ( .C (CLK), .D (signal_9776), .Q (signal_9777) ) ;
    buf_clk cell_7649 ( .C (CLK), .D (signal_9792), .Q (signal_9793) ) ;
    buf_clk cell_7665 ( .C (CLK), .D (signal_9808), .Q (signal_9809) ) ;
    buf_clk cell_7681 ( .C (CLK), .D (signal_9824), .Q (signal_9825) ) ;
    buf_clk cell_7697 ( .C (CLK), .D (signal_9840), .Q (signal_9841) ) ;
    buf_clk cell_7713 ( .C (CLK), .D (signal_9856), .Q (signal_9857) ) ;
    buf_clk cell_7729 ( .C (CLK), .D (signal_9872), .Q (signal_9873) ) ;
    buf_clk cell_7745 ( .C (CLK), .D (signal_9888), .Q (signal_9889) ) ;
    buf_clk cell_7753 ( .C (CLK), .D (signal_9896), .Q (signal_9897) ) ;
    buf_clk cell_7761 ( .C (CLK), .D (signal_9904), .Q (signal_9905) ) ;
    buf_clk cell_7769 ( .C (CLK), .D (signal_9912), .Q (signal_9913) ) ;
    buf_clk cell_7777 ( .C (CLK), .D (signal_9920), .Q (signal_9921) ) ;
    buf_clk cell_7785 ( .C (CLK), .D (signal_9928), .Q (signal_9929) ) ;
    buf_clk cell_7793 ( .C (CLK), .D (signal_9936), .Q (signal_9937) ) ;
    buf_clk cell_7801 ( .C (CLK), .D (signal_9944), .Q (signal_9945) ) ;
    buf_clk cell_7809 ( .C (CLK), .D (signal_9952), .Q (signal_9953) ) ;
    buf_clk cell_7817 ( .C (CLK), .D (signal_9960), .Q (signal_9961) ) ;
    buf_clk cell_7825 ( .C (CLK), .D (signal_9968), .Q (signal_9969) ) ;
    buf_clk cell_7833 ( .C (CLK), .D (signal_9976), .Q (signal_9977) ) ;
    buf_clk cell_7841 ( .C (CLK), .D (signal_9984), .Q (signal_9985) ) ;
    buf_clk cell_7849 ( .C (CLK), .D (signal_9992), .Q (signal_9993) ) ;
    buf_clk cell_7857 ( .C (CLK), .D (signal_10000), .Q (signal_10001) ) ;
    buf_clk cell_7865 ( .C (CLK), .D (signal_10008), .Q (signal_10009) ) ;
    buf_clk cell_7873 ( .C (CLK), .D (signal_10016), .Q (signal_10017) ) ;
    buf_clk cell_7881 ( .C (CLK), .D (signal_10024), .Q (signal_10025) ) ;
    buf_clk cell_7889 ( .C (CLK), .D (signal_10032), .Q (signal_10033) ) ;
    buf_clk cell_7897 ( .C (CLK), .D (signal_10040), .Q (signal_10041) ) ;
    buf_clk cell_7905 ( .C (CLK), .D (signal_10048), .Q (signal_10049) ) ;
    buf_clk cell_7913 ( .C (CLK), .D (signal_10056), .Q (signal_10057) ) ;
    buf_clk cell_7921 ( .C (CLK), .D (signal_10064), .Q (signal_10065) ) ;
    buf_clk cell_7929 ( .C (CLK), .D (signal_10072), .Q (signal_10073) ) ;
    buf_clk cell_7937 ( .C (CLK), .D (signal_10080), .Q (signal_10081) ) ;
    buf_clk cell_7953 ( .C (CLK), .D (signal_10096), .Q (signal_10097) ) ;

    /* cells in depth 13 */
    buf_clk cell_3442 ( .C (CLK), .D (signal_5585), .Q (signal_5586) ) ;
    buf_clk cell_3458 ( .C (CLK), .D (signal_5601), .Q (signal_5602) ) ;
    buf_clk cell_3474 ( .C (CLK), .D (signal_5617), .Q (signal_5618) ) ;
    buf_clk cell_3482 ( .C (CLK), .D (signal_5625), .Q (signal_5626) ) ;
    buf_clk cell_3498 ( .C (CLK), .D (signal_5641), .Q (signal_5642) ) ;
    buf_clk cell_3514 ( .C (CLK), .D (signal_5657), .Q (signal_5658) ) ;
    buf_clk cell_3522 ( .C (CLK), .D (signal_5665), .Q (signal_5666) ) ;
    buf_clk cell_3538 ( .C (CLK), .D (signal_5681), .Q (signal_5682) ) ;
    buf_clk cell_3554 ( .C (CLK), .D (signal_5697), .Q (signal_5698) ) ;
    buf_clk cell_3570 ( .C (CLK), .D (signal_5713), .Q (signal_5714) ) ;
    buf_clk cell_3586 ( .C (CLK), .D (signal_5729), .Q (signal_5730) ) ;
    buf_clk cell_3590 ( .C (CLK), .D (signal_5545), .Q (signal_5734) ) ;
    buf_clk cell_3594 ( .C (CLK), .D (signal_5549), .Q (signal_5738) ) ;
    buf_clk cell_3600 ( .C (CLK), .D (signal_5743), .Q (signal_5744) ) ;
    buf_clk cell_3606 ( .C (CLK), .D (signal_5749), .Q (signal_5750) ) ;
    buf_clk cell_3612 ( .C (CLK), .D (signal_5755), .Q (signal_5756) ) ;
    buf_clk cell_3618 ( .C (CLK), .D (signal_5761), .Q (signal_5762) ) ;
    buf_clk cell_3624 ( .C (CLK), .D (signal_5767), .Q (signal_5768) ) ;
    buf_clk cell_3630 ( .C (CLK), .D (signal_5773), .Q (signal_5774) ) ;
    buf_clk cell_3646 ( .C (CLK), .D (signal_5789), .Q (signal_5790) ) ;
    buf_clk cell_3662 ( .C (CLK), .D (signal_5805), .Q (signal_5806) ) ;
    buf_clk cell_3678 ( .C (CLK), .D (signal_5821), .Q (signal_5822) ) ;
    buf_clk cell_3694 ( .C (CLK), .D (signal_5837), .Q (signal_5838) ) ;
    buf_clk cell_3710 ( .C (CLK), .D (signal_5853), .Q (signal_5854) ) ;
    buf_clk cell_3726 ( .C (CLK), .D (signal_5869), .Q (signal_5870) ) ;
    buf_clk cell_3742 ( .C (CLK), .D (signal_5885), .Q (signal_5886) ) ;
    buf_clk cell_3758 ( .C (CLK), .D (signal_5901), .Q (signal_5902) ) ;
    buf_clk cell_3774 ( .C (CLK), .D (signal_5917), .Q (signal_5918) ) ;
    buf_clk cell_3790 ( .C (CLK), .D (signal_5933), .Q (signal_5934) ) ;
    buf_clk cell_3794 ( .C (CLK), .D (signal_5433), .Q (signal_5938) ) ;
    buf_clk cell_3798 ( .C (CLK), .D (signal_5437), .Q (signal_5942) ) ;
    buf_clk cell_3806 ( .C (CLK), .D (signal_5949), .Q (signal_5950) ) ;
    buf_clk cell_3814 ( .C (CLK), .D (signal_5957), .Q (signal_5958) ) ;
    buf_clk cell_3820 ( .C (CLK), .D (signal_5963), .Q (signal_5964) ) ;
    buf_clk cell_3826 ( .C (CLK), .D (signal_5969), .Q (signal_5970) ) ;
    buf_clk cell_3834 ( .C (CLK), .D (signal_5977), .Q (signal_5978) ) ;
    buf_clk cell_3842 ( .C (CLK), .D (signal_5985), .Q (signal_5986) ) ;
    buf_clk cell_3850 ( .C (CLK), .D (signal_5993), .Q (signal_5994) ) ;
    buf_clk cell_3858 ( .C (CLK), .D (signal_6001), .Q (signal_6002) ) ;
    buf_clk cell_3862 ( .C (CLK), .D (signal_5469), .Q (signal_6006) ) ;
    buf_clk cell_3866 ( .C (CLK), .D (signal_5477), .Q (signal_6010) ) ;
    buf_clk cell_3874 ( .C (CLK), .D (signal_6017), .Q (signal_6018) ) ;
    buf_clk cell_3882 ( .C (CLK), .D (signal_6025), .Q (signal_6026) ) ;
    buf_clk cell_3898 ( .C (CLK), .D (signal_6041), .Q (signal_6042) ) ;
    buf_clk cell_3914 ( .C (CLK), .D (signal_6057), .Q (signal_6058) ) ;
    buf_clk cell_3930 ( .C (CLK), .D (signal_6073), .Q (signal_6074) ) ;
    buf_clk cell_3946 ( .C (CLK), .D (signal_6089), .Q (signal_6090) ) ;
    buf_clk cell_3962 ( .C (CLK), .D (signal_6105), .Q (signal_6106) ) ;
    buf_clk cell_3978 ( .C (CLK), .D (signal_6121), .Q (signal_6122) ) ;
    buf_clk cell_3994 ( .C (CLK), .D (signal_6137), .Q (signal_6138) ) ;
    buf_clk cell_4010 ( .C (CLK), .D (signal_6153), .Q (signal_6154) ) ;
    buf_clk cell_4026 ( .C (CLK), .D (signal_6169), .Q (signal_6170) ) ;
    buf_clk cell_4042 ( .C (CLK), .D (signal_6185), .Q (signal_6186) ) ;
    buf_clk cell_4058 ( .C (CLK), .D (signal_6201), .Q (signal_6202) ) ;
    buf_clk cell_4074 ( .C (CLK), .D (signal_6217), .Q (signal_6218) ) ;
    buf_clk cell_4090 ( .C (CLK), .D (signal_6233), .Q (signal_6234) ) ;
    buf_clk cell_4106 ( .C (CLK), .D (signal_6249), .Q (signal_6250) ) ;
    buf_clk cell_4116 ( .C (CLK), .D (signal_6259), .Q (signal_6260) ) ;
    buf_clk cell_4126 ( .C (CLK), .D (signal_6269), .Q (signal_6270) ) ;
    buf_clk cell_4132 ( .C (CLK), .D (signal_6275), .Q (signal_6276) ) ;
    buf_clk cell_4138 ( .C (CLK), .D (signal_6281), .Q (signal_6282) ) ;
    buf_clk cell_4146 ( .C (CLK), .D (signal_6289), .Q (signal_6290) ) ;
    buf_clk cell_4154 ( .C (CLK), .D (signal_6297), .Q (signal_6298) ) ;
    buf_clk cell_4164 ( .C (CLK), .D (signal_6307), .Q (signal_6308) ) ;
    buf_clk cell_4174 ( .C (CLK), .D (signal_6317), .Q (signal_6318) ) ;
    buf_clk cell_4190 ( .C (CLK), .D (signal_6333), .Q (signal_6334) ) ;
    buf_clk cell_4202 ( .C (CLK), .D (signal_6345), .Q (signal_6346) ) ;
    buf_clk cell_4214 ( .C (CLK), .D (signal_6357), .Q (signal_6358) ) ;
    buf_clk cell_4222 ( .C (CLK), .D (signal_6365), .Q (signal_6366) ) ;
    buf_clk cell_4230 ( .C (CLK), .D (signal_6373), .Q (signal_6374) ) ;
    buf_clk cell_4242 ( .C (CLK), .D (signal_6385), .Q (signal_6386) ) ;
    buf_clk cell_4254 ( .C (CLK), .D (signal_6397), .Q (signal_6398) ) ;
    buf_clk cell_4268 ( .C (CLK), .D (signal_6411), .Q (signal_6412) ) ;
    buf_clk cell_4282 ( .C (CLK), .D (signal_6425), .Q (signal_6426) ) ;
    buf_clk cell_4298 ( .C (CLK), .D (signal_6441), .Q (signal_6442) ) ;
    buf_clk cell_4314 ( .C (CLK), .D (signal_6457), .Q (signal_6458) ) ;
    buf_clk cell_4330 ( .C (CLK), .D (signal_6473), .Q (signal_6474) ) ;
    buf_clk cell_4346 ( .C (CLK), .D (signal_6489), .Q (signal_6490) ) ;
    buf_clk cell_4362 ( .C (CLK), .D (signal_6505), .Q (signal_6506) ) ;
    buf_clk cell_4378 ( .C (CLK), .D (signal_6521), .Q (signal_6522) ) ;
    buf_clk cell_4394 ( .C (CLK), .D (signal_6537), .Q (signal_6538) ) ;
    buf_clk cell_4410 ( .C (CLK), .D (signal_6553), .Q (signal_6554) ) ;
    buf_clk cell_4426 ( .C (CLK), .D (signal_6569), .Q (signal_6570) ) ;
    buf_clk cell_4442 ( .C (CLK), .D (signal_6585), .Q (signal_6586) ) ;
    buf_clk cell_4458 ( .C (CLK), .D (signal_6601), .Q (signal_6602) ) ;
    buf_clk cell_4474 ( .C (CLK), .D (signal_6617), .Q (signal_6618) ) ;
    buf_clk cell_4490 ( .C (CLK), .D (signal_6633), .Q (signal_6634) ) ;
    buf_clk cell_4506 ( .C (CLK), .D (signal_6649), .Q (signal_6650) ) ;
    buf_clk cell_4522 ( .C (CLK), .D (signal_6665), .Q (signal_6666) ) ;
    buf_clk cell_4538 ( .C (CLK), .D (signal_6681), .Q (signal_6682) ) ;
    buf_clk cell_4548 ( .C (CLK), .D (signal_6691), .Q (signal_6692) ) ;
    buf_clk cell_4558 ( .C (CLK), .D (signal_6701), .Q (signal_6702) ) ;
    buf_clk cell_4566 ( .C (CLK), .D (signal_6709), .Q (signal_6710) ) ;
    buf_clk cell_4574 ( .C (CLK), .D (signal_6717), .Q (signal_6718) ) ;
    buf_clk cell_4586 ( .C (CLK), .D (signal_6729), .Q (signal_6730) ) ;
    buf_clk cell_4598 ( .C (CLK), .D (signal_6741), .Q (signal_6742) ) ;
    buf_clk cell_4612 ( .C (CLK), .D (signal_6755), .Q (signal_6756) ) ;
    buf_clk cell_4626 ( .C (CLK), .D (signal_6769), .Q (signal_6770) ) ;
    buf_clk cell_4642 ( .C (CLK), .D (signal_6785), .Q (signal_6786) ) ;
    buf_clk cell_4658 ( .C (CLK), .D (signal_6801), .Q (signal_6802) ) ;
    buf_clk cell_4664 ( .C (CLK), .D (signal_6807), .Q (signal_6808) ) ;
    buf_clk cell_4670 ( .C (CLK), .D (signal_6813), .Q (signal_6814) ) ;
    buf_clk cell_4678 ( .C (CLK), .D (signal_6821), .Q (signal_6822) ) ;
    buf_clk cell_4686 ( .C (CLK), .D (signal_6829), .Q (signal_6830) ) ;
    buf_clk cell_4696 ( .C (CLK), .D (signal_6839), .Q (signal_6840) ) ;
    buf_clk cell_4706 ( .C (CLK), .D (signal_6849), .Q (signal_6850) ) ;
    buf_clk cell_4718 ( .C (CLK), .D (signal_6861), .Q (signal_6862) ) ;
    buf_clk cell_4730 ( .C (CLK), .D (signal_6873), .Q (signal_6874) ) ;
    buf_clk cell_4738 ( .C (CLK), .D (signal_6881), .Q (signal_6882) ) ;
    buf_clk cell_4754 ( .C (CLK), .D (signal_6897), .Q (signal_6898) ) ;
    buf_clk cell_4770 ( .C (CLK), .D (signal_6913), .Q (signal_6914) ) ;
    buf_clk cell_4786 ( .C (CLK), .D (signal_6929), .Q (signal_6930) ) ;
    buf_clk cell_4802 ( .C (CLK), .D (signal_6945), .Q (signal_6946) ) ;
    buf_clk cell_4818 ( .C (CLK), .D (signal_6961), .Q (signal_6962) ) ;
    buf_clk cell_4834 ( .C (CLK), .D (signal_6977), .Q (signal_6978) ) ;
    buf_clk cell_4850 ( .C (CLK), .D (signal_6993), .Q (signal_6994) ) ;
    buf_clk cell_4866 ( .C (CLK), .D (signal_7009), .Q (signal_7010) ) ;
    buf_clk cell_4882 ( .C (CLK), .D (signal_7025), .Q (signal_7026) ) ;
    buf_clk cell_4898 ( .C (CLK), .D (signal_7041), .Q (signal_7042) ) ;
    buf_clk cell_4914 ( .C (CLK), .D (signal_7057), .Q (signal_7058) ) ;
    buf_clk cell_4930 ( .C (CLK), .D (signal_7073), .Q (signal_7074) ) ;
    buf_clk cell_4946 ( .C (CLK), .D (signal_7089), .Q (signal_7090) ) ;
    buf_clk cell_4962 ( .C (CLK), .D (signal_7105), .Q (signal_7106) ) ;
    buf_clk cell_4978 ( .C (CLK), .D (signal_7121), .Q (signal_7122) ) ;
    buf_clk cell_4994 ( .C (CLK), .D (signal_7137), .Q (signal_7138) ) ;
    buf_clk cell_5010 ( .C (CLK), .D (signal_7153), .Q (signal_7154) ) ;
    buf_clk cell_5026 ( .C (CLK), .D (signal_7169), .Q (signal_7170) ) ;
    buf_clk cell_5042 ( .C (CLK), .D (signal_7185), .Q (signal_7186) ) ;
    buf_clk cell_5058 ( .C (CLK), .D (signal_7201), .Q (signal_7202) ) ;
    buf_clk cell_5074 ( .C (CLK), .D (signal_7217), .Q (signal_7218) ) ;
    buf_clk cell_5090 ( .C (CLK), .D (signal_7233), .Q (signal_7234) ) ;
    buf_clk cell_5106 ( .C (CLK), .D (signal_7249), .Q (signal_7250) ) ;
    buf_clk cell_5122 ( .C (CLK), .D (signal_7265), .Q (signal_7266) ) ;
    buf_clk cell_5138 ( .C (CLK), .D (signal_7281), .Q (signal_7282) ) ;
    buf_clk cell_5154 ( .C (CLK), .D (signal_7297), .Q (signal_7298) ) ;
    buf_clk cell_5170 ( .C (CLK), .D (signal_7313), .Q (signal_7314) ) ;
    buf_clk cell_5186 ( .C (CLK), .D (signal_7329), .Q (signal_7330) ) ;
    buf_clk cell_5202 ( .C (CLK), .D (signal_7345), .Q (signal_7346) ) ;
    buf_clk cell_5218 ( .C (CLK), .D (signal_7361), .Q (signal_7362) ) ;
    buf_clk cell_5234 ( .C (CLK), .D (signal_7377), .Q (signal_7378) ) ;
    buf_clk cell_5250 ( .C (CLK), .D (signal_7393), .Q (signal_7394) ) ;
    buf_clk cell_5266 ( .C (CLK), .D (signal_7409), .Q (signal_7410) ) ;
    buf_clk cell_5282 ( .C (CLK), .D (signal_7425), .Q (signal_7426) ) ;
    buf_clk cell_5298 ( .C (CLK), .D (signal_7441), .Q (signal_7442) ) ;
    buf_clk cell_5314 ( .C (CLK), .D (signal_7457), .Q (signal_7458) ) ;
    buf_clk cell_5330 ( .C (CLK), .D (signal_7473), .Q (signal_7474) ) ;
    buf_clk cell_5346 ( .C (CLK), .D (signal_7489), .Q (signal_7490) ) ;
    buf_clk cell_5362 ( .C (CLK), .D (signal_7505), .Q (signal_7506) ) ;
    buf_clk cell_5378 ( .C (CLK), .D (signal_7521), .Q (signal_7522) ) ;
    buf_clk cell_5394 ( .C (CLK), .D (signal_7537), .Q (signal_7538) ) ;
    buf_clk cell_5410 ( .C (CLK), .D (signal_7553), .Q (signal_7554) ) ;
    buf_clk cell_5426 ( .C (CLK), .D (signal_7569), .Q (signal_7570) ) ;
    buf_clk cell_5442 ( .C (CLK), .D (signal_7585), .Q (signal_7586) ) ;
    buf_clk cell_5458 ( .C (CLK), .D (signal_7601), .Q (signal_7602) ) ;
    buf_clk cell_5474 ( .C (CLK), .D (signal_7617), .Q (signal_7618) ) ;
    buf_clk cell_5490 ( .C (CLK), .D (signal_7633), .Q (signal_7634) ) ;
    buf_clk cell_5506 ( .C (CLK), .D (signal_7649), .Q (signal_7650) ) ;
    buf_clk cell_5522 ( .C (CLK), .D (signal_7665), .Q (signal_7666) ) ;
    buf_clk cell_5538 ( .C (CLK), .D (signal_7681), .Q (signal_7682) ) ;
    buf_clk cell_5554 ( .C (CLK), .D (signal_7697), .Q (signal_7698) ) ;
    buf_clk cell_5570 ( .C (CLK), .D (signal_7713), .Q (signal_7714) ) ;
    buf_clk cell_5586 ( .C (CLK), .D (signal_7729), .Q (signal_7730) ) ;
    buf_clk cell_5602 ( .C (CLK), .D (signal_7745), .Q (signal_7746) ) ;
    buf_clk cell_5618 ( .C (CLK), .D (signal_7761), .Q (signal_7762) ) ;
    buf_clk cell_5634 ( .C (CLK), .D (signal_7777), .Q (signal_7778) ) ;
    buf_clk cell_5650 ( .C (CLK), .D (signal_7793), .Q (signal_7794) ) ;
    buf_clk cell_5666 ( .C (CLK), .D (signal_7809), .Q (signal_7810) ) ;
    buf_clk cell_5682 ( .C (CLK), .D (signal_7825), .Q (signal_7826) ) ;
    buf_clk cell_5698 ( .C (CLK), .D (signal_7841), .Q (signal_7842) ) ;
    buf_clk cell_5714 ( .C (CLK), .D (signal_7857), .Q (signal_7858) ) ;
    buf_clk cell_5730 ( .C (CLK), .D (signal_7873), .Q (signal_7874) ) ;
    buf_clk cell_5746 ( .C (CLK), .D (signal_7889), .Q (signal_7890) ) ;
    buf_clk cell_5762 ( .C (CLK), .D (signal_7905), .Q (signal_7906) ) ;
    buf_clk cell_5778 ( .C (CLK), .D (signal_7921), .Q (signal_7922) ) ;
    buf_clk cell_5794 ( .C (CLK), .D (signal_7937), .Q (signal_7938) ) ;
    buf_clk cell_5810 ( .C (CLK), .D (signal_7953), .Q (signal_7954) ) ;
    buf_clk cell_5826 ( .C (CLK), .D (signal_7969), .Q (signal_7970) ) ;
    buf_clk cell_5842 ( .C (CLK), .D (signal_7985), .Q (signal_7986) ) ;
    buf_clk cell_5858 ( .C (CLK), .D (signal_8001), .Q (signal_8002) ) ;
    buf_clk cell_5874 ( .C (CLK), .D (signal_8017), .Q (signal_8018) ) ;
    buf_clk cell_5890 ( .C (CLK), .D (signal_8033), .Q (signal_8034) ) ;
    buf_clk cell_5906 ( .C (CLK), .D (signal_8049), .Q (signal_8050) ) ;
    buf_clk cell_5922 ( .C (CLK), .D (signal_8065), .Q (signal_8066) ) ;
    buf_clk cell_5938 ( .C (CLK), .D (signal_8081), .Q (signal_8082) ) ;
    buf_clk cell_5954 ( .C (CLK), .D (signal_8097), .Q (signal_8098) ) ;
    buf_clk cell_5970 ( .C (CLK), .D (signal_8113), .Q (signal_8114) ) ;
    buf_clk cell_5986 ( .C (CLK), .D (signal_8129), .Q (signal_8130) ) ;
    buf_clk cell_6002 ( .C (CLK), .D (signal_8145), .Q (signal_8146) ) ;
    buf_clk cell_6018 ( .C (CLK), .D (signal_8161), .Q (signal_8162) ) ;
    buf_clk cell_6034 ( .C (CLK), .D (signal_8177), .Q (signal_8178) ) ;
    buf_clk cell_6050 ( .C (CLK), .D (signal_8193), .Q (signal_8194) ) ;
    buf_clk cell_6066 ( .C (CLK), .D (signal_8209), .Q (signal_8210) ) ;
    buf_clk cell_6082 ( .C (CLK), .D (signal_8225), .Q (signal_8226) ) ;
    buf_clk cell_6098 ( .C (CLK), .D (signal_8241), .Q (signal_8242) ) ;
    buf_clk cell_6114 ( .C (CLK), .D (signal_8257), .Q (signal_8258) ) ;
    buf_clk cell_6130 ( .C (CLK), .D (signal_8273), .Q (signal_8274) ) ;
    buf_clk cell_6146 ( .C (CLK), .D (signal_8289), .Q (signal_8290) ) ;
    buf_clk cell_6162 ( .C (CLK), .D (signal_8305), .Q (signal_8306) ) ;
    buf_clk cell_6178 ( .C (CLK), .D (signal_8321), .Q (signal_8322) ) ;
    buf_clk cell_6194 ( .C (CLK), .D (signal_8337), .Q (signal_8338) ) ;
    buf_clk cell_6210 ( .C (CLK), .D (signal_8353), .Q (signal_8354) ) ;
    buf_clk cell_6226 ( .C (CLK), .D (signal_8369), .Q (signal_8370) ) ;
    buf_clk cell_6242 ( .C (CLK), .D (signal_8385), .Q (signal_8386) ) ;
    buf_clk cell_6258 ( .C (CLK), .D (signal_8401), .Q (signal_8402) ) ;
    buf_clk cell_6274 ( .C (CLK), .D (signal_8417), .Q (signal_8418) ) ;
    buf_clk cell_6290 ( .C (CLK), .D (signal_8433), .Q (signal_8434) ) ;
    buf_clk cell_6306 ( .C (CLK), .D (signal_8449), .Q (signal_8450) ) ;
    buf_clk cell_6322 ( .C (CLK), .D (signal_8465), .Q (signal_8466) ) ;
    buf_clk cell_6338 ( .C (CLK), .D (signal_8481), .Q (signal_8482) ) ;
    buf_clk cell_6354 ( .C (CLK), .D (signal_8497), .Q (signal_8498) ) ;
    buf_clk cell_6370 ( .C (CLK), .D (signal_8513), .Q (signal_8514) ) ;
    buf_clk cell_6386 ( .C (CLK), .D (signal_8529), .Q (signal_8530) ) ;
    buf_clk cell_6402 ( .C (CLK), .D (signal_8545), .Q (signal_8546) ) ;
    buf_clk cell_6410 ( .C (CLK), .D (signal_8553), .Q (signal_8554) ) ;
    buf_clk cell_6418 ( .C (CLK), .D (signal_8561), .Q (signal_8562) ) ;
    buf_clk cell_6426 ( .C (CLK), .D (signal_8569), .Q (signal_8570) ) ;
    buf_clk cell_6434 ( .C (CLK), .D (signal_8577), .Q (signal_8578) ) ;
    buf_clk cell_6442 ( .C (CLK), .D (signal_8585), .Q (signal_8586) ) ;
    buf_clk cell_6450 ( .C (CLK), .D (signal_8593), .Q (signal_8594) ) ;
    buf_clk cell_6458 ( .C (CLK), .D (signal_8601), .Q (signal_8602) ) ;
    buf_clk cell_6466 ( .C (CLK), .D (signal_8609), .Q (signal_8610) ) ;
    buf_clk cell_6474 ( .C (CLK), .D (signal_8617), .Q (signal_8618) ) ;
    buf_clk cell_6482 ( .C (CLK), .D (signal_8625), .Q (signal_8626) ) ;
    buf_clk cell_6490 ( .C (CLK), .D (signal_8633), .Q (signal_8634) ) ;
    buf_clk cell_6498 ( .C (CLK), .D (signal_8641), .Q (signal_8642) ) ;
    buf_clk cell_6506 ( .C (CLK), .D (signal_8649), .Q (signal_8650) ) ;
    buf_clk cell_6514 ( .C (CLK), .D (signal_8657), .Q (signal_8658) ) ;
    buf_clk cell_6522 ( .C (CLK), .D (signal_8665), .Q (signal_8666) ) ;
    buf_clk cell_6530 ( .C (CLK), .D (signal_8673), .Q (signal_8674) ) ;
    buf_clk cell_6538 ( .C (CLK), .D (signal_8681), .Q (signal_8682) ) ;
    buf_clk cell_6546 ( .C (CLK), .D (signal_8689), .Q (signal_8690) ) ;
    buf_clk cell_6554 ( .C (CLK), .D (signal_8697), .Q (signal_8698) ) ;
    buf_clk cell_6562 ( .C (CLK), .D (signal_8705), .Q (signal_8706) ) ;
    buf_clk cell_6570 ( .C (CLK), .D (signal_8713), .Q (signal_8714) ) ;
    buf_clk cell_6578 ( .C (CLK), .D (signal_8721), .Q (signal_8722) ) ;
    buf_clk cell_6586 ( .C (CLK), .D (signal_8729), .Q (signal_8730) ) ;
    buf_clk cell_6594 ( .C (CLK), .D (signal_8737), .Q (signal_8738) ) ;
    buf_clk cell_6602 ( .C (CLK), .D (signal_8745), .Q (signal_8746) ) ;
    buf_clk cell_6610 ( .C (CLK), .D (signal_8753), .Q (signal_8754) ) ;
    buf_clk cell_6618 ( .C (CLK), .D (signal_8761), .Q (signal_8762) ) ;
    buf_clk cell_6626 ( .C (CLK), .D (signal_8769), .Q (signal_8770) ) ;
    buf_clk cell_6634 ( .C (CLK), .D (signal_8777), .Q (signal_8778) ) ;
    buf_clk cell_6642 ( .C (CLK), .D (signal_8785), .Q (signal_8786) ) ;
    buf_clk cell_6650 ( .C (CLK), .D (signal_8793), .Q (signal_8794) ) ;
    buf_clk cell_6658 ( .C (CLK), .D (signal_8801), .Q (signal_8802) ) ;
    buf_clk cell_6666 ( .C (CLK), .D (signal_8809), .Q (signal_8810) ) ;
    buf_clk cell_6674 ( .C (CLK), .D (signal_8817), .Q (signal_8818) ) ;
    buf_clk cell_6682 ( .C (CLK), .D (signal_8825), .Q (signal_8826) ) ;
    buf_clk cell_6690 ( .C (CLK), .D (signal_8833), .Q (signal_8834) ) ;
    buf_clk cell_6698 ( .C (CLK), .D (signal_8841), .Q (signal_8842) ) ;
    buf_clk cell_6706 ( .C (CLK), .D (signal_8849), .Q (signal_8850) ) ;
    buf_clk cell_6714 ( .C (CLK), .D (signal_8857), .Q (signal_8858) ) ;
    buf_clk cell_6722 ( .C (CLK), .D (signal_8865), .Q (signal_8866) ) ;
    buf_clk cell_6730 ( .C (CLK), .D (signal_8873), .Q (signal_8874) ) ;
    buf_clk cell_6738 ( .C (CLK), .D (signal_8881), .Q (signal_8882) ) ;
    buf_clk cell_6746 ( .C (CLK), .D (signal_8889), .Q (signal_8890) ) ;
    buf_clk cell_6754 ( .C (CLK), .D (signal_8897), .Q (signal_8898) ) ;
    buf_clk cell_6762 ( .C (CLK), .D (signal_8905), .Q (signal_8906) ) ;
    buf_clk cell_6770 ( .C (CLK), .D (signal_8913), .Q (signal_8914) ) ;
    buf_clk cell_6778 ( .C (CLK), .D (signal_8921), .Q (signal_8922) ) ;
    buf_clk cell_6786 ( .C (CLK), .D (signal_8929), .Q (signal_8930) ) ;
    buf_clk cell_6794 ( .C (CLK), .D (signal_8937), .Q (signal_8938) ) ;
    buf_clk cell_6802 ( .C (CLK), .D (signal_8945), .Q (signal_8946) ) ;
    buf_clk cell_6810 ( .C (CLK), .D (signal_8953), .Q (signal_8954) ) ;
    buf_clk cell_6818 ( .C (CLK), .D (signal_8961), .Q (signal_8962) ) ;
    buf_clk cell_6826 ( .C (CLK), .D (signal_8969), .Q (signal_8970) ) ;
    buf_clk cell_6834 ( .C (CLK), .D (signal_8977), .Q (signal_8978) ) ;
    buf_clk cell_6842 ( .C (CLK), .D (signal_8985), .Q (signal_8986) ) ;
    buf_clk cell_6850 ( .C (CLK), .D (signal_8993), .Q (signal_8994) ) ;
    buf_clk cell_6858 ( .C (CLK), .D (signal_9001), .Q (signal_9002) ) ;
    buf_clk cell_6866 ( .C (CLK), .D (signal_9009), .Q (signal_9010) ) ;
    buf_clk cell_6874 ( .C (CLK), .D (signal_9017), .Q (signal_9018) ) ;
    buf_clk cell_6882 ( .C (CLK), .D (signal_9025), .Q (signal_9026) ) ;
    buf_clk cell_6890 ( .C (CLK), .D (signal_9033), .Q (signal_9034) ) ;
    buf_clk cell_6898 ( .C (CLK), .D (signal_9041), .Q (signal_9042) ) ;
    buf_clk cell_6906 ( .C (CLK), .D (signal_9049), .Q (signal_9050) ) ;
    buf_clk cell_6914 ( .C (CLK), .D (signal_9057), .Q (signal_9058) ) ;
    buf_clk cell_6922 ( .C (CLK), .D (signal_9065), .Q (signal_9066) ) ;
    buf_clk cell_6930 ( .C (CLK), .D (signal_9073), .Q (signal_9074) ) ;
    buf_clk cell_6938 ( .C (CLK), .D (signal_9081), .Q (signal_9082) ) ;
    buf_clk cell_6946 ( .C (CLK), .D (signal_9089), .Q (signal_9090) ) ;
    buf_clk cell_6954 ( .C (CLK), .D (signal_9097), .Q (signal_9098) ) ;
    buf_clk cell_6962 ( .C (CLK), .D (signal_9105), .Q (signal_9106) ) ;
    buf_clk cell_6970 ( .C (CLK), .D (signal_9113), .Q (signal_9114) ) ;
    buf_clk cell_6978 ( .C (CLK), .D (signal_9121), .Q (signal_9122) ) ;
    buf_clk cell_6986 ( .C (CLK), .D (signal_9129), .Q (signal_9130) ) ;
    buf_clk cell_6994 ( .C (CLK), .D (signal_9137), .Q (signal_9138) ) ;
    buf_clk cell_7002 ( .C (CLK), .D (signal_9145), .Q (signal_9146) ) ;
    buf_clk cell_7010 ( .C (CLK), .D (signal_9153), .Q (signal_9154) ) ;
    buf_clk cell_7018 ( .C (CLK), .D (signal_9161), .Q (signal_9162) ) ;
    buf_clk cell_7026 ( .C (CLK), .D (signal_9169), .Q (signal_9170) ) ;
    buf_clk cell_7034 ( .C (CLK), .D (signal_9177), .Q (signal_9178) ) ;
    buf_clk cell_7042 ( .C (CLK), .D (signal_9185), .Q (signal_9186) ) ;
    buf_clk cell_7050 ( .C (CLK), .D (signal_9193), .Q (signal_9194) ) ;
    buf_clk cell_7058 ( .C (CLK), .D (signal_9201), .Q (signal_9202) ) ;
    buf_clk cell_7066 ( .C (CLK), .D (signal_9209), .Q (signal_9210) ) ;
    buf_clk cell_7074 ( .C (CLK), .D (signal_9217), .Q (signal_9218) ) ;
    buf_clk cell_7082 ( .C (CLK), .D (signal_9225), .Q (signal_9226) ) ;
    buf_clk cell_7090 ( .C (CLK), .D (signal_9233), .Q (signal_9234) ) ;
    buf_clk cell_7098 ( .C (CLK), .D (signal_9241), .Q (signal_9242) ) ;
    buf_clk cell_7106 ( .C (CLK), .D (signal_9249), .Q (signal_9250) ) ;
    buf_clk cell_7114 ( .C (CLK), .D (signal_9257), .Q (signal_9258) ) ;
    buf_clk cell_7122 ( .C (CLK), .D (signal_9265), .Q (signal_9266) ) ;
    buf_clk cell_7130 ( .C (CLK), .D (signal_9273), .Q (signal_9274) ) ;
    buf_clk cell_7138 ( .C (CLK), .D (signal_9281), .Q (signal_9282) ) ;
    buf_clk cell_7146 ( .C (CLK), .D (signal_9289), .Q (signal_9290) ) ;
    buf_clk cell_7154 ( .C (CLK), .D (signal_9297), .Q (signal_9298) ) ;
    buf_clk cell_7162 ( .C (CLK), .D (signal_9305), .Q (signal_9306) ) ;
    buf_clk cell_7170 ( .C (CLK), .D (signal_9313), .Q (signal_9314) ) ;
    buf_clk cell_7178 ( .C (CLK), .D (signal_9321), .Q (signal_9322) ) ;
    buf_clk cell_7186 ( .C (CLK), .D (signal_9329), .Q (signal_9330) ) ;
    buf_clk cell_7194 ( .C (CLK), .D (signal_9337), .Q (signal_9338) ) ;
    buf_clk cell_7202 ( .C (CLK), .D (signal_9345), .Q (signal_9346) ) ;
    buf_clk cell_7210 ( .C (CLK), .D (signal_9353), .Q (signal_9354) ) ;
    buf_clk cell_7218 ( .C (CLK), .D (signal_9361), .Q (signal_9362) ) ;
    buf_clk cell_7226 ( .C (CLK), .D (signal_9369), .Q (signal_9370) ) ;
    buf_clk cell_7234 ( .C (CLK), .D (signal_9377), .Q (signal_9378) ) ;
    buf_clk cell_7242 ( .C (CLK), .D (signal_9385), .Q (signal_9386) ) ;
    buf_clk cell_7250 ( .C (CLK), .D (signal_9393), .Q (signal_9394) ) ;
    buf_clk cell_7258 ( .C (CLK), .D (signal_9401), .Q (signal_9402) ) ;
    buf_clk cell_7266 ( .C (CLK), .D (signal_9409), .Q (signal_9410) ) ;
    buf_clk cell_7274 ( .C (CLK), .D (signal_9417), .Q (signal_9418) ) ;
    buf_clk cell_7282 ( .C (CLK), .D (signal_9425), .Q (signal_9426) ) ;
    buf_clk cell_7290 ( .C (CLK), .D (signal_9433), .Q (signal_9434) ) ;
    buf_clk cell_7298 ( .C (CLK), .D (signal_9441), .Q (signal_9442) ) ;
    buf_clk cell_7306 ( .C (CLK), .D (signal_9449), .Q (signal_9450) ) ;
    buf_clk cell_7314 ( .C (CLK), .D (signal_9457), .Q (signal_9458) ) ;
    buf_clk cell_7322 ( .C (CLK), .D (signal_9465), .Q (signal_9466) ) ;
    buf_clk cell_7330 ( .C (CLK), .D (signal_9473), .Q (signal_9474) ) ;
    buf_clk cell_7338 ( .C (CLK), .D (signal_9481), .Q (signal_9482) ) ;
    buf_clk cell_7346 ( .C (CLK), .D (signal_9489), .Q (signal_9490) ) ;
    buf_clk cell_7354 ( .C (CLK), .D (signal_9497), .Q (signal_9498) ) ;
    buf_clk cell_7362 ( .C (CLK), .D (signal_9505), .Q (signal_9506) ) ;
    buf_clk cell_7370 ( .C (CLK), .D (signal_9513), .Q (signal_9514) ) ;
    buf_clk cell_7378 ( .C (CLK), .D (signal_9521), .Q (signal_9522) ) ;
    buf_clk cell_7386 ( .C (CLK), .D (signal_9529), .Q (signal_9530) ) ;
    buf_clk cell_7394 ( .C (CLK), .D (signal_9537), .Q (signal_9538) ) ;
    buf_clk cell_7402 ( .C (CLK), .D (signal_9545), .Q (signal_9546) ) ;
    buf_clk cell_7410 ( .C (CLK), .D (signal_9553), .Q (signal_9554) ) ;
    buf_clk cell_7418 ( .C (CLK), .D (signal_9561), .Q (signal_9562) ) ;
    buf_clk cell_7426 ( .C (CLK), .D (signal_9569), .Q (signal_9570) ) ;
    buf_clk cell_7434 ( .C (CLK), .D (signal_9577), .Q (signal_9578) ) ;
    buf_clk cell_7442 ( .C (CLK), .D (signal_9585), .Q (signal_9586) ) ;
    buf_clk cell_7450 ( .C (CLK), .D (signal_9593), .Q (signal_9594) ) ;
    buf_clk cell_7458 ( .C (CLK), .D (signal_9601), .Q (signal_9602) ) ;
    buf_clk cell_7466 ( .C (CLK), .D (signal_9609), .Q (signal_9610) ) ;
    buf_clk cell_7474 ( .C (CLK), .D (signal_9617), .Q (signal_9618) ) ;
    buf_clk cell_7482 ( .C (CLK), .D (signal_9625), .Q (signal_9626) ) ;
    buf_clk cell_7490 ( .C (CLK), .D (signal_9633), .Q (signal_9634) ) ;
    buf_clk cell_7498 ( .C (CLK), .D (signal_9641), .Q (signal_9642) ) ;
    buf_clk cell_7506 ( .C (CLK), .D (signal_9649), .Q (signal_9650) ) ;
    buf_clk cell_7514 ( .C (CLK), .D (signal_9657), .Q (signal_9658) ) ;
    buf_clk cell_7522 ( .C (CLK), .D (signal_9665), .Q (signal_9666) ) ;
    buf_clk cell_7530 ( .C (CLK), .D (signal_9673), .Q (signal_9674) ) ;
    buf_clk cell_7538 ( .C (CLK), .D (signal_9681), .Q (signal_9682) ) ;
    buf_clk cell_7546 ( .C (CLK), .D (signal_9689), .Q (signal_9690) ) ;
    buf_clk cell_7554 ( .C (CLK), .D (signal_9697), .Q (signal_9698) ) ;
    buf_clk cell_7558 ( .C (CLK), .D (signal_5447), .Q (signal_9702) ) ;
    buf_clk cell_7560 ( .C (CLK), .D (signal_5453), .Q (signal_9704) ) ;
    buf_clk cell_7568 ( .C (CLK), .D (signal_9711), .Q (signal_9712) ) ;
    buf_clk cell_7576 ( .C (CLK), .D (signal_9719), .Q (signal_9720) ) ;
    buf_clk cell_7580 ( .C (CLK), .D (signal_9723), .Q (signal_9724) ) ;
    buf_clk cell_7584 ( .C (CLK), .D (signal_9727), .Q (signal_9728) ) ;
    buf_clk cell_7586 ( .C (CLK), .D (signal_5487), .Q (signal_9730) ) ;
    buf_clk cell_7588 ( .C (CLK), .D (signal_5493), .Q (signal_9732) ) ;
    buf_clk cell_7602 ( .C (CLK), .D (signal_9745), .Q (signal_9746) ) ;
    buf_clk cell_7618 ( .C (CLK), .D (signal_9761), .Q (signal_9762) ) ;
    buf_clk cell_7634 ( .C (CLK), .D (signal_9777), .Q (signal_9778) ) ;
    buf_clk cell_7650 ( .C (CLK), .D (signal_9793), .Q (signal_9794) ) ;
    buf_clk cell_7666 ( .C (CLK), .D (signal_9809), .Q (signal_9810) ) ;
    buf_clk cell_7682 ( .C (CLK), .D (signal_9825), .Q (signal_9826) ) ;
    buf_clk cell_7698 ( .C (CLK), .D (signal_9841), .Q (signal_9842) ) ;
    buf_clk cell_7714 ( .C (CLK), .D (signal_9857), .Q (signal_9858) ) ;
    buf_clk cell_7730 ( .C (CLK), .D (signal_9873), .Q (signal_9874) ) ;
    buf_clk cell_7746 ( .C (CLK), .D (signal_9889), .Q (signal_9890) ) ;
    buf_clk cell_7754 ( .C (CLK), .D (signal_9897), .Q (signal_9898) ) ;
    buf_clk cell_7762 ( .C (CLK), .D (signal_9905), .Q (signal_9906) ) ;
    buf_clk cell_7770 ( .C (CLK), .D (signal_9913), .Q (signal_9914) ) ;
    buf_clk cell_7778 ( .C (CLK), .D (signal_9921), .Q (signal_9922) ) ;
    buf_clk cell_7786 ( .C (CLK), .D (signal_9929), .Q (signal_9930) ) ;
    buf_clk cell_7794 ( .C (CLK), .D (signal_9937), .Q (signal_9938) ) ;
    buf_clk cell_7802 ( .C (CLK), .D (signal_9945), .Q (signal_9946) ) ;
    buf_clk cell_7810 ( .C (CLK), .D (signal_9953), .Q (signal_9954) ) ;
    buf_clk cell_7818 ( .C (CLK), .D (signal_9961), .Q (signal_9962) ) ;
    buf_clk cell_7826 ( .C (CLK), .D (signal_9969), .Q (signal_9970) ) ;
    buf_clk cell_7834 ( .C (CLK), .D (signal_9977), .Q (signal_9978) ) ;
    buf_clk cell_7842 ( .C (CLK), .D (signal_9985), .Q (signal_9986) ) ;
    buf_clk cell_7850 ( .C (CLK), .D (signal_9993), .Q (signal_9994) ) ;
    buf_clk cell_7858 ( .C (CLK), .D (signal_10001), .Q (signal_10002) ) ;
    buf_clk cell_7866 ( .C (CLK), .D (signal_10009), .Q (signal_10010) ) ;
    buf_clk cell_7874 ( .C (CLK), .D (signal_10017), .Q (signal_10018) ) ;
    buf_clk cell_7882 ( .C (CLK), .D (signal_10025), .Q (signal_10026) ) ;
    buf_clk cell_7890 ( .C (CLK), .D (signal_10033), .Q (signal_10034) ) ;
    buf_clk cell_7898 ( .C (CLK), .D (signal_10041), .Q (signal_10042) ) ;
    buf_clk cell_7906 ( .C (CLK), .D (signal_10049), .Q (signal_10050) ) ;
    buf_clk cell_7914 ( .C (CLK), .D (signal_10057), .Q (signal_10058) ) ;
    buf_clk cell_7922 ( .C (CLK), .D (signal_10065), .Q (signal_10066) ) ;
    buf_clk cell_7930 ( .C (CLK), .D (signal_10073), .Q (signal_10074) ) ;
    buf_clk cell_7938 ( .C (CLK), .D (signal_10081), .Q (signal_10082) ) ;
    buf_clk cell_7954 ( .C (CLK), .D (signal_10097), .Q (signal_10098) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1678 ( .s ({signal_5425, signal_5421}), .b ({signal_5429, signal_5427}), .a ({signal_2803, signal_1778}), .clk (CLK), .r (Fresh[550]), .c ({signal_2870, signal_1822}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1679 ( .s ({signal_5425, signal_5421}), .b ({signal_2805, signal_1780}), .a ({signal_2804, signal_1779}), .clk (CLK), .r (Fresh[551]), .c ({signal_2871, signal_1823}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1680 ( .s ({signal_5437, signal_5433}), .b ({signal_2838, signal_1781}), .a ({signal_5441, signal_5439}), .clk (CLK), .r (Fresh[552]), .c ({signal_2890, signal_1824}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1681 ( .s ({signal_5437, signal_5433}), .b ({signal_2840, signal_1783}), .a ({signal_2839, signal_1782}), .clk (CLK), .r (Fresh[553]), .c ({signal_2891, signal_1825}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1682 ( .s ({signal_5453, signal_5447}), .b ({signal_5457, signal_5455}), .a ({signal_2841, signal_1784}), .clk (CLK), .r (Fresh[554]), .c ({signal_2892, signal_1826}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1683 ( .s ({signal_5453, signal_5447}), .b ({signal_5461, signal_5459}), .a ({signal_2842, signal_1785}), .clk (CLK), .r (Fresh[555]), .c ({signal_2893, signal_1827}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1684 ( .s ({signal_5477, signal_5469}), .b ({signal_2844, signal_1787}), .a ({signal_2843, signal_1786}), .clk (CLK), .r (Fresh[556]), .c ({signal_2894, signal_1828}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1685 ( .s ({signal_5477, signal_5469}), .b ({signal_2845, signal_1788}), .a ({signal_5481, signal_5479}), .clk (CLK), .r (Fresh[557]), .c ({signal_2895, signal_1829}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1686 ( .s ({signal_5493, signal_5487}), .b ({signal_2847, signal_1790}), .a ({signal_2846, signal_1789}), .clk (CLK), .r (Fresh[558]), .c ({signal_2896, signal_1830}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1687 ( .s ({signal_5493, signal_5487}), .b ({signal_2849, signal_1792}), .a ({signal_2848, signal_1791}), .clk (CLK), .r (Fresh[559]), .c ({signal_2897, signal_1831}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1688 ( .s ({signal_5497, signal_5495}), .b ({signal_2851, signal_1794}), .a ({signal_2850, signal_1793}), .clk (CLK), .r (Fresh[560]), .c ({signal_2898, signal_1832}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1689 ( .s ({signal_5497, signal_5495}), .b ({signal_2850, signal_1793}), .a ({signal_2851, signal_1794}), .clk (CLK), .r (Fresh[561]), .c ({signal_2899, signal_1833}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1690 ( .s ({signal_5513, signal_5505}), .b ({signal_5517, signal_5515}), .a ({signal_2852, signal_1795}), .clk (CLK), .r (Fresh[562]), .c ({signal_2900, signal_1834}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1691 ( .s ({signal_5513, signal_5505}), .b ({signal_5521, signal_5519}), .a ({signal_2853, signal_1796}), .clk (CLK), .r (Fresh[563]), .c ({signal_2901, signal_1835}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1692 ( .s ({signal_5425, signal_5421}), .b ({signal_5525, signal_5523}), .a ({signal_2854, signal_1797}), .clk (CLK), .r (Fresh[564]), .c ({signal_2902, signal_1836}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1693 ( .s ({signal_5425, signal_5421}), .b ({signal_5529, signal_5527}), .a ({signal_2855, signal_1798}), .clk (CLK), .r (Fresh[565]), .c ({signal_2903, signal_1837}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1694 ( .s ({signal_5533, signal_5531}), .b ({signal_2856, signal_1799}), .a ({signal_5537, signal_5535}), .clk (CLK), .r (Fresh[566]), .c ({signal_2904, signal_1838}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1695 ( .s ({signal_5533, signal_5531}), .b ({signal_2857, signal_1800}), .a ({signal_5541, signal_5539}), .clk (CLK), .r (Fresh[567]), .c ({signal_2905, signal_1839}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1696 ( .s ({signal_5549, signal_5545}), .b ({signal_2807, signal_1802}), .a ({signal_2806, signal_1801}), .clk (CLK), .r (Fresh[568]), .c ({signal_2872, signal_1840}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1697 ( .s ({signal_5549, signal_5545}), .b ({signal_2809, signal_1804}), .a ({signal_2808, signal_1803}), .clk (CLK), .r (Fresh[569]), .c ({signal_2873, signal_1841}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1698 ( .s ({signal_5557, signal_5553}), .b ({signal_2810, signal_1805}), .a ({signal_5561, signal_5559}), .clk (CLK), .r (Fresh[570]), .c ({signal_2874, signal_1842}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1699 ( .s ({signal_5557, signal_5553}), .b ({signal_2811, signal_1806}), .a ({signal_5565, signal_5563}), .clk (CLK), .r (Fresh[571]), .c ({signal_2875, signal_1843}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1700 ( .s ({signal_5569, signal_5567}), .b ({signal_2859, signal_1808}), .a ({signal_2858, signal_1807}), .clk (CLK), .r (Fresh[572]), .c ({signal_2906, signal_1844}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1701 ( .s ({signal_5569, signal_5567}), .b ({signal_2858, signal_1807}), .a ({signal_2859, signal_1808}), .clk (CLK), .r (Fresh[573]), .c ({signal_2907, signal_1845}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1702 ( .s ({signal_5425, signal_5421}), .b ({signal_5573, signal_5571}), .a ({signal_2812, signal_1809}), .clk (CLK), .r (Fresh[574]), .c ({signal_2876, signal_1846}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1703 ( .s ({signal_5425, signal_5421}), .b ({signal_2814, signal_1811}), .a ({signal_2813, signal_1810}), .clk (CLK), .r (Fresh[575]), .c ({signal_2877, signal_1847}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1704 ( .s ({signal_5477, signal_5469}), .b ({signal_2861, signal_1813}), .a ({signal_2860, signal_1812}), .clk (CLK), .r (Fresh[576]), .c ({signal_2908, signal_1848}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1705 ( .s ({signal_5477, signal_5469}), .b ({signal_2862, signal_1814}), .a ({signal_5577, signal_5575}), .clk (CLK), .r (Fresh[577]), .c ({signal_2909, signal_1849}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1706 ( .s ({signal_5437, signal_5433}), .b ({signal_2863, signal_1815}), .a ({signal_5581, signal_5579}), .clk (CLK), .r (Fresh[578]), .c ({signal_2910, signal_1850}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1707 ( .s ({signal_5437, signal_5433}), .b ({signal_2865, signal_1817}), .a ({signal_2864, signal_1816}), .clk (CLK), .r (Fresh[579]), .c ({signal_2911, signal_1851}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1708 ( .s ({signal_5493, signal_5487}), .b ({signal_2867, signal_1819}), .a ({signal_2866, signal_1818}), .clk (CLK), .r (Fresh[580]), .c ({signal_2912, signal_1852}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1709 ( .s ({signal_5493, signal_5487}), .b ({signal_2869, signal_1821}), .a ({signal_2868, signal_1820}), .clk (CLK), .r (Fresh[581]), .c ({signal_2913, signal_1853}) ) ;
    buf_clk cell_3443 ( .C (CLK), .D (signal_5586), .Q (signal_5587) ) ;
    buf_clk cell_3459 ( .C (CLK), .D (signal_5602), .Q (signal_5603) ) ;
    buf_clk cell_3475 ( .C (CLK), .D (signal_5618), .Q (signal_5619) ) ;
    buf_clk cell_3483 ( .C (CLK), .D (signal_5626), .Q (signal_5627) ) ;
    buf_clk cell_3499 ( .C (CLK), .D (signal_5642), .Q (signal_5643) ) ;
    buf_clk cell_3515 ( .C (CLK), .D (signal_5658), .Q (signal_5659) ) ;
    buf_clk cell_3523 ( .C (CLK), .D (signal_5666), .Q (signal_5667) ) ;
    buf_clk cell_3539 ( .C (CLK), .D (signal_5682), .Q (signal_5683) ) ;
    buf_clk cell_3555 ( .C (CLK), .D (signal_5698), .Q (signal_5699) ) ;
    buf_clk cell_3571 ( .C (CLK), .D (signal_5714), .Q (signal_5715) ) ;
    buf_clk cell_3587 ( .C (CLK), .D (signal_5730), .Q (signal_5731) ) ;
    buf_clk cell_3591 ( .C (CLK), .D (signal_5734), .Q (signal_5735) ) ;
    buf_clk cell_3595 ( .C (CLK), .D (signal_5738), .Q (signal_5739) ) ;
    buf_clk cell_3601 ( .C (CLK), .D (signal_5744), .Q (signal_5745) ) ;
    buf_clk cell_3607 ( .C (CLK), .D (signal_5750), .Q (signal_5751) ) ;
    buf_clk cell_3613 ( .C (CLK), .D (signal_5756), .Q (signal_5757) ) ;
    buf_clk cell_3619 ( .C (CLK), .D (signal_5762), .Q (signal_5763) ) ;
    buf_clk cell_3625 ( .C (CLK), .D (signal_5768), .Q (signal_5769) ) ;
    buf_clk cell_3631 ( .C (CLK), .D (signal_5774), .Q (signal_5775) ) ;
    buf_clk cell_3647 ( .C (CLK), .D (signal_5790), .Q (signal_5791) ) ;
    buf_clk cell_3663 ( .C (CLK), .D (signal_5806), .Q (signal_5807) ) ;
    buf_clk cell_3679 ( .C (CLK), .D (signal_5822), .Q (signal_5823) ) ;
    buf_clk cell_3695 ( .C (CLK), .D (signal_5838), .Q (signal_5839) ) ;
    buf_clk cell_3711 ( .C (CLK), .D (signal_5854), .Q (signal_5855) ) ;
    buf_clk cell_3727 ( .C (CLK), .D (signal_5870), .Q (signal_5871) ) ;
    buf_clk cell_3743 ( .C (CLK), .D (signal_5886), .Q (signal_5887) ) ;
    buf_clk cell_3759 ( .C (CLK), .D (signal_5902), .Q (signal_5903) ) ;
    buf_clk cell_3775 ( .C (CLK), .D (signal_5918), .Q (signal_5919) ) ;
    buf_clk cell_3791 ( .C (CLK), .D (signal_5934), .Q (signal_5935) ) ;
    buf_clk cell_3795 ( .C (CLK), .D (signal_5938), .Q (signal_5939) ) ;
    buf_clk cell_3799 ( .C (CLK), .D (signal_5942), .Q (signal_5943) ) ;
    buf_clk cell_3807 ( .C (CLK), .D (signal_5950), .Q (signal_5951) ) ;
    buf_clk cell_3815 ( .C (CLK), .D (signal_5958), .Q (signal_5959) ) ;
    buf_clk cell_3821 ( .C (CLK), .D (signal_5964), .Q (signal_5965) ) ;
    buf_clk cell_3827 ( .C (CLK), .D (signal_5970), .Q (signal_5971) ) ;
    buf_clk cell_3835 ( .C (CLK), .D (signal_5978), .Q (signal_5979) ) ;
    buf_clk cell_3843 ( .C (CLK), .D (signal_5986), .Q (signal_5987) ) ;
    buf_clk cell_3851 ( .C (CLK), .D (signal_5994), .Q (signal_5995) ) ;
    buf_clk cell_3859 ( .C (CLK), .D (signal_6002), .Q (signal_6003) ) ;
    buf_clk cell_3863 ( .C (CLK), .D (signal_6006), .Q (signal_6007) ) ;
    buf_clk cell_3867 ( .C (CLK), .D (signal_6010), .Q (signal_6011) ) ;
    buf_clk cell_3875 ( .C (CLK), .D (signal_6018), .Q (signal_6019) ) ;
    buf_clk cell_3883 ( .C (CLK), .D (signal_6026), .Q (signal_6027) ) ;
    buf_clk cell_3899 ( .C (CLK), .D (signal_6042), .Q (signal_6043) ) ;
    buf_clk cell_3915 ( .C (CLK), .D (signal_6058), .Q (signal_6059) ) ;
    buf_clk cell_3931 ( .C (CLK), .D (signal_6074), .Q (signal_6075) ) ;
    buf_clk cell_3947 ( .C (CLK), .D (signal_6090), .Q (signal_6091) ) ;
    buf_clk cell_3963 ( .C (CLK), .D (signal_6106), .Q (signal_6107) ) ;
    buf_clk cell_3979 ( .C (CLK), .D (signal_6122), .Q (signal_6123) ) ;
    buf_clk cell_3995 ( .C (CLK), .D (signal_6138), .Q (signal_6139) ) ;
    buf_clk cell_4011 ( .C (CLK), .D (signal_6154), .Q (signal_6155) ) ;
    buf_clk cell_4027 ( .C (CLK), .D (signal_6170), .Q (signal_6171) ) ;
    buf_clk cell_4043 ( .C (CLK), .D (signal_6186), .Q (signal_6187) ) ;
    buf_clk cell_4059 ( .C (CLK), .D (signal_6202), .Q (signal_6203) ) ;
    buf_clk cell_4075 ( .C (CLK), .D (signal_6218), .Q (signal_6219) ) ;
    buf_clk cell_4091 ( .C (CLK), .D (signal_6234), .Q (signal_6235) ) ;
    buf_clk cell_4107 ( .C (CLK), .D (signal_6250), .Q (signal_6251) ) ;
    buf_clk cell_4117 ( .C (CLK), .D (signal_6260), .Q (signal_6261) ) ;
    buf_clk cell_4127 ( .C (CLK), .D (signal_6270), .Q (signal_6271) ) ;
    buf_clk cell_4133 ( .C (CLK), .D (signal_6276), .Q (signal_6277) ) ;
    buf_clk cell_4139 ( .C (CLK), .D (signal_6282), .Q (signal_6283) ) ;
    buf_clk cell_4147 ( .C (CLK), .D (signal_6290), .Q (signal_6291) ) ;
    buf_clk cell_4155 ( .C (CLK), .D (signal_6298), .Q (signal_6299) ) ;
    buf_clk cell_4165 ( .C (CLK), .D (signal_6308), .Q (signal_6309) ) ;
    buf_clk cell_4175 ( .C (CLK), .D (signal_6318), .Q (signal_6319) ) ;
    buf_clk cell_4191 ( .C (CLK), .D (signal_6334), .Q (signal_6335) ) ;
    buf_clk cell_4203 ( .C (CLK), .D (signal_6346), .Q (signal_6347) ) ;
    buf_clk cell_4215 ( .C (CLK), .D (signal_6358), .Q (signal_6359) ) ;
    buf_clk cell_4223 ( .C (CLK), .D (signal_6366), .Q (signal_6367) ) ;
    buf_clk cell_4231 ( .C (CLK), .D (signal_6374), .Q (signal_6375) ) ;
    buf_clk cell_4243 ( .C (CLK), .D (signal_6386), .Q (signal_6387) ) ;
    buf_clk cell_4255 ( .C (CLK), .D (signal_6398), .Q (signal_6399) ) ;
    buf_clk cell_4269 ( .C (CLK), .D (signal_6412), .Q (signal_6413) ) ;
    buf_clk cell_4283 ( .C (CLK), .D (signal_6426), .Q (signal_6427) ) ;
    buf_clk cell_4299 ( .C (CLK), .D (signal_6442), .Q (signal_6443) ) ;
    buf_clk cell_4315 ( .C (CLK), .D (signal_6458), .Q (signal_6459) ) ;
    buf_clk cell_4331 ( .C (CLK), .D (signal_6474), .Q (signal_6475) ) ;
    buf_clk cell_4347 ( .C (CLK), .D (signal_6490), .Q (signal_6491) ) ;
    buf_clk cell_4363 ( .C (CLK), .D (signal_6506), .Q (signal_6507) ) ;
    buf_clk cell_4379 ( .C (CLK), .D (signal_6522), .Q (signal_6523) ) ;
    buf_clk cell_4395 ( .C (CLK), .D (signal_6538), .Q (signal_6539) ) ;
    buf_clk cell_4411 ( .C (CLK), .D (signal_6554), .Q (signal_6555) ) ;
    buf_clk cell_4427 ( .C (CLK), .D (signal_6570), .Q (signal_6571) ) ;
    buf_clk cell_4443 ( .C (CLK), .D (signal_6586), .Q (signal_6587) ) ;
    buf_clk cell_4459 ( .C (CLK), .D (signal_6602), .Q (signal_6603) ) ;
    buf_clk cell_4475 ( .C (CLK), .D (signal_6618), .Q (signal_6619) ) ;
    buf_clk cell_4491 ( .C (CLK), .D (signal_6634), .Q (signal_6635) ) ;
    buf_clk cell_4507 ( .C (CLK), .D (signal_6650), .Q (signal_6651) ) ;
    buf_clk cell_4523 ( .C (CLK), .D (signal_6666), .Q (signal_6667) ) ;
    buf_clk cell_4539 ( .C (CLK), .D (signal_6682), .Q (signal_6683) ) ;
    buf_clk cell_4549 ( .C (CLK), .D (signal_6692), .Q (signal_6693) ) ;
    buf_clk cell_4559 ( .C (CLK), .D (signal_6702), .Q (signal_6703) ) ;
    buf_clk cell_4567 ( .C (CLK), .D (signal_6710), .Q (signal_6711) ) ;
    buf_clk cell_4575 ( .C (CLK), .D (signal_6718), .Q (signal_6719) ) ;
    buf_clk cell_4587 ( .C (CLK), .D (signal_6730), .Q (signal_6731) ) ;
    buf_clk cell_4599 ( .C (CLK), .D (signal_6742), .Q (signal_6743) ) ;
    buf_clk cell_4613 ( .C (CLK), .D (signal_6756), .Q (signal_6757) ) ;
    buf_clk cell_4627 ( .C (CLK), .D (signal_6770), .Q (signal_6771) ) ;
    buf_clk cell_4643 ( .C (CLK), .D (signal_6786), .Q (signal_6787) ) ;
    buf_clk cell_4659 ( .C (CLK), .D (signal_6802), .Q (signal_6803) ) ;
    buf_clk cell_4665 ( .C (CLK), .D (signal_6808), .Q (signal_6809) ) ;
    buf_clk cell_4671 ( .C (CLK), .D (signal_6814), .Q (signal_6815) ) ;
    buf_clk cell_4679 ( .C (CLK), .D (signal_6822), .Q (signal_6823) ) ;
    buf_clk cell_4687 ( .C (CLK), .D (signal_6830), .Q (signal_6831) ) ;
    buf_clk cell_4697 ( .C (CLK), .D (signal_6840), .Q (signal_6841) ) ;
    buf_clk cell_4707 ( .C (CLK), .D (signal_6850), .Q (signal_6851) ) ;
    buf_clk cell_4719 ( .C (CLK), .D (signal_6862), .Q (signal_6863) ) ;
    buf_clk cell_4731 ( .C (CLK), .D (signal_6874), .Q (signal_6875) ) ;
    buf_clk cell_4739 ( .C (CLK), .D (signal_6882), .Q (signal_6883) ) ;
    buf_clk cell_4755 ( .C (CLK), .D (signal_6898), .Q (signal_6899) ) ;
    buf_clk cell_4771 ( .C (CLK), .D (signal_6914), .Q (signal_6915) ) ;
    buf_clk cell_4787 ( .C (CLK), .D (signal_6930), .Q (signal_6931) ) ;
    buf_clk cell_4803 ( .C (CLK), .D (signal_6946), .Q (signal_6947) ) ;
    buf_clk cell_4819 ( .C (CLK), .D (signal_6962), .Q (signal_6963) ) ;
    buf_clk cell_4835 ( .C (CLK), .D (signal_6978), .Q (signal_6979) ) ;
    buf_clk cell_4851 ( .C (CLK), .D (signal_6994), .Q (signal_6995) ) ;
    buf_clk cell_4867 ( .C (CLK), .D (signal_7010), .Q (signal_7011) ) ;
    buf_clk cell_4883 ( .C (CLK), .D (signal_7026), .Q (signal_7027) ) ;
    buf_clk cell_4899 ( .C (CLK), .D (signal_7042), .Q (signal_7043) ) ;
    buf_clk cell_4915 ( .C (CLK), .D (signal_7058), .Q (signal_7059) ) ;
    buf_clk cell_4931 ( .C (CLK), .D (signal_7074), .Q (signal_7075) ) ;
    buf_clk cell_4947 ( .C (CLK), .D (signal_7090), .Q (signal_7091) ) ;
    buf_clk cell_4963 ( .C (CLK), .D (signal_7106), .Q (signal_7107) ) ;
    buf_clk cell_4979 ( .C (CLK), .D (signal_7122), .Q (signal_7123) ) ;
    buf_clk cell_4995 ( .C (CLK), .D (signal_7138), .Q (signal_7139) ) ;
    buf_clk cell_5011 ( .C (CLK), .D (signal_7154), .Q (signal_7155) ) ;
    buf_clk cell_5027 ( .C (CLK), .D (signal_7170), .Q (signal_7171) ) ;
    buf_clk cell_5043 ( .C (CLK), .D (signal_7186), .Q (signal_7187) ) ;
    buf_clk cell_5059 ( .C (CLK), .D (signal_7202), .Q (signal_7203) ) ;
    buf_clk cell_5075 ( .C (CLK), .D (signal_7218), .Q (signal_7219) ) ;
    buf_clk cell_5091 ( .C (CLK), .D (signal_7234), .Q (signal_7235) ) ;
    buf_clk cell_5107 ( .C (CLK), .D (signal_7250), .Q (signal_7251) ) ;
    buf_clk cell_5123 ( .C (CLK), .D (signal_7266), .Q (signal_7267) ) ;
    buf_clk cell_5139 ( .C (CLK), .D (signal_7282), .Q (signal_7283) ) ;
    buf_clk cell_5155 ( .C (CLK), .D (signal_7298), .Q (signal_7299) ) ;
    buf_clk cell_5171 ( .C (CLK), .D (signal_7314), .Q (signal_7315) ) ;
    buf_clk cell_5187 ( .C (CLK), .D (signal_7330), .Q (signal_7331) ) ;
    buf_clk cell_5203 ( .C (CLK), .D (signal_7346), .Q (signal_7347) ) ;
    buf_clk cell_5219 ( .C (CLK), .D (signal_7362), .Q (signal_7363) ) ;
    buf_clk cell_5235 ( .C (CLK), .D (signal_7378), .Q (signal_7379) ) ;
    buf_clk cell_5251 ( .C (CLK), .D (signal_7394), .Q (signal_7395) ) ;
    buf_clk cell_5267 ( .C (CLK), .D (signal_7410), .Q (signal_7411) ) ;
    buf_clk cell_5283 ( .C (CLK), .D (signal_7426), .Q (signal_7427) ) ;
    buf_clk cell_5299 ( .C (CLK), .D (signal_7442), .Q (signal_7443) ) ;
    buf_clk cell_5315 ( .C (CLK), .D (signal_7458), .Q (signal_7459) ) ;
    buf_clk cell_5331 ( .C (CLK), .D (signal_7474), .Q (signal_7475) ) ;
    buf_clk cell_5347 ( .C (CLK), .D (signal_7490), .Q (signal_7491) ) ;
    buf_clk cell_5363 ( .C (CLK), .D (signal_7506), .Q (signal_7507) ) ;
    buf_clk cell_5379 ( .C (CLK), .D (signal_7522), .Q (signal_7523) ) ;
    buf_clk cell_5395 ( .C (CLK), .D (signal_7538), .Q (signal_7539) ) ;
    buf_clk cell_5411 ( .C (CLK), .D (signal_7554), .Q (signal_7555) ) ;
    buf_clk cell_5427 ( .C (CLK), .D (signal_7570), .Q (signal_7571) ) ;
    buf_clk cell_5443 ( .C (CLK), .D (signal_7586), .Q (signal_7587) ) ;
    buf_clk cell_5459 ( .C (CLK), .D (signal_7602), .Q (signal_7603) ) ;
    buf_clk cell_5475 ( .C (CLK), .D (signal_7618), .Q (signal_7619) ) ;
    buf_clk cell_5491 ( .C (CLK), .D (signal_7634), .Q (signal_7635) ) ;
    buf_clk cell_5507 ( .C (CLK), .D (signal_7650), .Q (signal_7651) ) ;
    buf_clk cell_5523 ( .C (CLK), .D (signal_7666), .Q (signal_7667) ) ;
    buf_clk cell_5539 ( .C (CLK), .D (signal_7682), .Q (signal_7683) ) ;
    buf_clk cell_5555 ( .C (CLK), .D (signal_7698), .Q (signal_7699) ) ;
    buf_clk cell_5571 ( .C (CLK), .D (signal_7714), .Q (signal_7715) ) ;
    buf_clk cell_5587 ( .C (CLK), .D (signal_7730), .Q (signal_7731) ) ;
    buf_clk cell_5603 ( .C (CLK), .D (signal_7746), .Q (signal_7747) ) ;
    buf_clk cell_5619 ( .C (CLK), .D (signal_7762), .Q (signal_7763) ) ;
    buf_clk cell_5635 ( .C (CLK), .D (signal_7778), .Q (signal_7779) ) ;
    buf_clk cell_5651 ( .C (CLK), .D (signal_7794), .Q (signal_7795) ) ;
    buf_clk cell_5667 ( .C (CLK), .D (signal_7810), .Q (signal_7811) ) ;
    buf_clk cell_5683 ( .C (CLK), .D (signal_7826), .Q (signal_7827) ) ;
    buf_clk cell_5699 ( .C (CLK), .D (signal_7842), .Q (signal_7843) ) ;
    buf_clk cell_5715 ( .C (CLK), .D (signal_7858), .Q (signal_7859) ) ;
    buf_clk cell_5731 ( .C (CLK), .D (signal_7874), .Q (signal_7875) ) ;
    buf_clk cell_5747 ( .C (CLK), .D (signal_7890), .Q (signal_7891) ) ;
    buf_clk cell_5763 ( .C (CLK), .D (signal_7906), .Q (signal_7907) ) ;
    buf_clk cell_5779 ( .C (CLK), .D (signal_7922), .Q (signal_7923) ) ;
    buf_clk cell_5795 ( .C (CLK), .D (signal_7938), .Q (signal_7939) ) ;
    buf_clk cell_5811 ( .C (CLK), .D (signal_7954), .Q (signal_7955) ) ;
    buf_clk cell_5827 ( .C (CLK), .D (signal_7970), .Q (signal_7971) ) ;
    buf_clk cell_5843 ( .C (CLK), .D (signal_7986), .Q (signal_7987) ) ;
    buf_clk cell_5859 ( .C (CLK), .D (signal_8002), .Q (signal_8003) ) ;
    buf_clk cell_5875 ( .C (CLK), .D (signal_8018), .Q (signal_8019) ) ;
    buf_clk cell_5891 ( .C (CLK), .D (signal_8034), .Q (signal_8035) ) ;
    buf_clk cell_5907 ( .C (CLK), .D (signal_8050), .Q (signal_8051) ) ;
    buf_clk cell_5923 ( .C (CLK), .D (signal_8066), .Q (signal_8067) ) ;
    buf_clk cell_5939 ( .C (CLK), .D (signal_8082), .Q (signal_8083) ) ;
    buf_clk cell_5955 ( .C (CLK), .D (signal_8098), .Q (signal_8099) ) ;
    buf_clk cell_5971 ( .C (CLK), .D (signal_8114), .Q (signal_8115) ) ;
    buf_clk cell_5987 ( .C (CLK), .D (signal_8130), .Q (signal_8131) ) ;
    buf_clk cell_6003 ( .C (CLK), .D (signal_8146), .Q (signal_8147) ) ;
    buf_clk cell_6019 ( .C (CLK), .D (signal_8162), .Q (signal_8163) ) ;
    buf_clk cell_6035 ( .C (CLK), .D (signal_8178), .Q (signal_8179) ) ;
    buf_clk cell_6051 ( .C (CLK), .D (signal_8194), .Q (signal_8195) ) ;
    buf_clk cell_6067 ( .C (CLK), .D (signal_8210), .Q (signal_8211) ) ;
    buf_clk cell_6083 ( .C (CLK), .D (signal_8226), .Q (signal_8227) ) ;
    buf_clk cell_6099 ( .C (CLK), .D (signal_8242), .Q (signal_8243) ) ;
    buf_clk cell_6115 ( .C (CLK), .D (signal_8258), .Q (signal_8259) ) ;
    buf_clk cell_6131 ( .C (CLK), .D (signal_8274), .Q (signal_8275) ) ;
    buf_clk cell_6147 ( .C (CLK), .D (signal_8290), .Q (signal_8291) ) ;
    buf_clk cell_6163 ( .C (CLK), .D (signal_8306), .Q (signal_8307) ) ;
    buf_clk cell_6179 ( .C (CLK), .D (signal_8322), .Q (signal_8323) ) ;
    buf_clk cell_6195 ( .C (CLK), .D (signal_8338), .Q (signal_8339) ) ;
    buf_clk cell_6211 ( .C (CLK), .D (signal_8354), .Q (signal_8355) ) ;
    buf_clk cell_6227 ( .C (CLK), .D (signal_8370), .Q (signal_8371) ) ;
    buf_clk cell_6243 ( .C (CLK), .D (signal_8386), .Q (signal_8387) ) ;
    buf_clk cell_6259 ( .C (CLK), .D (signal_8402), .Q (signal_8403) ) ;
    buf_clk cell_6275 ( .C (CLK), .D (signal_8418), .Q (signal_8419) ) ;
    buf_clk cell_6291 ( .C (CLK), .D (signal_8434), .Q (signal_8435) ) ;
    buf_clk cell_6307 ( .C (CLK), .D (signal_8450), .Q (signal_8451) ) ;
    buf_clk cell_6323 ( .C (CLK), .D (signal_8466), .Q (signal_8467) ) ;
    buf_clk cell_6339 ( .C (CLK), .D (signal_8482), .Q (signal_8483) ) ;
    buf_clk cell_6355 ( .C (CLK), .D (signal_8498), .Q (signal_8499) ) ;
    buf_clk cell_6371 ( .C (CLK), .D (signal_8514), .Q (signal_8515) ) ;
    buf_clk cell_6387 ( .C (CLK), .D (signal_8530), .Q (signal_8531) ) ;
    buf_clk cell_6403 ( .C (CLK), .D (signal_8546), .Q (signal_8547) ) ;
    buf_clk cell_6411 ( .C (CLK), .D (signal_8554), .Q (signal_8555) ) ;
    buf_clk cell_6419 ( .C (CLK), .D (signal_8562), .Q (signal_8563) ) ;
    buf_clk cell_6427 ( .C (CLK), .D (signal_8570), .Q (signal_8571) ) ;
    buf_clk cell_6435 ( .C (CLK), .D (signal_8578), .Q (signal_8579) ) ;
    buf_clk cell_6443 ( .C (CLK), .D (signal_8586), .Q (signal_8587) ) ;
    buf_clk cell_6451 ( .C (CLK), .D (signal_8594), .Q (signal_8595) ) ;
    buf_clk cell_6459 ( .C (CLK), .D (signal_8602), .Q (signal_8603) ) ;
    buf_clk cell_6467 ( .C (CLK), .D (signal_8610), .Q (signal_8611) ) ;
    buf_clk cell_6475 ( .C (CLK), .D (signal_8618), .Q (signal_8619) ) ;
    buf_clk cell_6483 ( .C (CLK), .D (signal_8626), .Q (signal_8627) ) ;
    buf_clk cell_6491 ( .C (CLK), .D (signal_8634), .Q (signal_8635) ) ;
    buf_clk cell_6499 ( .C (CLK), .D (signal_8642), .Q (signal_8643) ) ;
    buf_clk cell_6507 ( .C (CLK), .D (signal_8650), .Q (signal_8651) ) ;
    buf_clk cell_6515 ( .C (CLK), .D (signal_8658), .Q (signal_8659) ) ;
    buf_clk cell_6523 ( .C (CLK), .D (signal_8666), .Q (signal_8667) ) ;
    buf_clk cell_6531 ( .C (CLK), .D (signal_8674), .Q (signal_8675) ) ;
    buf_clk cell_6539 ( .C (CLK), .D (signal_8682), .Q (signal_8683) ) ;
    buf_clk cell_6547 ( .C (CLK), .D (signal_8690), .Q (signal_8691) ) ;
    buf_clk cell_6555 ( .C (CLK), .D (signal_8698), .Q (signal_8699) ) ;
    buf_clk cell_6563 ( .C (CLK), .D (signal_8706), .Q (signal_8707) ) ;
    buf_clk cell_6571 ( .C (CLK), .D (signal_8714), .Q (signal_8715) ) ;
    buf_clk cell_6579 ( .C (CLK), .D (signal_8722), .Q (signal_8723) ) ;
    buf_clk cell_6587 ( .C (CLK), .D (signal_8730), .Q (signal_8731) ) ;
    buf_clk cell_6595 ( .C (CLK), .D (signal_8738), .Q (signal_8739) ) ;
    buf_clk cell_6603 ( .C (CLK), .D (signal_8746), .Q (signal_8747) ) ;
    buf_clk cell_6611 ( .C (CLK), .D (signal_8754), .Q (signal_8755) ) ;
    buf_clk cell_6619 ( .C (CLK), .D (signal_8762), .Q (signal_8763) ) ;
    buf_clk cell_6627 ( .C (CLK), .D (signal_8770), .Q (signal_8771) ) ;
    buf_clk cell_6635 ( .C (CLK), .D (signal_8778), .Q (signal_8779) ) ;
    buf_clk cell_6643 ( .C (CLK), .D (signal_8786), .Q (signal_8787) ) ;
    buf_clk cell_6651 ( .C (CLK), .D (signal_8794), .Q (signal_8795) ) ;
    buf_clk cell_6659 ( .C (CLK), .D (signal_8802), .Q (signal_8803) ) ;
    buf_clk cell_6667 ( .C (CLK), .D (signal_8810), .Q (signal_8811) ) ;
    buf_clk cell_6675 ( .C (CLK), .D (signal_8818), .Q (signal_8819) ) ;
    buf_clk cell_6683 ( .C (CLK), .D (signal_8826), .Q (signal_8827) ) ;
    buf_clk cell_6691 ( .C (CLK), .D (signal_8834), .Q (signal_8835) ) ;
    buf_clk cell_6699 ( .C (CLK), .D (signal_8842), .Q (signal_8843) ) ;
    buf_clk cell_6707 ( .C (CLK), .D (signal_8850), .Q (signal_8851) ) ;
    buf_clk cell_6715 ( .C (CLK), .D (signal_8858), .Q (signal_8859) ) ;
    buf_clk cell_6723 ( .C (CLK), .D (signal_8866), .Q (signal_8867) ) ;
    buf_clk cell_6731 ( .C (CLK), .D (signal_8874), .Q (signal_8875) ) ;
    buf_clk cell_6739 ( .C (CLK), .D (signal_8882), .Q (signal_8883) ) ;
    buf_clk cell_6747 ( .C (CLK), .D (signal_8890), .Q (signal_8891) ) ;
    buf_clk cell_6755 ( .C (CLK), .D (signal_8898), .Q (signal_8899) ) ;
    buf_clk cell_6763 ( .C (CLK), .D (signal_8906), .Q (signal_8907) ) ;
    buf_clk cell_6771 ( .C (CLK), .D (signal_8914), .Q (signal_8915) ) ;
    buf_clk cell_6779 ( .C (CLK), .D (signal_8922), .Q (signal_8923) ) ;
    buf_clk cell_6787 ( .C (CLK), .D (signal_8930), .Q (signal_8931) ) ;
    buf_clk cell_6795 ( .C (CLK), .D (signal_8938), .Q (signal_8939) ) ;
    buf_clk cell_6803 ( .C (CLK), .D (signal_8946), .Q (signal_8947) ) ;
    buf_clk cell_6811 ( .C (CLK), .D (signal_8954), .Q (signal_8955) ) ;
    buf_clk cell_6819 ( .C (CLK), .D (signal_8962), .Q (signal_8963) ) ;
    buf_clk cell_6827 ( .C (CLK), .D (signal_8970), .Q (signal_8971) ) ;
    buf_clk cell_6835 ( .C (CLK), .D (signal_8978), .Q (signal_8979) ) ;
    buf_clk cell_6843 ( .C (CLK), .D (signal_8986), .Q (signal_8987) ) ;
    buf_clk cell_6851 ( .C (CLK), .D (signal_8994), .Q (signal_8995) ) ;
    buf_clk cell_6859 ( .C (CLK), .D (signal_9002), .Q (signal_9003) ) ;
    buf_clk cell_6867 ( .C (CLK), .D (signal_9010), .Q (signal_9011) ) ;
    buf_clk cell_6875 ( .C (CLK), .D (signal_9018), .Q (signal_9019) ) ;
    buf_clk cell_6883 ( .C (CLK), .D (signal_9026), .Q (signal_9027) ) ;
    buf_clk cell_6891 ( .C (CLK), .D (signal_9034), .Q (signal_9035) ) ;
    buf_clk cell_6899 ( .C (CLK), .D (signal_9042), .Q (signal_9043) ) ;
    buf_clk cell_6907 ( .C (CLK), .D (signal_9050), .Q (signal_9051) ) ;
    buf_clk cell_6915 ( .C (CLK), .D (signal_9058), .Q (signal_9059) ) ;
    buf_clk cell_6923 ( .C (CLK), .D (signal_9066), .Q (signal_9067) ) ;
    buf_clk cell_6931 ( .C (CLK), .D (signal_9074), .Q (signal_9075) ) ;
    buf_clk cell_6939 ( .C (CLK), .D (signal_9082), .Q (signal_9083) ) ;
    buf_clk cell_6947 ( .C (CLK), .D (signal_9090), .Q (signal_9091) ) ;
    buf_clk cell_6955 ( .C (CLK), .D (signal_9098), .Q (signal_9099) ) ;
    buf_clk cell_6963 ( .C (CLK), .D (signal_9106), .Q (signal_9107) ) ;
    buf_clk cell_6971 ( .C (CLK), .D (signal_9114), .Q (signal_9115) ) ;
    buf_clk cell_6979 ( .C (CLK), .D (signal_9122), .Q (signal_9123) ) ;
    buf_clk cell_6987 ( .C (CLK), .D (signal_9130), .Q (signal_9131) ) ;
    buf_clk cell_6995 ( .C (CLK), .D (signal_9138), .Q (signal_9139) ) ;
    buf_clk cell_7003 ( .C (CLK), .D (signal_9146), .Q (signal_9147) ) ;
    buf_clk cell_7011 ( .C (CLK), .D (signal_9154), .Q (signal_9155) ) ;
    buf_clk cell_7019 ( .C (CLK), .D (signal_9162), .Q (signal_9163) ) ;
    buf_clk cell_7027 ( .C (CLK), .D (signal_9170), .Q (signal_9171) ) ;
    buf_clk cell_7035 ( .C (CLK), .D (signal_9178), .Q (signal_9179) ) ;
    buf_clk cell_7043 ( .C (CLK), .D (signal_9186), .Q (signal_9187) ) ;
    buf_clk cell_7051 ( .C (CLK), .D (signal_9194), .Q (signal_9195) ) ;
    buf_clk cell_7059 ( .C (CLK), .D (signal_9202), .Q (signal_9203) ) ;
    buf_clk cell_7067 ( .C (CLK), .D (signal_9210), .Q (signal_9211) ) ;
    buf_clk cell_7075 ( .C (CLK), .D (signal_9218), .Q (signal_9219) ) ;
    buf_clk cell_7083 ( .C (CLK), .D (signal_9226), .Q (signal_9227) ) ;
    buf_clk cell_7091 ( .C (CLK), .D (signal_9234), .Q (signal_9235) ) ;
    buf_clk cell_7099 ( .C (CLK), .D (signal_9242), .Q (signal_9243) ) ;
    buf_clk cell_7107 ( .C (CLK), .D (signal_9250), .Q (signal_9251) ) ;
    buf_clk cell_7115 ( .C (CLK), .D (signal_9258), .Q (signal_9259) ) ;
    buf_clk cell_7123 ( .C (CLK), .D (signal_9266), .Q (signal_9267) ) ;
    buf_clk cell_7131 ( .C (CLK), .D (signal_9274), .Q (signal_9275) ) ;
    buf_clk cell_7139 ( .C (CLK), .D (signal_9282), .Q (signal_9283) ) ;
    buf_clk cell_7147 ( .C (CLK), .D (signal_9290), .Q (signal_9291) ) ;
    buf_clk cell_7155 ( .C (CLK), .D (signal_9298), .Q (signal_9299) ) ;
    buf_clk cell_7163 ( .C (CLK), .D (signal_9306), .Q (signal_9307) ) ;
    buf_clk cell_7171 ( .C (CLK), .D (signal_9314), .Q (signal_9315) ) ;
    buf_clk cell_7179 ( .C (CLK), .D (signal_9322), .Q (signal_9323) ) ;
    buf_clk cell_7187 ( .C (CLK), .D (signal_9330), .Q (signal_9331) ) ;
    buf_clk cell_7195 ( .C (CLK), .D (signal_9338), .Q (signal_9339) ) ;
    buf_clk cell_7203 ( .C (CLK), .D (signal_9346), .Q (signal_9347) ) ;
    buf_clk cell_7211 ( .C (CLK), .D (signal_9354), .Q (signal_9355) ) ;
    buf_clk cell_7219 ( .C (CLK), .D (signal_9362), .Q (signal_9363) ) ;
    buf_clk cell_7227 ( .C (CLK), .D (signal_9370), .Q (signal_9371) ) ;
    buf_clk cell_7235 ( .C (CLK), .D (signal_9378), .Q (signal_9379) ) ;
    buf_clk cell_7243 ( .C (CLK), .D (signal_9386), .Q (signal_9387) ) ;
    buf_clk cell_7251 ( .C (CLK), .D (signal_9394), .Q (signal_9395) ) ;
    buf_clk cell_7259 ( .C (CLK), .D (signal_9402), .Q (signal_9403) ) ;
    buf_clk cell_7267 ( .C (CLK), .D (signal_9410), .Q (signal_9411) ) ;
    buf_clk cell_7275 ( .C (CLK), .D (signal_9418), .Q (signal_9419) ) ;
    buf_clk cell_7283 ( .C (CLK), .D (signal_9426), .Q (signal_9427) ) ;
    buf_clk cell_7291 ( .C (CLK), .D (signal_9434), .Q (signal_9435) ) ;
    buf_clk cell_7299 ( .C (CLK), .D (signal_9442), .Q (signal_9443) ) ;
    buf_clk cell_7307 ( .C (CLK), .D (signal_9450), .Q (signal_9451) ) ;
    buf_clk cell_7315 ( .C (CLK), .D (signal_9458), .Q (signal_9459) ) ;
    buf_clk cell_7323 ( .C (CLK), .D (signal_9466), .Q (signal_9467) ) ;
    buf_clk cell_7331 ( .C (CLK), .D (signal_9474), .Q (signal_9475) ) ;
    buf_clk cell_7339 ( .C (CLK), .D (signal_9482), .Q (signal_9483) ) ;
    buf_clk cell_7347 ( .C (CLK), .D (signal_9490), .Q (signal_9491) ) ;
    buf_clk cell_7355 ( .C (CLK), .D (signal_9498), .Q (signal_9499) ) ;
    buf_clk cell_7363 ( .C (CLK), .D (signal_9506), .Q (signal_9507) ) ;
    buf_clk cell_7371 ( .C (CLK), .D (signal_9514), .Q (signal_9515) ) ;
    buf_clk cell_7379 ( .C (CLK), .D (signal_9522), .Q (signal_9523) ) ;
    buf_clk cell_7387 ( .C (CLK), .D (signal_9530), .Q (signal_9531) ) ;
    buf_clk cell_7395 ( .C (CLK), .D (signal_9538), .Q (signal_9539) ) ;
    buf_clk cell_7403 ( .C (CLK), .D (signal_9546), .Q (signal_9547) ) ;
    buf_clk cell_7411 ( .C (CLK), .D (signal_9554), .Q (signal_9555) ) ;
    buf_clk cell_7419 ( .C (CLK), .D (signal_9562), .Q (signal_9563) ) ;
    buf_clk cell_7427 ( .C (CLK), .D (signal_9570), .Q (signal_9571) ) ;
    buf_clk cell_7435 ( .C (CLK), .D (signal_9578), .Q (signal_9579) ) ;
    buf_clk cell_7443 ( .C (CLK), .D (signal_9586), .Q (signal_9587) ) ;
    buf_clk cell_7451 ( .C (CLK), .D (signal_9594), .Q (signal_9595) ) ;
    buf_clk cell_7459 ( .C (CLK), .D (signal_9602), .Q (signal_9603) ) ;
    buf_clk cell_7467 ( .C (CLK), .D (signal_9610), .Q (signal_9611) ) ;
    buf_clk cell_7475 ( .C (CLK), .D (signal_9618), .Q (signal_9619) ) ;
    buf_clk cell_7483 ( .C (CLK), .D (signal_9626), .Q (signal_9627) ) ;
    buf_clk cell_7491 ( .C (CLK), .D (signal_9634), .Q (signal_9635) ) ;
    buf_clk cell_7499 ( .C (CLK), .D (signal_9642), .Q (signal_9643) ) ;
    buf_clk cell_7507 ( .C (CLK), .D (signal_9650), .Q (signal_9651) ) ;
    buf_clk cell_7515 ( .C (CLK), .D (signal_9658), .Q (signal_9659) ) ;
    buf_clk cell_7523 ( .C (CLK), .D (signal_9666), .Q (signal_9667) ) ;
    buf_clk cell_7531 ( .C (CLK), .D (signal_9674), .Q (signal_9675) ) ;
    buf_clk cell_7539 ( .C (CLK), .D (signal_9682), .Q (signal_9683) ) ;
    buf_clk cell_7547 ( .C (CLK), .D (signal_9690), .Q (signal_9691) ) ;
    buf_clk cell_7555 ( .C (CLK), .D (signal_9698), .Q (signal_9699) ) ;
    buf_clk cell_7559 ( .C (CLK), .D (signal_9702), .Q (signal_9703) ) ;
    buf_clk cell_7561 ( .C (CLK), .D (signal_9704), .Q (signal_9705) ) ;
    buf_clk cell_7569 ( .C (CLK), .D (signal_9712), .Q (signal_9713) ) ;
    buf_clk cell_7577 ( .C (CLK), .D (signal_9720), .Q (signal_9721) ) ;
    buf_clk cell_7581 ( .C (CLK), .D (signal_9724), .Q (signal_9725) ) ;
    buf_clk cell_7585 ( .C (CLK), .D (signal_9728), .Q (signal_9729) ) ;
    buf_clk cell_7587 ( .C (CLK), .D (signal_9730), .Q (signal_9731) ) ;
    buf_clk cell_7589 ( .C (CLK), .D (signal_9732), .Q (signal_9733) ) ;
    buf_clk cell_7603 ( .C (CLK), .D (signal_9746), .Q (signal_9747) ) ;
    buf_clk cell_7619 ( .C (CLK), .D (signal_9762), .Q (signal_9763) ) ;
    buf_clk cell_7635 ( .C (CLK), .D (signal_9778), .Q (signal_9779) ) ;
    buf_clk cell_7651 ( .C (CLK), .D (signal_9794), .Q (signal_9795) ) ;
    buf_clk cell_7667 ( .C (CLK), .D (signal_9810), .Q (signal_9811) ) ;
    buf_clk cell_7683 ( .C (CLK), .D (signal_9826), .Q (signal_9827) ) ;
    buf_clk cell_7699 ( .C (CLK), .D (signal_9842), .Q (signal_9843) ) ;
    buf_clk cell_7715 ( .C (CLK), .D (signal_9858), .Q (signal_9859) ) ;
    buf_clk cell_7731 ( .C (CLK), .D (signal_9874), .Q (signal_9875) ) ;
    buf_clk cell_7747 ( .C (CLK), .D (signal_9890), .Q (signal_9891) ) ;
    buf_clk cell_7755 ( .C (CLK), .D (signal_9898), .Q (signal_9899) ) ;
    buf_clk cell_7763 ( .C (CLK), .D (signal_9906), .Q (signal_9907) ) ;
    buf_clk cell_7771 ( .C (CLK), .D (signal_9914), .Q (signal_9915) ) ;
    buf_clk cell_7779 ( .C (CLK), .D (signal_9922), .Q (signal_9923) ) ;
    buf_clk cell_7787 ( .C (CLK), .D (signal_9930), .Q (signal_9931) ) ;
    buf_clk cell_7795 ( .C (CLK), .D (signal_9938), .Q (signal_9939) ) ;
    buf_clk cell_7803 ( .C (CLK), .D (signal_9946), .Q (signal_9947) ) ;
    buf_clk cell_7811 ( .C (CLK), .D (signal_9954), .Q (signal_9955) ) ;
    buf_clk cell_7819 ( .C (CLK), .D (signal_9962), .Q (signal_9963) ) ;
    buf_clk cell_7827 ( .C (CLK), .D (signal_9970), .Q (signal_9971) ) ;
    buf_clk cell_7835 ( .C (CLK), .D (signal_9978), .Q (signal_9979) ) ;
    buf_clk cell_7843 ( .C (CLK), .D (signal_9986), .Q (signal_9987) ) ;
    buf_clk cell_7851 ( .C (CLK), .D (signal_9994), .Q (signal_9995) ) ;
    buf_clk cell_7859 ( .C (CLK), .D (signal_10002), .Q (signal_10003) ) ;
    buf_clk cell_7867 ( .C (CLK), .D (signal_10010), .Q (signal_10011) ) ;
    buf_clk cell_7875 ( .C (CLK), .D (signal_10018), .Q (signal_10019) ) ;
    buf_clk cell_7883 ( .C (CLK), .D (signal_10026), .Q (signal_10027) ) ;
    buf_clk cell_7891 ( .C (CLK), .D (signal_10034), .Q (signal_10035) ) ;
    buf_clk cell_7899 ( .C (CLK), .D (signal_10042), .Q (signal_10043) ) ;
    buf_clk cell_7907 ( .C (CLK), .D (signal_10050), .Q (signal_10051) ) ;
    buf_clk cell_7915 ( .C (CLK), .D (signal_10058), .Q (signal_10059) ) ;
    buf_clk cell_7923 ( .C (CLK), .D (signal_10066), .Q (signal_10067) ) ;
    buf_clk cell_7931 ( .C (CLK), .D (signal_10074), .Q (signal_10075) ) ;
    buf_clk cell_7939 ( .C (CLK), .D (signal_10082), .Q (signal_10083) ) ;
    buf_clk cell_7955 ( .C (CLK), .D (signal_10098), .Q (signal_10099) ) ;

    /* cells in depth 15 */
    buf_clk cell_3444 ( .C (CLK), .D (signal_5587), .Q (signal_5588) ) ;
    buf_clk cell_3460 ( .C (CLK), .D (signal_5603), .Q (signal_5604) ) ;
    buf_clk cell_3476 ( .C (CLK), .D (signal_5619), .Q (signal_5620) ) ;
    buf_clk cell_3484 ( .C (CLK), .D (signal_5627), .Q (signal_5628) ) ;
    buf_clk cell_3500 ( .C (CLK), .D (signal_5643), .Q (signal_5644) ) ;
    buf_clk cell_3516 ( .C (CLK), .D (signal_5659), .Q (signal_5660) ) ;
    buf_clk cell_3524 ( .C (CLK), .D (signal_5667), .Q (signal_5668) ) ;
    buf_clk cell_3540 ( .C (CLK), .D (signal_5683), .Q (signal_5684) ) ;
    buf_clk cell_3556 ( .C (CLK), .D (signal_5699), .Q (signal_5700) ) ;
    buf_clk cell_3572 ( .C (CLK), .D (signal_5715), .Q (signal_5716) ) ;
    buf_clk cell_3588 ( .C (CLK), .D (signal_5731), .Q (signal_5732) ) ;
    buf_clk cell_3592 ( .C (CLK), .D (signal_5735), .Q (signal_5736) ) ;
    buf_clk cell_3596 ( .C (CLK), .D (signal_5739), .Q (signal_5740) ) ;
    buf_clk cell_3602 ( .C (CLK), .D (signal_5745), .Q (signal_5746) ) ;
    buf_clk cell_3608 ( .C (CLK), .D (signal_5751), .Q (signal_5752) ) ;
    buf_clk cell_3614 ( .C (CLK), .D (signal_5757), .Q (signal_5758) ) ;
    buf_clk cell_3620 ( .C (CLK), .D (signal_5763), .Q (signal_5764) ) ;
    buf_clk cell_3626 ( .C (CLK), .D (signal_5769), .Q (signal_5770) ) ;
    buf_clk cell_3632 ( .C (CLK), .D (signal_5775), .Q (signal_5776) ) ;
    buf_clk cell_3648 ( .C (CLK), .D (signal_5791), .Q (signal_5792) ) ;
    buf_clk cell_3664 ( .C (CLK), .D (signal_5807), .Q (signal_5808) ) ;
    buf_clk cell_3680 ( .C (CLK), .D (signal_5823), .Q (signal_5824) ) ;
    buf_clk cell_3696 ( .C (CLK), .D (signal_5839), .Q (signal_5840) ) ;
    buf_clk cell_3712 ( .C (CLK), .D (signal_5855), .Q (signal_5856) ) ;
    buf_clk cell_3728 ( .C (CLK), .D (signal_5871), .Q (signal_5872) ) ;
    buf_clk cell_3744 ( .C (CLK), .D (signal_5887), .Q (signal_5888) ) ;
    buf_clk cell_3760 ( .C (CLK), .D (signal_5903), .Q (signal_5904) ) ;
    buf_clk cell_3776 ( .C (CLK), .D (signal_5919), .Q (signal_5920) ) ;
    buf_clk cell_3792 ( .C (CLK), .D (signal_5935), .Q (signal_5936) ) ;
    buf_clk cell_3796 ( .C (CLK), .D (signal_5939), .Q (signal_5940) ) ;
    buf_clk cell_3800 ( .C (CLK), .D (signal_5943), .Q (signal_5944) ) ;
    buf_clk cell_3808 ( .C (CLK), .D (signal_5951), .Q (signal_5952) ) ;
    buf_clk cell_3816 ( .C (CLK), .D (signal_5959), .Q (signal_5960) ) ;
    buf_clk cell_3822 ( .C (CLK), .D (signal_5965), .Q (signal_5966) ) ;
    buf_clk cell_3828 ( .C (CLK), .D (signal_5971), .Q (signal_5972) ) ;
    buf_clk cell_3836 ( .C (CLK), .D (signal_5979), .Q (signal_5980) ) ;
    buf_clk cell_3844 ( .C (CLK), .D (signal_5987), .Q (signal_5988) ) ;
    buf_clk cell_3852 ( .C (CLK), .D (signal_5995), .Q (signal_5996) ) ;
    buf_clk cell_3860 ( .C (CLK), .D (signal_6003), .Q (signal_6004) ) ;
    buf_clk cell_3864 ( .C (CLK), .D (signal_6007), .Q (signal_6008) ) ;
    buf_clk cell_3868 ( .C (CLK), .D (signal_6011), .Q (signal_6012) ) ;
    buf_clk cell_3876 ( .C (CLK), .D (signal_6019), .Q (signal_6020) ) ;
    buf_clk cell_3884 ( .C (CLK), .D (signal_6027), .Q (signal_6028) ) ;
    buf_clk cell_3900 ( .C (CLK), .D (signal_6043), .Q (signal_6044) ) ;
    buf_clk cell_3916 ( .C (CLK), .D (signal_6059), .Q (signal_6060) ) ;
    buf_clk cell_3932 ( .C (CLK), .D (signal_6075), .Q (signal_6076) ) ;
    buf_clk cell_3948 ( .C (CLK), .D (signal_6091), .Q (signal_6092) ) ;
    buf_clk cell_3964 ( .C (CLK), .D (signal_6107), .Q (signal_6108) ) ;
    buf_clk cell_3980 ( .C (CLK), .D (signal_6123), .Q (signal_6124) ) ;
    buf_clk cell_3996 ( .C (CLK), .D (signal_6139), .Q (signal_6140) ) ;
    buf_clk cell_4012 ( .C (CLK), .D (signal_6155), .Q (signal_6156) ) ;
    buf_clk cell_4028 ( .C (CLK), .D (signal_6171), .Q (signal_6172) ) ;
    buf_clk cell_4044 ( .C (CLK), .D (signal_6187), .Q (signal_6188) ) ;
    buf_clk cell_4060 ( .C (CLK), .D (signal_6203), .Q (signal_6204) ) ;
    buf_clk cell_4076 ( .C (CLK), .D (signal_6219), .Q (signal_6220) ) ;
    buf_clk cell_4092 ( .C (CLK), .D (signal_6235), .Q (signal_6236) ) ;
    buf_clk cell_4108 ( .C (CLK), .D (signal_6251), .Q (signal_6252) ) ;
    buf_clk cell_4118 ( .C (CLK), .D (signal_6261), .Q (signal_6262) ) ;
    buf_clk cell_4128 ( .C (CLK), .D (signal_6271), .Q (signal_6272) ) ;
    buf_clk cell_4134 ( .C (CLK), .D (signal_6277), .Q (signal_6278) ) ;
    buf_clk cell_4140 ( .C (CLK), .D (signal_6283), .Q (signal_6284) ) ;
    buf_clk cell_4148 ( .C (CLK), .D (signal_6291), .Q (signal_6292) ) ;
    buf_clk cell_4156 ( .C (CLK), .D (signal_6299), .Q (signal_6300) ) ;
    buf_clk cell_4166 ( .C (CLK), .D (signal_6309), .Q (signal_6310) ) ;
    buf_clk cell_4176 ( .C (CLK), .D (signal_6319), .Q (signal_6320) ) ;
    buf_clk cell_4192 ( .C (CLK), .D (signal_6335), .Q (signal_6336) ) ;
    buf_clk cell_4204 ( .C (CLK), .D (signal_6347), .Q (signal_6348) ) ;
    buf_clk cell_4216 ( .C (CLK), .D (signal_6359), .Q (signal_6360) ) ;
    buf_clk cell_4224 ( .C (CLK), .D (signal_6367), .Q (signal_6368) ) ;
    buf_clk cell_4232 ( .C (CLK), .D (signal_6375), .Q (signal_6376) ) ;
    buf_clk cell_4244 ( .C (CLK), .D (signal_6387), .Q (signal_6388) ) ;
    buf_clk cell_4256 ( .C (CLK), .D (signal_6399), .Q (signal_6400) ) ;
    buf_clk cell_4270 ( .C (CLK), .D (signal_6413), .Q (signal_6414) ) ;
    buf_clk cell_4284 ( .C (CLK), .D (signal_6427), .Q (signal_6428) ) ;
    buf_clk cell_4300 ( .C (CLK), .D (signal_6443), .Q (signal_6444) ) ;
    buf_clk cell_4316 ( .C (CLK), .D (signal_6459), .Q (signal_6460) ) ;
    buf_clk cell_4332 ( .C (CLK), .D (signal_6475), .Q (signal_6476) ) ;
    buf_clk cell_4348 ( .C (CLK), .D (signal_6491), .Q (signal_6492) ) ;
    buf_clk cell_4364 ( .C (CLK), .D (signal_6507), .Q (signal_6508) ) ;
    buf_clk cell_4380 ( .C (CLK), .D (signal_6523), .Q (signal_6524) ) ;
    buf_clk cell_4396 ( .C (CLK), .D (signal_6539), .Q (signal_6540) ) ;
    buf_clk cell_4412 ( .C (CLK), .D (signal_6555), .Q (signal_6556) ) ;
    buf_clk cell_4428 ( .C (CLK), .D (signal_6571), .Q (signal_6572) ) ;
    buf_clk cell_4444 ( .C (CLK), .D (signal_6587), .Q (signal_6588) ) ;
    buf_clk cell_4460 ( .C (CLK), .D (signal_6603), .Q (signal_6604) ) ;
    buf_clk cell_4476 ( .C (CLK), .D (signal_6619), .Q (signal_6620) ) ;
    buf_clk cell_4492 ( .C (CLK), .D (signal_6635), .Q (signal_6636) ) ;
    buf_clk cell_4508 ( .C (CLK), .D (signal_6651), .Q (signal_6652) ) ;
    buf_clk cell_4524 ( .C (CLK), .D (signal_6667), .Q (signal_6668) ) ;
    buf_clk cell_4540 ( .C (CLK), .D (signal_6683), .Q (signal_6684) ) ;
    buf_clk cell_4550 ( .C (CLK), .D (signal_6693), .Q (signal_6694) ) ;
    buf_clk cell_4560 ( .C (CLK), .D (signal_6703), .Q (signal_6704) ) ;
    buf_clk cell_4568 ( .C (CLK), .D (signal_6711), .Q (signal_6712) ) ;
    buf_clk cell_4576 ( .C (CLK), .D (signal_6719), .Q (signal_6720) ) ;
    buf_clk cell_4588 ( .C (CLK), .D (signal_6731), .Q (signal_6732) ) ;
    buf_clk cell_4600 ( .C (CLK), .D (signal_6743), .Q (signal_6744) ) ;
    buf_clk cell_4614 ( .C (CLK), .D (signal_6757), .Q (signal_6758) ) ;
    buf_clk cell_4628 ( .C (CLK), .D (signal_6771), .Q (signal_6772) ) ;
    buf_clk cell_4644 ( .C (CLK), .D (signal_6787), .Q (signal_6788) ) ;
    buf_clk cell_4660 ( .C (CLK), .D (signal_6803), .Q (signal_6804) ) ;
    buf_clk cell_4666 ( .C (CLK), .D (signal_6809), .Q (signal_6810) ) ;
    buf_clk cell_4672 ( .C (CLK), .D (signal_6815), .Q (signal_6816) ) ;
    buf_clk cell_4680 ( .C (CLK), .D (signal_6823), .Q (signal_6824) ) ;
    buf_clk cell_4688 ( .C (CLK), .D (signal_6831), .Q (signal_6832) ) ;
    buf_clk cell_4698 ( .C (CLK), .D (signal_6841), .Q (signal_6842) ) ;
    buf_clk cell_4708 ( .C (CLK), .D (signal_6851), .Q (signal_6852) ) ;
    buf_clk cell_4720 ( .C (CLK), .D (signal_6863), .Q (signal_6864) ) ;
    buf_clk cell_4732 ( .C (CLK), .D (signal_6875), .Q (signal_6876) ) ;
    buf_clk cell_4740 ( .C (CLK), .D (signal_6883), .Q (signal_6884) ) ;
    buf_clk cell_4756 ( .C (CLK), .D (signal_6899), .Q (signal_6900) ) ;
    buf_clk cell_4772 ( .C (CLK), .D (signal_6915), .Q (signal_6916) ) ;
    buf_clk cell_4788 ( .C (CLK), .D (signal_6931), .Q (signal_6932) ) ;
    buf_clk cell_4804 ( .C (CLK), .D (signal_6947), .Q (signal_6948) ) ;
    buf_clk cell_4820 ( .C (CLK), .D (signal_6963), .Q (signal_6964) ) ;
    buf_clk cell_4836 ( .C (CLK), .D (signal_6979), .Q (signal_6980) ) ;
    buf_clk cell_4852 ( .C (CLK), .D (signal_6995), .Q (signal_6996) ) ;
    buf_clk cell_4868 ( .C (CLK), .D (signal_7011), .Q (signal_7012) ) ;
    buf_clk cell_4884 ( .C (CLK), .D (signal_7027), .Q (signal_7028) ) ;
    buf_clk cell_4900 ( .C (CLK), .D (signal_7043), .Q (signal_7044) ) ;
    buf_clk cell_4916 ( .C (CLK), .D (signal_7059), .Q (signal_7060) ) ;
    buf_clk cell_4932 ( .C (CLK), .D (signal_7075), .Q (signal_7076) ) ;
    buf_clk cell_4948 ( .C (CLK), .D (signal_7091), .Q (signal_7092) ) ;
    buf_clk cell_4964 ( .C (CLK), .D (signal_7107), .Q (signal_7108) ) ;
    buf_clk cell_4980 ( .C (CLK), .D (signal_7123), .Q (signal_7124) ) ;
    buf_clk cell_4996 ( .C (CLK), .D (signal_7139), .Q (signal_7140) ) ;
    buf_clk cell_5012 ( .C (CLK), .D (signal_7155), .Q (signal_7156) ) ;
    buf_clk cell_5028 ( .C (CLK), .D (signal_7171), .Q (signal_7172) ) ;
    buf_clk cell_5044 ( .C (CLK), .D (signal_7187), .Q (signal_7188) ) ;
    buf_clk cell_5060 ( .C (CLK), .D (signal_7203), .Q (signal_7204) ) ;
    buf_clk cell_5076 ( .C (CLK), .D (signal_7219), .Q (signal_7220) ) ;
    buf_clk cell_5092 ( .C (CLK), .D (signal_7235), .Q (signal_7236) ) ;
    buf_clk cell_5108 ( .C (CLK), .D (signal_7251), .Q (signal_7252) ) ;
    buf_clk cell_5124 ( .C (CLK), .D (signal_7267), .Q (signal_7268) ) ;
    buf_clk cell_5140 ( .C (CLK), .D (signal_7283), .Q (signal_7284) ) ;
    buf_clk cell_5156 ( .C (CLK), .D (signal_7299), .Q (signal_7300) ) ;
    buf_clk cell_5172 ( .C (CLK), .D (signal_7315), .Q (signal_7316) ) ;
    buf_clk cell_5188 ( .C (CLK), .D (signal_7331), .Q (signal_7332) ) ;
    buf_clk cell_5204 ( .C (CLK), .D (signal_7347), .Q (signal_7348) ) ;
    buf_clk cell_5220 ( .C (CLK), .D (signal_7363), .Q (signal_7364) ) ;
    buf_clk cell_5236 ( .C (CLK), .D (signal_7379), .Q (signal_7380) ) ;
    buf_clk cell_5252 ( .C (CLK), .D (signal_7395), .Q (signal_7396) ) ;
    buf_clk cell_5268 ( .C (CLK), .D (signal_7411), .Q (signal_7412) ) ;
    buf_clk cell_5284 ( .C (CLK), .D (signal_7427), .Q (signal_7428) ) ;
    buf_clk cell_5300 ( .C (CLK), .D (signal_7443), .Q (signal_7444) ) ;
    buf_clk cell_5316 ( .C (CLK), .D (signal_7459), .Q (signal_7460) ) ;
    buf_clk cell_5332 ( .C (CLK), .D (signal_7475), .Q (signal_7476) ) ;
    buf_clk cell_5348 ( .C (CLK), .D (signal_7491), .Q (signal_7492) ) ;
    buf_clk cell_5364 ( .C (CLK), .D (signal_7507), .Q (signal_7508) ) ;
    buf_clk cell_5380 ( .C (CLK), .D (signal_7523), .Q (signal_7524) ) ;
    buf_clk cell_5396 ( .C (CLK), .D (signal_7539), .Q (signal_7540) ) ;
    buf_clk cell_5412 ( .C (CLK), .D (signal_7555), .Q (signal_7556) ) ;
    buf_clk cell_5428 ( .C (CLK), .D (signal_7571), .Q (signal_7572) ) ;
    buf_clk cell_5444 ( .C (CLK), .D (signal_7587), .Q (signal_7588) ) ;
    buf_clk cell_5460 ( .C (CLK), .D (signal_7603), .Q (signal_7604) ) ;
    buf_clk cell_5476 ( .C (CLK), .D (signal_7619), .Q (signal_7620) ) ;
    buf_clk cell_5492 ( .C (CLK), .D (signal_7635), .Q (signal_7636) ) ;
    buf_clk cell_5508 ( .C (CLK), .D (signal_7651), .Q (signal_7652) ) ;
    buf_clk cell_5524 ( .C (CLK), .D (signal_7667), .Q (signal_7668) ) ;
    buf_clk cell_5540 ( .C (CLK), .D (signal_7683), .Q (signal_7684) ) ;
    buf_clk cell_5556 ( .C (CLK), .D (signal_7699), .Q (signal_7700) ) ;
    buf_clk cell_5572 ( .C (CLK), .D (signal_7715), .Q (signal_7716) ) ;
    buf_clk cell_5588 ( .C (CLK), .D (signal_7731), .Q (signal_7732) ) ;
    buf_clk cell_5604 ( .C (CLK), .D (signal_7747), .Q (signal_7748) ) ;
    buf_clk cell_5620 ( .C (CLK), .D (signal_7763), .Q (signal_7764) ) ;
    buf_clk cell_5636 ( .C (CLK), .D (signal_7779), .Q (signal_7780) ) ;
    buf_clk cell_5652 ( .C (CLK), .D (signal_7795), .Q (signal_7796) ) ;
    buf_clk cell_5668 ( .C (CLK), .D (signal_7811), .Q (signal_7812) ) ;
    buf_clk cell_5684 ( .C (CLK), .D (signal_7827), .Q (signal_7828) ) ;
    buf_clk cell_5700 ( .C (CLK), .D (signal_7843), .Q (signal_7844) ) ;
    buf_clk cell_5716 ( .C (CLK), .D (signal_7859), .Q (signal_7860) ) ;
    buf_clk cell_5732 ( .C (CLK), .D (signal_7875), .Q (signal_7876) ) ;
    buf_clk cell_5748 ( .C (CLK), .D (signal_7891), .Q (signal_7892) ) ;
    buf_clk cell_5764 ( .C (CLK), .D (signal_7907), .Q (signal_7908) ) ;
    buf_clk cell_5780 ( .C (CLK), .D (signal_7923), .Q (signal_7924) ) ;
    buf_clk cell_5796 ( .C (CLK), .D (signal_7939), .Q (signal_7940) ) ;
    buf_clk cell_5812 ( .C (CLK), .D (signal_7955), .Q (signal_7956) ) ;
    buf_clk cell_5828 ( .C (CLK), .D (signal_7971), .Q (signal_7972) ) ;
    buf_clk cell_5844 ( .C (CLK), .D (signal_7987), .Q (signal_7988) ) ;
    buf_clk cell_5860 ( .C (CLK), .D (signal_8003), .Q (signal_8004) ) ;
    buf_clk cell_5876 ( .C (CLK), .D (signal_8019), .Q (signal_8020) ) ;
    buf_clk cell_5892 ( .C (CLK), .D (signal_8035), .Q (signal_8036) ) ;
    buf_clk cell_5908 ( .C (CLK), .D (signal_8051), .Q (signal_8052) ) ;
    buf_clk cell_5924 ( .C (CLK), .D (signal_8067), .Q (signal_8068) ) ;
    buf_clk cell_5940 ( .C (CLK), .D (signal_8083), .Q (signal_8084) ) ;
    buf_clk cell_5956 ( .C (CLK), .D (signal_8099), .Q (signal_8100) ) ;
    buf_clk cell_5972 ( .C (CLK), .D (signal_8115), .Q (signal_8116) ) ;
    buf_clk cell_5988 ( .C (CLK), .D (signal_8131), .Q (signal_8132) ) ;
    buf_clk cell_6004 ( .C (CLK), .D (signal_8147), .Q (signal_8148) ) ;
    buf_clk cell_6020 ( .C (CLK), .D (signal_8163), .Q (signal_8164) ) ;
    buf_clk cell_6036 ( .C (CLK), .D (signal_8179), .Q (signal_8180) ) ;
    buf_clk cell_6052 ( .C (CLK), .D (signal_8195), .Q (signal_8196) ) ;
    buf_clk cell_6068 ( .C (CLK), .D (signal_8211), .Q (signal_8212) ) ;
    buf_clk cell_6084 ( .C (CLK), .D (signal_8227), .Q (signal_8228) ) ;
    buf_clk cell_6100 ( .C (CLK), .D (signal_8243), .Q (signal_8244) ) ;
    buf_clk cell_6116 ( .C (CLK), .D (signal_8259), .Q (signal_8260) ) ;
    buf_clk cell_6132 ( .C (CLK), .D (signal_8275), .Q (signal_8276) ) ;
    buf_clk cell_6148 ( .C (CLK), .D (signal_8291), .Q (signal_8292) ) ;
    buf_clk cell_6164 ( .C (CLK), .D (signal_8307), .Q (signal_8308) ) ;
    buf_clk cell_6180 ( .C (CLK), .D (signal_8323), .Q (signal_8324) ) ;
    buf_clk cell_6196 ( .C (CLK), .D (signal_8339), .Q (signal_8340) ) ;
    buf_clk cell_6212 ( .C (CLK), .D (signal_8355), .Q (signal_8356) ) ;
    buf_clk cell_6228 ( .C (CLK), .D (signal_8371), .Q (signal_8372) ) ;
    buf_clk cell_6244 ( .C (CLK), .D (signal_8387), .Q (signal_8388) ) ;
    buf_clk cell_6260 ( .C (CLK), .D (signal_8403), .Q (signal_8404) ) ;
    buf_clk cell_6276 ( .C (CLK), .D (signal_8419), .Q (signal_8420) ) ;
    buf_clk cell_6292 ( .C (CLK), .D (signal_8435), .Q (signal_8436) ) ;
    buf_clk cell_6308 ( .C (CLK), .D (signal_8451), .Q (signal_8452) ) ;
    buf_clk cell_6324 ( .C (CLK), .D (signal_8467), .Q (signal_8468) ) ;
    buf_clk cell_6340 ( .C (CLK), .D (signal_8483), .Q (signal_8484) ) ;
    buf_clk cell_6356 ( .C (CLK), .D (signal_8499), .Q (signal_8500) ) ;
    buf_clk cell_6372 ( .C (CLK), .D (signal_8515), .Q (signal_8516) ) ;
    buf_clk cell_6388 ( .C (CLK), .D (signal_8531), .Q (signal_8532) ) ;
    buf_clk cell_6404 ( .C (CLK), .D (signal_8547), .Q (signal_8548) ) ;
    buf_clk cell_6412 ( .C (CLK), .D (signal_8555), .Q (signal_8556) ) ;
    buf_clk cell_6420 ( .C (CLK), .D (signal_8563), .Q (signal_8564) ) ;
    buf_clk cell_6428 ( .C (CLK), .D (signal_8571), .Q (signal_8572) ) ;
    buf_clk cell_6436 ( .C (CLK), .D (signal_8579), .Q (signal_8580) ) ;
    buf_clk cell_6444 ( .C (CLK), .D (signal_8587), .Q (signal_8588) ) ;
    buf_clk cell_6452 ( .C (CLK), .D (signal_8595), .Q (signal_8596) ) ;
    buf_clk cell_6460 ( .C (CLK), .D (signal_8603), .Q (signal_8604) ) ;
    buf_clk cell_6468 ( .C (CLK), .D (signal_8611), .Q (signal_8612) ) ;
    buf_clk cell_6476 ( .C (CLK), .D (signal_8619), .Q (signal_8620) ) ;
    buf_clk cell_6484 ( .C (CLK), .D (signal_8627), .Q (signal_8628) ) ;
    buf_clk cell_6492 ( .C (CLK), .D (signal_8635), .Q (signal_8636) ) ;
    buf_clk cell_6500 ( .C (CLK), .D (signal_8643), .Q (signal_8644) ) ;
    buf_clk cell_6508 ( .C (CLK), .D (signal_8651), .Q (signal_8652) ) ;
    buf_clk cell_6516 ( .C (CLK), .D (signal_8659), .Q (signal_8660) ) ;
    buf_clk cell_6524 ( .C (CLK), .D (signal_8667), .Q (signal_8668) ) ;
    buf_clk cell_6532 ( .C (CLK), .D (signal_8675), .Q (signal_8676) ) ;
    buf_clk cell_6540 ( .C (CLK), .D (signal_8683), .Q (signal_8684) ) ;
    buf_clk cell_6548 ( .C (CLK), .D (signal_8691), .Q (signal_8692) ) ;
    buf_clk cell_6556 ( .C (CLK), .D (signal_8699), .Q (signal_8700) ) ;
    buf_clk cell_6564 ( .C (CLK), .D (signal_8707), .Q (signal_8708) ) ;
    buf_clk cell_6572 ( .C (CLK), .D (signal_8715), .Q (signal_8716) ) ;
    buf_clk cell_6580 ( .C (CLK), .D (signal_8723), .Q (signal_8724) ) ;
    buf_clk cell_6588 ( .C (CLK), .D (signal_8731), .Q (signal_8732) ) ;
    buf_clk cell_6596 ( .C (CLK), .D (signal_8739), .Q (signal_8740) ) ;
    buf_clk cell_6604 ( .C (CLK), .D (signal_8747), .Q (signal_8748) ) ;
    buf_clk cell_6612 ( .C (CLK), .D (signal_8755), .Q (signal_8756) ) ;
    buf_clk cell_6620 ( .C (CLK), .D (signal_8763), .Q (signal_8764) ) ;
    buf_clk cell_6628 ( .C (CLK), .D (signal_8771), .Q (signal_8772) ) ;
    buf_clk cell_6636 ( .C (CLK), .D (signal_8779), .Q (signal_8780) ) ;
    buf_clk cell_6644 ( .C (CLK), .D (signal_8787), .Q (signal_8788) ) ;
    buf_clk cell_6652 ( .C (CLK), .D (signal_8795), .Q (signal_8796) ) ;
    buf_clk cell_6660 ( .C (CLK), .D (signal_8803), .Q (signal_8804) ) ;
    buf_clk cell_6668 ( .C (CLK), .D (signal_8811), .Q (signal_8812) ) ;
    buf_clk cell_6676 ( .C (CLK), .D (signal_8819), .Q (signal_8820) ) ;
    buf_clk cell_6684 ( .C (CLK), .D (signal_8827), .Q (signal_8828) ) ;
    buf_clk cell_6692 ( .C (CLK), .D (signal_8835), .Q (signal_8836) ) ;
    buf_clk cell_6700 ( .C (CLK), .D (signal_8843), .Q (signal_8844) ) ;
    buf_clk cell_6708 ( .C (CLK), .D (signal_8851), .Q (signal_8852) ) ;
    buf_clk cell_6716 ( .C (CLK), .D (signal_8859), .Q (signal_8860) ) ;
    buf_clk cell_6724 ( .C (CLK), .D (signal_8867), .Q (signal_8868) ) ;
    buf_clk cell_6732 ( .C (CLK), .D (signal_8875), .Q (signal_8876) ) ;
    buf_clk cell_6740 ( .C (CLK), .D (signal_8883), .Q (signal_8884) ) ;
    buf_clk cell_6748 ( .C (CLK), .D (signal_8891), .Q (signal_8892) ) ;
    buf_clk cell_6756 ( .C (CLK), .D (signal_8899), .Q (signal_8900) ) ;
    buf_clk cell_6764 ( .C (CLK), .D (signal_8907), .Q (signal_8908) ) ;
    buf_clk cell_6772 ( .C (CLK), .D (signal_8915), .Q (signal_8916) ) ;
    buf_clk cell_6780 ( .C (CLK), .D (signal_8923), .Q (signal_8924) ) ;
    buf_clk cell_6788 ( .C (CLK), .D (signal_8931), .Q (signal_8932) ) ;
    buf_clk cell_6796 ( .C (CLK), .D (signal_8939), .Q (signal_8940) ) ;
    buf_clk cell_6804 ( .C (CLK), .D (signal_8947), .Q (signal_8948) ) ;
    buf_clk cell_6812 ( .C (CLK), .D (signal_8955), .Q (signal_8956) ) ;
    buf_clk cell_6820 ( .C (CLK), .D (signal_8963), .Q (signal_8964) ) ;
    buf_clk cell_6828 ( .C (CLK), .D (signal_8971), .Q (signal_8972) ) ;
    buf_clk cell_6836 ( .C (CLK), .D (signal_8979), .Q (signal_8980) ) ;
    buf_clk cell_6844 ( .C (CLK), .D (signal_8987), .Q (signal_8988) ) ;
    buf_clk cell_6852 ( .C (CLK), .D (signal_8995), .Q (signal_8996) ) ;
    buf_clk cell_6860 ( .C (CLK), .D (signal_9003), .Q (signal_9004) ) ;
    buf_clk cell_6868 ( .C (CLK), .D (signal_9011), .Q (signal_9012) ) ;
    buf_clk cell_6876 ( .C (CLK), .D (signal_9019), .Q (signal_9020) ) ;
    buf_clk cell_6884 ( .C (CLK), .D (signal_9027), .Q (signal_9028) ) ;
    buf_clk cell_6892 ( .C (CLK), .D (signal_9035), .Q (signal_9036) ) ;
    buf_clk cell_6900 ( .C (CLK), .D (signal_9043), .Q (signal_9044) ) ;
    buf_clk cell_6908 ( .C (CLK), .D (signal_9051), .Q (signal_9052) ) ;
    buf_clk cell_6916 ( .C (CLK), .D (signal_9059), .Q (signal_9060) ) ;
    buf_clk cell_6924 ( .C (CLK), .D (signal_9067), .Q (signal_9068) ) ;
    buf_clk cell_6932 ( .C (CLK), .D (signal_9075), .Q (signal_9076) ) ;
    buf_clk cell_6940 ( .C (CLK), .D (signal_9083), .Q (signal_9084) ) ;
    buf_clk cell_6948 ( .C (CLK), .D (signal_9091), .Q (signal_9092) ) ;
    buf_clk cell_6956 ( .C (CLK), .D (signal_9099), .Q (signal_9100) ) ;
    buf_clk cell_6964 ( .C (CLK), .D (signal_9107), .Q (signal_9108) ) ;
    buf_clk cell_6972 ( .C (CLK), .D (signal_9115), .Q (signal_9116) ) ;
    buf_clk cell_6980 ( .C (CLK), .D (signal_9123), .Q (signal_9124) ) ;
    buf_clk cell_6988 ( .C (CLK), .D (signal_9131), .Q (signal_9132) ) ;
    buf_clk cell_6996 ( .C (CLK), .D (signal_9139), .Q (signal_9140) ) ;
    buf_clk cell_7004 ( .C (CLK), .D (signal_9147), .Q (signal_9148) ) ;
    buf_clk cell_7012 ( .C (CLK), .D (signal_9155), .Q (signal_9156) ) ;
    buf_clk cell_7020 ( .C (CLK), .D (signal_9163), .Q (signal_9164) ) ;
    buf_clk cell_7028 ( .C (CLK), .D (signal_9171), .Q (signal_9172) ) ;
    buf_clk cell_7036 ( .C (CLK), .D (signal_9179), .Q (signal_9180) ) ;
    buf_clk cell_7044 ( .C (CLK), .D (signal_9187), .Q (signal_9188) ) ;
    buf_clk cell_7052 ( .C (CLK), .D (signal_9195), .Q (signal_9196) ) ;
    buf_clk cell_7060 ( .C (CLK), .D (signal_9203), .Q (signal_9204) ) ;
    buf_clk cell_7068 ( .C (CLK), .D (signal_9211), .Q (signal_9212) ) ;
    buf_clk cell_7076 ( .C (CLK), .D (signal_9219), .Q (signal_9220) ) ;
    buf_clk cell_7084 ( .C (CLK), .D (signal_9227), .Q (signal_9228) ) ;
    buf_clk cell_7092 ( .C (CLK), .D (signal_9235), .Q (signal_9236) ) ;
    buf_clk cell_7100 ( .C (CLK), .D (signal_9243), .Q (signal_9244) ) ;
    buf_clk cell_7108 ( .C (CLK), .D (signal_9251), .Q (signal_9252) ) ;
    buf_clk cell_7116 ( .C (CLK), .D (signal_9259), .Q (signal_9260) ) ;
    buf_clk cell_7124 ( .C (CLK), .D (signal_9267), .Q (signal_9268) ) ;
    buf_clk cell_7132 ( .C (CLK), .D (signal_9275), .Q (signal_9276) ) ;
    buf_clk cell_7140 ( .C (CLK), .D (signal_9283), .Q (signal_9284) ) ;
    buf_clk cell_7148 ( .C (CLK), .D (signal_9291), .Q (signal_9292) ) ;
    buf_clk cell_7156 ( .C (CLK), .D (signal_9299), .Q (signal_9300) ) ;
    buf_clk cell_7164 ( .C (CLK), .D (signal_9307), .Q (signal_9308) ) ;
    buf_clk cell_7172 ( .C (CLK), .D (signal_9315), .Q (signal_9316) ) ;
    buf_clk cell_7180 ( .C (CLK), .D (signal_9323), .Q (signal_9324) ) ;
    buf_clk cell_7188 ( .C (CLK), .D (signal_9331), .Q (signal_9332) ) ;
    buf_clk cell_7196 ( .C (CLK), .D (signal_9339), .Q (signal_9340) ) ;
    buf_clk cell_7204 ( .C (CLK), .D (signal_9347), .Q (signal_9348) ) ;
    buf_clk cell_7212 ( .C (CLK), .D (signal_9355), .Q (signal_9356) ) ;
    buf_clk cell_7220 ( .C (CLK), .D (signal_9363), .Q (signal_9364) ) ;
    buf_clk cell_7228 ( .C (CLK), .D (signal_9371), .Q (signal_9372) ) ;
    buf_clk cell_7236 ( .C (CLK), .D (signal_9379), .Q (signal_9380) ) ;
    buf_clk cell_7244 ( .C (CLK), .D (signal_9387), .Q (signal_9388) ) ;
    buf_clk cell_7252 ( .C (CLK), .D (signal_9395), .Q (signal_9396) ) ;
    buf_clk cell_7260 ( .C (CLK), .D (signal_9403), .Q (signal_9404) ) ;
    buf_clk cell_7268 ( .C (CLK), .D (signal_9411), .Q (signal_9412) ) ;
    buf_clk cell_7276 ( .C (CLK), .D (signal_9419), .Q (signal_9420) ) ;
    buf_clk cell_7284 ( .C (CLK), .D (signal_9427), .Q (signal_9428) ) ;
    buf_clk cell_7292 ( .C (CLK), .D (signal_9435), .Q (signal_9436) ) ;
    buf_clk cell_7300 ( .C (CLK), .D (signal_9443), .Q (signal_9444) ) ;
    buf_clk cell_7308 ( .C (CLK), .D (signal_9451), .Q (signal_9452) ) ;
    buf_clk cell_7316 ( .C (CLK), .D (signal_9459), .Q (signal_9460) ) ;
    buf_clk cell_7324 ( .C (CLK), .D (signal_9467), .Q (signal_9468) ) ;
    buf_clk cell_7332 ( .C (CLK), .D (signal_9475), .Q (signal_9476) ) ;
    buf_clk cell_7340 ( .C (CLK), .D (signal_9483), .Q (signal_9484) ) ;
    buf_clk cell_7348 ( .C (CLK), .D (signal_9491), .Q (signal_9492) ) ;
    buf_clk cell_7356 ( .C (CLK), .D (signal_9499), .Q (signal_9500) ) ;
    buf_clk cell_7364 ( .C (CLK), .D (signal_9507), .Q (signal_9508) ) ;
    buf_clk cell_7372 ( .C (CLK), .D (signal_9515), .Q (signal_9516) ) ;
    buf_clk cell_7380 ( .C (CLK), .D (signal_9523), .Q (signal_9524) ) ;
    buf_clk cell_7388 ( .C (CLK), .D (signal_9531), .Q (signal_9532) ) ;
    buf_clk cell_7396 ( .C (CLK), .D (signal_9539), .Q (signal_9540) ) ;
    buf_clk cell_7404 ( .C (CLK), .D (signal_9547), .Q (signal_9548) ) ;
    buf_clk cell_7412 ( .C (CLK), .D (signal_9555), .Q (signal_9556) ) ;
    buf_clk cell_7420 ( .C (CLK), .D (signal_9563), .Q (signal_9564) ) ;
    buf_clk cell_7428 ( .C (CLK), .D (signal_9571), .Q (signal_9572) ) ;
    buf_clk cell_7436 ( .C (CLK), .D (signal_9579), .Q (signal_9580) ) ;
    buf_clk cell_7444 ( .C (CLK), .D (signal_9587), .Q (signal_9588) ) ;
    buf_clk cell_7452 ( .C (CLK), .D (signal_9595), .Q (signal_9596) ) ;
    buf_clk cell_7460 ( .C (CLK), .D (signal_9603), .Q (signal_9604) ) ;
    buf_clk cell_7468 ( .C (CLK), .D (signal_9611), .Q (signal_9612) ) ;
    buf_clk cell_7476 ( .C (CLK), .D (signal_9619), .Q (signal_9620) ) ;
    buf_clk cell_7484 ( .C (CLK), .D (signal_9627), .Q (signal_9628) ) ;
    buf_clk cell_7492 ( .C (CLK), .D (signal_9635), .Q (signal_9636) ) ;
    buf_clk cell_7500 ( .C (CLK), .D (signal_9643), .Q (signal_9644) ) ;
    buf_clk cell_7508 ( .C (CLK), .D (signal_9651), .Q (signal_9652) ) ;
    buf_clk cell_7516 ( .C (CLK), .D (signal_9659), .Q (signal_9660) ) ;
    buf_clk cell_7524 ( .C (CLK), .D (signal_9667), .Q (signal_9668) ) ;
    buf_clk cell_7532 ( .C (CLK), .D (signal_9675), .Q (signal_9676) ) ;
    buf_clk cell_7540 ( .C (CLK), .D (signal_9683), .Q (signal_9684) ) ;
    buf_clk cell_7548 ( .C (CLK), .D (signal_9691), .Q (signal_9692) ) ;
    buf_clk cell_7556 ( .C (CLK), .D (signal_9699), .Q (signal_9700) ) ;
    buf_clk cell_7604 ( .C (CLK), .D (signal_9747), .Q (signal_9748) ) ;
    buf_clk cell_7620 ( .C (CLK), .D (signal_9763), .Q (signal_9764) ) ;
    buf_clk cell_7636 ( .C (CLK), .D (signal_9779), .Q (signal_9780) ) ;
    buf_clk cell_7652 ( .C (CLK), .D (signal_9795), .Q (signal_9796) ) ;
    buf_clk cell_7668 ( .C (CLK), .D (signal_9811), .Q (signal_9812) ) ;
    buf_clk cell_7684 ( .C (CLK), .D (signal_9827), .Q (signal_9828) ) ;
    buf_clk cell_7700 ( .C (CLK), .D (signal_9843), .Q (signal_9844) ) ;
    buf_clk cell_7716 ( .C (CLK), .D (signal_9859), .Q (signal_9860) ) ;
    buf_clk cell_7732 ( .C (CLK), .D (signal_9875), .Q (signal_9876) ) ;
    buf_clk cell_7748 ( .C (CLK), .D (signal_9891), .Q (signal_9892) ) ;
    buf_clk cell_7756 ( .C (CLK), .D (signal_9899), .Q (signal_9900) ) ;
    buf_clk cell_7764 ( .C (CLK), .D (signal_9907), .Q (signal_9908) ) ;
    buf_clk cell_7772 ( .C (CLK), .D (signal_9915), .Q (signal_9916) ) ;
    buf_clk cell_7780 ( .C (CLK), .D (signal_9923), .Q (signal_9924) ) ;
    buf_clk cell_7788 ( .C (CLK), .D (signal_9931), .Q (signal_9932) ) ;
    buf_clk cell_7796 ( .C (CLK), .D (signal_9939), .Q (signal_9940) ) ;
    buf_clk cell_7804 ( .C (CLK), .D (signal_9947), .Q (signal_9948) ) ;
    buf_clk cell_7812 ( .C (CLK), .D (signal_9955), .Q (signal_9956) ) ;
    buf_clk cell_7820 ( .C (CLK), .D (signal_9963), .Q (signal_9964) ) ;
    buf_clk cell_7828 ( .C (CLK), .D (signal_9971), .Q (signal_9972) ) ;
    buf_clk cell_7836 ( .C (CLK), .D (signal_9979), .Q (signal_9980) ) ;
    buf_clk cell_7844 ( .C (CLK), .D (signal_9987), .Q (signal_9988) ) ;
    buf_clk cell_7852 ( .C (CLK), .D (signal_9995), .Q (signal_9996) ) ;
    buf_clk cell_7860 ( .C (CLK), .D (signal_10003), .Q (signal_10004) ) ;
    buf_clk cell_7868 ( .C (CLK), .D (signal_10011), .Q (signal_10012) ) ;
    buf_clk cell_7876 ( .C (CLK), .D (signal_10019), .Q (signal_10020) ) ;
    buf_clk cell_7884 ( .C (CLK), .D (signal_10027), .Q (signal_10028) ) ;
    buf_clk cell_7892 ( .C (CLK), .D (signal_10035), .Q (signal_10036) ) ;
    buf_clk cell_7900 ( .C (CLK), .D (signal_10043), .Q (signal_10044) ) ;
    buf_clk cell_7908 ( .C (CLK), .D (signal_10051), .Q (signal_10052) ) ;
    buf_clk cell_7916 ( .C (CLK), .D (signal_10059), .Q (signal_10060) ) ;
    buf_clk cell_7924 ( .C (CLK), .D (signal_10067), .Q (signal_10068) ) ;
    buf_clk cell_7932 ( .C (CLK), .D (signal_10075), .Q (signal_10076) ) ;
    buf_clk cell_7940 ( .C (CLK), .D (signal_10083), .Q (signal_10084) ) ;
    buf_clk cell_7956 ( .C (CLK), .D (signal_10099), .Q (signal_10100) ) ;

    /* cells in depth 16 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_39 ( .s (signal_5589), .b ({signal_2964, signal_1327}), .a ({signal_5621, signal_5605}), .c ({signal_2983, signal_1263}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_41 ( .s (signal_5629), .b ({signal_3004, signal_1325}), .a ({signal_5661, signal_5645}), .c ({signal_3018, signal_1261}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_43 ( .s (signal_5669), .b ({signal_2968, signal_1323}), .a ({signal_5701, signal_5685}), .c ({signal_2985, signal_1259}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_45 ( .s (signal_5669), .b ({signal_2967, signal_1321}), .a ({signal_5733, signal_5717}), .c ({signal_2987, signal_1257}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_47 ( .s (signal_5669), .b ({signal_2934, signal_1319}), .a ({signal_5741, signal_5737}), .c ({signal_2950, signal_1255}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_49 ( .s (signal_5669), .b ({signal_3012, signal_1317}), .a ({signal_5753, signal_5747}), .c ({signal_3019, signal_1253}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_51 ( .s (signal_5669), .b ({signal_2982, signal_1315}), .a ({signal_5765, signal_5759}), .c ({signal_2988, signal_1251}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_53 ( .s (signal_5669), .b ({signal_3016, signal_1313}), .a ({signal_5777, signal_5771}), .c ({signal_3020, signal_1249}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_55 ( .s (signal_5589), .b ({signal_3003, signal_1311}), .a ({signal_5809, signal_5793}), .c ({signal_3021, signal_1247}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_56 ( .s (signal_5589), .b ({signal_3083, signal_1310}), .a ({signal_5841, signal_5825}), .c ({signal_3100, signal_1246}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_58 ( .s (signal_5589), .b ({signal_3082, signal_1308}), .a ({signal_5873, signal_5857}), .c ({signal_3101, signal_1244}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_59 ( .s (signal_5589), .b ({signal_2966, signal_1307}), .a ({signal_5905, signal_5889}), .c ({signal_2989, signal_1243}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_60 ( .s (signal_5589), .b ({signal_3090, signal_1306}), .a ({signal_5937, signal_5921}), .c ({signal_3102, signal_1242}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_62 ( .s (signal_5589), .b ({signal_3047, signal_1304}), .a ({signal_5945, signal_5941}), .c ({signal_3061, signal_1240}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_63 ( .s (signal_5589), .b ({signal_2971, signal_1303}), .a ({signal_5961, signal_5953}), .c ({signal_2990, signal_1239}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_64 ( .s (signal_5589), .b ({signal_3054, signal_1302}), .a ({signal_5973, signal_5967}), .c ({signal_3062, signal_1238}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_66 ( .s (signal_5589), .b ({signal_3093, signal_1300}), .a ({signal_5989, signal_5981}), .c ({signal_3103, signal_1236}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_67 ( .s (signal_5629), .b ({signal_3015, signal_1299}), .a ({signal_6005, signal_5997}), .c ({signal_3023, signal_1235}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_68 ( .s (signal_5629), .b ({signal_3099, signal_1298}), .a ({signal_6013, signal_6009}), .c ({signal_3104, signal_1234}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_70 ( .s (signal_5629), .b ({signal_3098, signal_1296}), .a ({signal_6029, signal_6021}), .c ({signal_3105, signal_1232}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_71 ( .s (signal_5629), .b ({signal_3165, signal_1295}), .a ({signal_6061, signal_6045}), .c ({signal_3178, signal_1231}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_72 ( .s (signal_5629), .b ({signal_3167, signal_1294}), .a ({signal_6093, signal_6077}), .c ({signal_3179, signal_1230}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_73 ( .s (signal_5629), .b ({signal_3078, signal_1293}), .a ({signal_6125, signal_6109}), .c ({signal_3106, signal_1229}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_74 ( .s (signal_5629), .b ({signal_3123, signal_1292}), .a ({signal_6157, signal_6141}), .c ({signal_3137, signal_1228}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_75 ( .s (signal_5629), .b ({signal_3126, signal_1291}), .a ({signal_6189, signal_6173}), .c ({signal_3138, signal_1227}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_76 ( .s (signal_5629), .b ({signal_3128, signal_1290}), .a ({signal_6221, signal_6205}), .c ({signal_3139, signal_1226}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_77 ( .s (signal_5629), .b ({signal_3084, signal_1289}), .a ({signal_6253, signal_6237}), .c ({signal_3107, signal_1225}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_78 ( .s (signal_5629), .b ({signal_3127, signal_1288}), .a ({signal_6273, signal_6263}), .c ({signal_3140, signal_1224}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_79 ( .s (signal_5629), .b ({signal_3171, signal_1287}), .a ({signal_6285, signal_6279}), .c ({signal_3180, signal_1223}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_80 ( .s (signal_5589), .b ({signal_3173, signal_1286}), .a ({signal_6301, signal_6293}), .c ({signal_3181, signal_1222}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_81 ( .s (signal_5669), .b ({signal_3049, signal_1285}), .a ({signal_6321, signal_6311}), .c ({signal_3063, signal_1221}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_82 ( .s (signal_6337), .b ({signal_3092, signal_1284}), .a ({signal_6361, signal_6349}), .c ({signal_3108, signal_1220}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_83 ( .s (signal_5589), .b ({signal_3175, signal_1283}), .a ({signal_6377, signal_6369}), .c ({signal_3182, signal_1219}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_84 ( .s (signal_5669), .b ({signal_3177, signal_1282}), .a ({signal_6401, signal_6389}), .c ({signal_3183, signal_1218}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_85 ( .s (signal_5629), .b ({signal_3094, signal_1281}), .a ({signal_6429, signal_6415}), .c ({signal_3109, signal_1217}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_86 ( .s (signal_6337), .b ({signal_3096, signal_1280}), .a ({signal_6461, signal_6445}), .c ({signal_3110, signal_1216}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_87 ( .s (signal_6337), .b ({signal_3235, signal_1279}), .a ({signal_6493, signal_6477}), .c ({signal_3240, signal_1215}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_88 ( .s (signal_6337), .b ({signal_3252, signal_1278}), .a ({signal_6525, signal_6509}), .c ({signal_3256, signal_1214}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_89 ( .s (signal_6337), .b ({signal_3198, signal_1277}), .a ({signal_6557, signal_6541}), .c ({signal_3209, signal_1213}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_90 ( .s (signal_6337), .b ({signal_3164, signal_1276}), .a ({signal_6589, signal_6573}), .c ({signal_3184, signal_1212}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_91 ( .s (signal_6337), .b ({signal_3237, signal_1275}), .a ({signal_6621, signal_6605}), .c ({signal_3241, signal_1211}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_92 ( .s (signal_6337), .b ({signal_3253, signal_1274}), .a ({signal_6653, signal_6637}), .c ({signal_3257, signal_1210}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_93 ( .s (signal_5629), .b ({signal_3169, signal_1273}), .a ({signal_6685, signal_6669}), .c ({signal_3185, signal_1209}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_94 ( .s (signal_5589), .b ({signal_3168, signal_1272}), .a ({signal_6705, signal_6695}), .c ({signal_3186, signal_1208}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_95 ( .s (signal_5669), .b ({signal_3205, signal_1271}), .a ({signal_6721, signal_6713}), .c ({signal_3210, signal_1207}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_96 ( .s (signal_5629), .b ({signal_3254, signal_1270}), .a ({signal_6745, signal_6733}), .c ({signal_3258, signal_1206}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_97 ( .s (signal_5589), .b ({signal_3203, signal_1269}), .a ({signal_6773, signal_6759}), .c ({signal_3211, signal_1205}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_98 ( .s (signal_5669), .b ({signal_3129, signal_1268}), .a ({signal_6805, signal_6789}), .c ({signal_3141, signal_1204}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_99 ( .s (signal_5589), .b ({signal_3208, signal_1267}), .a ({signal_6817, signal_6811}), .c ({signal_3212, signal_1203}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_100 ( .s (signal_5669), .b ({signal_3255, signal_1266}), .a ({signal_6833, signal_6825}), .c ({signal_3259, signal_1202}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_101 ( .s (signal_5629), .b ({signal_3206, signal_1265}), .a ({signal_6853, signal_6843}), .c ({signal_3213, signal_1201}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_102 ( .s (signal_5629), .b ({signal_3174, signal_1264}), .a ({signal_6877, signal_6865}), .c ({signal_3187, signal_1200}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_103 ( .s (signal_6885), .b ({signal_2983, signal_1263}), .a ({signal_6917, signal_6901}), .c ({signal_3026, signal_1199}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_105 ( .s (signal_6885), .b ({signal_3018, signal_1261}), .a ({signal_6949, signal_6933}), .c ({signal_3065, signal_1197}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_107 ( .s (signal_6885), .b ({signal_2985, signal_1259}), .a ({signal_6981, signal_6965}), .c ({signal_3030, signal_1195}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_109 ( .s (signal_6885), .b ({signal_2987, signal_1257}), .a ({signal_7013, signal_6997}), .c ({signal_3034, signal_1193}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_111 ( .s (signal_6885), .b ({signal_2950, signal_1255}), .a ({signal_7045, signal_7029}), .c ({signal_2994, signal_1191}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_113 ( .s (signal_6885), .b ({signal_3019, signal_1253}), .a ({signal_7077, signal_7061}), .c ({signal_3067, signal_1189}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_115 ( .s (signal_6885), .b ({signal_2988, signal_1251}), .a ({signal_7109, signal_7093}), .c ({signal_3036, signal_1187}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_117 ( .s (signal_6885), .b ({signal_3020, signal_1249}), .a ({signal_7141, signal_7125}), .c ({signal_3069, signal_1185}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_119 ( .s (signal_6885), .b ({signal_3021, signal_1247}), .a ({signal_7173, signal_7157}), .c ({signal_3071, signal_1183}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_120 ( .s (signal_6885), .b ({signal_3100, signal_1246}), .a ({signal_7205, signal_7189}), .c ({signal_3143, signal_1182}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_122 ( .s (signal_6885), .b ({signal_3101, signal_1244}), .a ({signal_7237, signal_7221}), .c ({signal_3145, signal_1180}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_123 ( .s (signal_6885), .b ({signal_2989, signal_1243}), .a ({signal_7269, signal_7253}), .c ({signal_3038, signal_1179}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_124 ( .s (signal_6885), .b ({signal_3102, signal_1242}), .a ({signal_7301, signal_7285}), .c ({signal_3147, signal_1178}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_126 ( .s (signal_6885), .b ({signal_3061, signal_1240}), .a ({signal_7333, signal_7317}), .c ({signal_3116, signal_1176}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_127 ( .s (signal_6885), .b ({signal_2990, signal_1239}), .a ({signal_7365, signal_7349}), .c ({signal_3040, signal_1175}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_128 ( .s (signal_6885), .b ({signal_3062, signal_1238}), .a ({signal_7397, signal_7381}), .c ({signal_3118, signal_1174}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_130 ( .s (signal_6885), .b ({signal_3103, signal_1236}), .a ({signal_7429, signal_7413}), .c ({signal_3149, signal_1172}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_131 ( .s (signal_6885), .b ({signal_3023, signal_1235}), .a ({signal_7461, signal_7445}), .c ({signal_3075, signal_1171}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_132 ( .s (signal_6885), .b ({signal_3104, signal_1234}), .a ({signal_7493, signal_7477}), .c ({signal_3151, signal_1170}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_134 ( .s (signal_6885), .b ({signal_3105, signal_1232}), .a ({signal_7525, signal_7509}), .c ({signal_3153, signal_1168}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_135 ( .s (signal_6885), .b ({signal_3178, signal_1231}), .a ({signal_7557, signal_7541}), .c ({signal_3215, signal_1167}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_136 ( .s (signal_6885), .b ({signal_3179, signal_1230}), .a ({signal_7589, signal_7573}), .c ({signal_3217, signal_1166}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_137 ( .s (signal_6885), .b ({signal_3106, signal_1229}), .a ({signal_7621, signal_7605}), .c ({signal_3155, signal_1165}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_138 ( .s (signal_6885), .b ({signal_3137, signal_1228}), .a ({signal_7653, signal_7637}), .c ({signal_3189, signal_1164}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_139 ( .s (signal_6885), .b ({signal_3138, signal_1227}), .a ({signal_7685, signal_7669}), .c ({signal_3191, signal_1163}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_140 ( .s (signal_6885), .b ({signal_3139, signal_1226}), .a ({signal_7717, signal_7701}), .c ({signal_3193, signal_1162}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_141 ( .s (signal_6885), .b ({signal_3107, signal_1225}), .a ({signal_7749, signal_7733}), .c ({signal_3157, signal_1161}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_142 ( .s (signal_6885), .b ({signal_3140, signal_1224}), .a ({signal_7781, signal_7765}), .c ({signal_3195, signal_1160}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_143 ( .s (signal_6885), .b ({signal_3180, signal_1223}), .a ({signal_7813, signal_7797}), .c ({signal_3219, signal_1159}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_144 ( .s (signal_6885), .b ({signal_3181, signal_1222}), .a ({signal_7845, signal_7829}), .c ({signal_3221, signal_1158}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_145 ( .s (signal_6885), .b ({signal_3063, signal_1221}), .a ({signal_7877, signal_7861}), .c ({signal_3120, signal_1157}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_146 ( .s (signal_6885), .b ({signal_3108, signal_1220}), .a ({signal_7909, signal_7893}), .c ({signal_3159, signal_1156}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_147 ( .s (signal_6885), .b ({signal_3182, signal_1219}), .a ({signal_7941, signal_7925}), .c ({signal_3223, signal_1155}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_148 ( .s (signal_6885), .b ({signal_3183, signal_1218}), .a ({signal_7973, signal_7957}), .c ({signal_3225, signal_1154}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_149 ( .s (signal_6885), .b ({signal_3109, signal_1217}), .a ({signal_8005, signal_7989}), .c ({signal_3161, signal_1153}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_150 ( .s (signal_6885), .b ({signal_3110, signal_1216}), .a ({signal_8037, signal_8021}), .c ({signal_3163, signal_1152}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_151 ( .s (signal_6885), .b ({signal_3240, signal_1215}), .a ({signal_8069, signal_8053}), .c ({signal_3261, signal_1151}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_152 ( .s (signal_6885), .b ({signal_3256, signal_1214}), .a ({signal_8101, signal_8085}), .c ({signal_3265, signal_1150}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_153 ( .s (signal_6885), .b ({signal_3209, signal_1213}), .a ({signal_8133, signal_8117}), .c ({signal_3243, signal_1149}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_154 ( .s (signal_6885), .b ({signal_3184, signal_1212}), .a ({signal_8165, signal_8149}), .c ({signal_3227, signal_1148}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_155 ( .s (signal_6885), .b ({signal_3241, signal_1211}), .a ({signal_8197, signal_8181}), .c ({signal_3263, signal_1147}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_156 ( .s (signal_6885), .b ({signal_3257, signal_1210}), .a ({signal_8229, signal_8213}), .c ({signal_3267, signal_1146}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_157 ( .s (signal_6885), .b ({signal_3185, signal_1209}), .a ({signal_8261, signal_8245}), .c ({signal_3229, signal_1145}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_158 ( .s (signal_6885), .b ({signal_3186, signal_1208}), .a ({signal_8293, signal_8277}), .c ({signal_3231, signal_1144}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_159 ( .s (signal_6885), .b ({signal_3210, signal_1207}), .a ({signal_8325, signal_8309}), .c ({signal_3245, signal_1143}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_160 ( .s (signal_6885), .b ({signal_3258, signal_1206}), .a ({signal_8357, signal_8341}), .c ({signal_3269, signal_1142}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_161 ( .s (signal_6885), .b ({signal_3211, signal_1205}), .a ({signal_8389, signal_8373}), .c ({signal_3247, signal_1141}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_162 ( .s (signal_6885), .b ({signal_3141, signal_1204}), .a ({signal_8421, signal_8405}), .c ({signal_3197, signal_1140}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_163 ( .s (signal_6885), .b ({signal_3212, signal_1203}), .a ({signal_8453, signal_8437}), .c ({signal_3249, signal_1139}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_164 ( .s (signal_6885), .b ({signal_3259, signal_1202}), .a ({signal_8485, signal_8469}), .c ({signal_3271, signal_1138}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_165 ( .s (signal_6885), .b ({signal_3213, signal_1201}), .a ({signal_8517, signal_8501}), .c ({signal_3251, signal_1137}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_166 ( .s (signal_6885), .b ({signal_3187, signal_1200}), .a ({signal_8549, signal_8533}), .c ({signal_3233, signal_1136}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_762 ( .a ({signal_3121, signal_656}), .b ({signal_8565, signal_8557}), .c ({signal_3164, signal_1276}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_764 ( .a ({signal_3078, signal_1293}), .b ({signal_8581, signal_8573}), .c ({signal_3121, signal_656}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_765 ( .a ({signal_8597, signal_8589}), .b ({signal_3044, signal_659}), .c ({signal_3078, signal_1293}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_767 ( .a ({signal_3079, signal_661}), .b ({signal_3167, signal_1294}), .c ({signal_3198, signal_1277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_768 ( .a ({signal_3004, signal_1325}), .b ({signal_3044, signal_659}), .c ({signal_3079, signal_661}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_769 ( .a ({signal_3234, signal_662}), .b ({signal_3124, signal_663}), .c ({signal_3252, signal_1278}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_770 ( .a ({signal_3199, signal_664}), .b ({signal_8613, signal_8605}), .c ({signal_3234, signal_662}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_772 ( .a ({signal_3165, signal_1295}), .b ({signal_3166, signal_666}), .c ({signal_3199, signal_664}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_773 ( .a ({signal_3122, signal_667}), .b ({signal_8629, signal_8621}), .c ({signal_3165, signal_1295}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_775 ( .a ({signal_8645, signal_8637}), .b ({signal_3082, signal_1308}), .c ({signal_3122, signal_667}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_776 ( .a ({signal_3200, signal_669}), .b ({signal_2964, signal_1327}), .c ({signal_3235, signal_1279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_777 ( .a ({signal_3082, signal_1308}), .b ({signal_3166, signal_666}), .c ({signal_3200, signal_669}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_778 ( .a ({signal_8661, signal_8653}), .b ({signal_3123, signal_1292}), .c ({signal_3166, signal_666}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_779 ( .a ({signal_3080, signal_670}), .b ({signal_8677, signal_8669}), .c ({signal_3123, signal_1292}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_781 ( .a ({signal_8581, signal_8573}), .b ({signal_3004, signal_1325}), .c ({signal_3080, signal_670}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_790 ( .a ({signal_3081, signal_679}), .b ({signal_3124, signal_663}), .c ({signal_3167, signal_1294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_791 ( .a ({signal_3003, signal_1311}), .b ({signal_3082, signal_1308}), .c ({signal_3124, signal_663}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_792 ( .a ({signal_3042, signal_680}), .b ({signal_8693, signal_8685}), .c ({signal_3081, signal_679}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_794 ( .a ({signal_3005, signal_682}), .b ({signal_8709, signal_8701}), .c ({signal_3042, signal_680}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_795 ( .a ({signal_2947, signal_683}), .b ({signal_8725, signal_8717}), .c ({signal_3003, signal_1311}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_798 ( .a ({signal_3043, signal_685}), .b ({signal_8741, signal_8733}), .c ({signal_3082, signal_1308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_800 ( .a ({signal_3004, signal_1325}), .b ({signal_8757, signal_8749}), .c ({signal_3043, signal_685}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_801 ( .a ({signal_2941, signal_687}), .b ({signal_2962, signal_688}), .c ({signal_3004, signal_1325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_802 ( .a ({signal_2937, signal_689}), .b ({signal_8773, signal_8765}), .c ({signal_2962, signal_688}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_804 ( .a ({signal_8789, signal_8781}), .b ({signal_3044, signal_659}), .c ({signal_3083, signal_1310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_805 ( .a ({signal_2963, signal_690}), .b ({signal_3005, signal_682}), .c ({signal_3044, signal_659}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_806 ( .a ({signal_8805, signal_8797}), .b ({signal_2964, signal_1327}), .c ({signal_3005, signal_682}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_807 ( .a ({signal_8821, signal_8813}), .b ({signal_2937, signal_689}), .c ({signal_2963, signal_690}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_810 ( .a ({signal_2938, signal_691}), .b ({signal_8837, signal_8829}), .c ({signal_2964, signal_1327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_816 ( .a ({signal_3125, signal_694}), .b ({signal_8853, signal_8845}), .c ({signal_3168, signal_1272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_818 ( .a ({signal_3084, signal_1289}), .b ({signal_8869, signal_8861}), .c ({signal_3125, signal_694}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_819 ( .a ({signal_8885, signal_8877}), .b ({signal_3048, signal_697}), .c ({signal_3084, signal_1289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_821 ( .a ({signal_3085, signal_699}), .b ({signal_3128, signal_1290}), .c ({signal_3169, signal_1273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_822 ( .a ({signal_2967, signal_1321}), .b ({signal_3048, signal_697}), .c ({signal_3085, signal_699}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_823 ( .a ({signal_3236, signal_700}), .b ({signal_3088, signal_701}), .c ({signal_3253, signal_1274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_824 ( .a ({signal_3201, signal_702}), .b ({signal_8901, signal_8893}), .c ({signal_3236, signal_700}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_826 ( .a ({signal_3126, signal_1291}), .b ({signal_3170, signal_704}), .c ({signal_3201, signal_702}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_827 ( .a ({signal_3086, signal_705}), .b ({signal_8917, signal_8909}), .c ({signal_3126, signal_1291}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_829 ( .a ({signal_8933, signal_8925}), .b ({signal_3047, signal_1304}), .c ({signal_3086, signal_705}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_830 ( .a ({signal_3202, signal_707}), .b ({signal_2968, signal_1323}), .c ({signal_3237, signal_1275}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_831 ( .a ({signal_3047, signal_1304}), .b ({signal_3170, signal_704}), .c ({signal_3202, signal_707}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_832 ( .a ({signal_8949, signal_8941}), .b ({signal_3127, signal_1288}), .c ({signal_3170, signal_704}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_833 ( .a ({signal_3087, signal_708}), .b ({signal_8965, signal_8957}), .c ({signal_3127, signal_1288}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_835 ( .a ({signal_8869, signal_8861}), .b ({signal_2967, signal_1321}), .c ({signal_3087, signal_708}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_844 ( .a ({signal_3089, signal_717}), .b ({signal_3088, signal_701}), .c ({signal_3128, signal_1290}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_845 ( .a ({signal_2966, signal_1307}), .b ({signal_3047, signal_1304}), .c ({signal_3088, signal_701}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_846 ( .a ({signal_3046, signal_718}), .b ({signal_8981, signal_8973}), .c ({signal_3089, signal_717}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_848 ( .a ({signal_3009, signal_720}), .b ({signal_8997, signal_8989}), .c ({signal_3046, signal_718}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_849 ( .a ({signal_2917, signal_721}), .b ({signal_9013, signal_9005}), .c ({signal_2966, signal_1307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_852 ( .a ({signal_3008, signal_723}), .b ({signal_9029, signal_9021}), .c ({signal_3047, signal_1304}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_854 ( .a ({signal_2967, signal_1321}), .b ({signal_9045, signal_9037}), .c ({signal_3008, signal_723}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_855 ( .a ({signal_2942, signal_725}), .b ({signal_2928, signal_726}), .c ({signal_2967, signal_1321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_856 ( .a ({signal_2914, signal_727}), .b ({signal_9061, signal_9053}), .c ({signal_2928, signal_726}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_858 ( .a ({signal_9077, signal_9069}), .b ({signal_3048, signal_697}), .c ({signal_3090, signal_1306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_859 ( .a ({signal_2929, signal_728}), .b ({signal_3009, signal_720}), .c ({signal_3048, signal_697}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_860 ( .a ({signal_9093, signal_9085}), .b ({signal_2968, signal_1323}), .c ({signal_3009, signal_720}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_861 ( .a ({signal_9109, signal_9101}), .b ({signal_2914, signal_727}), .c ({signal_2929, signal_728}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_864 ( .a ({signal_2943, signal_729}), .b ({signal_9125, signal_9117}), .c ({signal_2968, signal_1323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_870 ( .a ({signal_3091, signal_732}), .b ({signal_9141, signal_9133}), .c ({signal_3129, signal_1268}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_872 ( .a ({signal_3049, signal_1285}), .b ({signal_9157, signal_9149}), .c ({signal_3091, signal_732}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_873 ( .a ({signal_9173, signal_9165}), .b ({signal_3013, signal_735}), .c ({signal_3049, signal_1285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_875 ( .a ({signal_3050, signal_737}), .b ({signal_3173, signal_1286}), .c ({signal_3203, signal_1269}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_876 ( .a ({signal_3012, signal_1317}), .b ({signal_3013, signal_735}), .c ({signal_3050, signal_737}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_877 ( .a ({signal_3238, signal_738}), .b ({signal_3132, signal_739}), .c ({signal_3254, signal_1270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_878 ( .a ({signal_3204, signal_740}), .b ({signal_9189, signal_9181}), .c ({signal_3238, signal_738}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_880 ( .a ({signal_3171, signal_1287}), .b ({signal_3131, signal_742}), .c ({signal_3204, signal_740}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_881 ( .a ({signal_3130, signal_743}), .b ({signal_9205, signal_9197}), .c ({signal_3171, signal_1287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_883 ( .a ({signal_9221, signal_9213}), .b ({signal_3093, signal_1300}), .c ({signal_3130, signal_743}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_884 ( .a ({signal_3172, signal_745}), .b ({signal_2934, signal_1319}), .c ({signal_3205, signal_1271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_885 ( .a ({signal_3093, signal_1300}), .b ({signal_3131, signal_742}), .c ({signal_3172, signal_745}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_886 ( .a ({signal_9237, signal_9229}), .b ({signal_3092, signal_1284}), .c ({signal_3131, signal_742}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_887 ( .a ({signal_3051, signal_746}), .b ({signal_9253, signal_9245}), .c ({signal_3092, signal_1284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_889 ( .a ({signal_9157, signal_9149}), .b ({signal_3012, signal_1317}), .c ({signal_3051, signal_746}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_898 ( .a ({signal_3052, signal_755}), .b ({signal_3132, signal_739}), .c ({signal_3173, signal_1286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_899 ( .a ({signal_2971, signal_1303}), .b ({signal_3093, signal_1300}), .c ({signal_3132, signal_739}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_900 ( .a ({signal_3011, signal_756}), .b ({signal_9269, signal_9261}), .c ({signal_3052, signal_755}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_902 ( .a ({signal_2973, signal_758}), .b ({signal_9285, signal_9277}), .c ({signal_3011, signal_756}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_903 ( .a ({signal_2946, signal_759}), .b ({signal_9301, signal_9293}), .c ({signal_2971, signal_1303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_906 ( .a ({signal_3053, signal_761}), .b ({signal_9317, signal_9309}), .c ({signal_3093, signal_1300}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_908 ( .a ({signal_3012, signal_1317}), .b ({signal_9333, signal_9325}), .c ({signal_3053, signal_761}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_909 ( .a ({signal_2944, signal_763}), .b ({signal_2972, signal_764}), .c ({signal_3012, signal_1317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_910 ( .a ({signal_2939, signal_765}), .b ({signal_9349, signal_9341}), .c ({signal_2972, signal_764}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_912 ( .a ({signal_9365, signal_9357}), .b ({signal_3013, signal_735}), .c ({signal_3054, signal_1302}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_913 ( .a ({signal_2974, signal_766}), .b ({signal_2973, signal_758}), .c ({signal_3013, signal_735}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_914 ( .a ({signal_9381, signal_9373}), .b ({signal_2934, signal_1319}), .c ({signal_2973, signal_758}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_915 ( .a ({signal_9397, signal_9389}), .b ({signal_2939, signal_765}), .c ({signal_2974, signal_766}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_918 ( .a ({signal_2915, signal_767}), .b ({signal_9413, signal_9405}), .c ({signal_2934, signal_1319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_924 ( .a ({signal_3133, signal_770}), .b ({signal_9429, signal_9421}), .c ({signal_3174, signal_1264}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_926 ( .a ({signal_3094, signal_1281}), .b ({signal_9445, signal_9437}), .c ({signal_3133, signal_770}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_927 ( .a ({signal_9461, signal_9453}), .b ({signal_3058, signal_773}), .c ({signal_3094, signal_1281}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_929 ( .a ({signal_3095, signal_775}), .b ({signal_3177, signal_1282}), .c ({signal_3206, signal_1265}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_930 ( .a ({signal_3016, signal_1313}), .b ({signal_3058, signal_773}), .c ({signal_3095, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_931 ( .a ({signal_3239, signal_776}), .b ({signal_3136, signal_777}), .c ({signal_3255, signal_1266}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_932 ( .a ({signal_3207, signal_778}), .b ({signal_9477, signal_9469}), .c ({signal_3239, signal_776}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_934 ( .a ({signal_3175, signal_1283}), .b ({signal_3135, signal_780}), .c ({signal_3207, signal_778}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_935 ( .a ({signal_3134, signal_781}), .b ({signal_9493, signal_9485}), .c ({signal_3175, signal_1283}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_937 ( .a ({signal_9509, signal_9501}), .b ({signal_3098, signal_1296}), .c ({signal_3134, signal_781}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_938 ( .a ({signal_3176, signal_783}), .b ({signal_2982, signal_1315}), .c ({signal_3208, signal_1267}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_939 ( .a ({signal_3098, signal_1296}), .b ({signal_3135, signal_780}), .c ({signal_3176, signal_783}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_940 ( .a ({signal_9525, signal_9517}), .b ({signal_3096, signal_1280}), .c ({signal_3135, signal_780}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_941 ( .a ({signal_3055, signal_784}), .b ({signal_9541, signal_9533}), .c ({signal_3096, signal_1280}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_943 ( .a ({signal_9445, signal_9437}), .b ({signal_3016, signal_1313}), .c ({signal_3055, signal_784}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_952 ( .a ({signal_3097, signal_793}), .b ({signal_3136, signal_777}), .c ({signal_3177, signal_1282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_953 ( .a ({signal_3015, signal_1299}), .b ({signal_3098, signal_1296}), .c ({signal_3136, signal_777}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_954 ( .a ({signal_3056, signal_794}), .b ({signal_9557, signal_9549}), .c ({signal_3097, signal_793}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_956 ( .a ({signal_3017, signal_796}), .b ({signal_9573, signal_9565}), .c ({signal_3056, signal_794}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_957 ( .a ({signal_2948, signal_797}), .b ({signal_9589, signal_9581}), .c ({signal_3015, signal_1299}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_960 ( .a ({signal_3057, signal_799}), .b ({signal_9605, signal_9597}), .c ({signal_3098, signal_1296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_962 ( .a ({signal_3016, signal_1313}), .b ({signal_9621, signal_9613}), .c ({signal_3057, signal_799}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_963 ( .a ({signal_2916, signal_801}), .b ({signal_2980, signal_802}), .c ({signal_3016, signal_1313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_964 ( .a ({signal_2940, signal_803}), .b ({signal_9637, signal_9629}), .c ({signal_2980, signal_802}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_966 ( .a ({signal_9653, signal_9645}), .b ({signal_3058, signal_773}), .c ({signal_3099, signal_1298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_967 ( .a ({signal_2981, signal_804}), .b ({signal_3017, signal_796}), .c ({signal_3058, signal_773}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_968 ( .a ({signal_9669, signal_9661}), .b ({signal_2982, signal_1315}), .c ({signal_3017, signal_796}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_969 ( .a ({signal_9685, signal_9677}), .b ({signal_2940, signal_803}), .c ({signal_2981, signal_804}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_972 ( .a ({signal_2945, signal_805}), .b ({signal_9701, signal_9693}), .c ({signal_2982, signal_1315}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1710 ( .s ({signal_5959, signal_5951}), .b ({signal_2871, signal_1823}), .a ({signal_2870, signal_1822}), .clk (CLK), .r (Fresh[582]), .c ({signal_2914, signal_727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1711 ( .s ({signal_9705, signal_9703}), .b ({signal_2891, signal_1825}), .a ({signal_2890, signal_1824}), .clk (CLK), .r (Fresh[583]), .c ({signal_2937, signal_689}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1712 ( .s ({signal_9721, signal_9713}), .b ({signal_2893, signal_1827}), .a ({signal_2892, signal_1826}), .clk (CLK), .r (Fresh[584]), .c ({signal_2938, signal_691}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1713 ( .s ({signal_6003, signal_5995}), .b ({signal_2895, signal_1829}), .a ({signal_2894, signal_1828}), .clk (CLK), .r (Fresh[585]), .c ({signal_2939, signal_765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1714 ( .s ({signal_6271, signal_6261}), .b ({signal_2897, signal_1831}), .a ({signal_2896, signal_1830}), .clk (CLK), .r (Fresh[586]), .c ({signal_2940, signal_803}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1715 ( .s ({signal_9721, signal_9713}), .b ({signal_2899, signal_1833}), .a ({signal_2898, signal_1832}), .clk (CLK), .r (Fresh[587]), .c ({signal_2941, signal_687}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1716 ( .s ({signal_9729, signal_9725}), .b ({signal_2901, signal_1835}), .a ({signal_2900, signal_1834}), .clk (CLK), .r (Fresh[588]), .c ({signal_2942, signal_725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1717 ( .s ({signal_5959, signal_5951}), .b ({signal_2903, signal_1837}), .a ({signal_2902, signal_1836}), .clk (CLK), .r (Fresh[589]), .c ({signal_2943, signal_729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1718 ( .s ({signal_5739, signal_5735}), .b ({signal_2905, signal_1839}), .a ({signal_2904, signal_1838}), .clk (CLK), .r (Fresh[590]), .c ({signal_2944, signal_763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1719 ( .s ({signal_6003, signal_5995}), .b ({signal_2873, signal_1841}), .a ({signal_2872, signal_1840}), .clk (CLK), .r (Fresh[591]), .c ({signal_2915, signal_767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1720 ( .s ({signal_5763, signal_5757}), .b ({signal_2875, signal_1843}), .a ({signal_2874, signal_1842}), .clk (CLK), .r (Fresh[592]), .c ({signal_2916, signal_801}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1721 ( .s ({signal_9733, signal_9731}), .b ({signal_2907, signal_1845}), .a ({signal_2906, signal_1844}), .clk (CLK), .r (Fresh[593]), .c ({signal_2945, signal_805}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1722 ( .s ({signal_5959, signal_5951}), .b ({signal_2877, signal_1847}), .a ({signal_2876, signal_1846}), .clk (CLK), .r (Fresh[594]), .c ({signal_2917, signal_721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1723 ( .s ({signal_6003, signal_5995}), .b ({signal_2909, signal_1849}), .a ({signal_2908, signal_1848}), .clk (CLK), .r (Fresh[595]), .c ({signal_2946, signal_759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1724 ( .s ({signal_9705, signal_9703}), .b ({signal_2911, signal_1851}), .a ({signal_2910, signal_1850}), .clk (CLK), .r (Fresh[596]), .c ({signal_2947, signal_683}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1725 ( .s ({signal_6271, signal_6261}), .b ({signal_2913, signal_1853}), .a ({signal_2912, signal_1852}), .clk (CLK), .r (Fresh[597]), .c ({signal_2948, signal_797}) ) ;
    buf_clk cell_3445 ( .C (CLK), .D (signal_5588), .Q (signal_5589) ) ;
    buf_clk cell_3461 ( .C (CLK), .D (signal_5604), .Q (signal_5605) ) ;
    buf_clk cell_3477 ( .C (CLK), .D (signal_5620), .Q (signal_5621) ) ;
    buf_clk cell_3485 ( .C (CLK), .D (signal_5628), .Q (signal_5629) ) ;
    buf_clk cell_3501 ( .C (CLK), .D (signal_5644), .Q (signal_5645) ) ;
    buf_clk cell_3517 ( .C (CLK), .D (signal_5660), .Q (signal_5661) ) ;
    buf_clk cell_3525 ( .C (CLK), .D (signal_5668), .Q (signal_5669) ) ;
    buf_clk cell_3541 ( .C (CLK), .D (signal_5684), .Q (signal_5685) ) ;
    buf_clk cell_3557 ( .C (CLK), .D (signal_5700), .Q (signal_5701) ) ;
    buf_clk cell_3573 ( .C (CLK), .D (signal_5716), .Q (signal_5717) ) ;
    buf_clk cell_3589 ( .C (CLK), .D (signal_5732), .Q (signal_5733) ) ;
    buf_clk cell_3593 ( .C (CLK), .D (signal_5736), .Q (signal_5737) ) ;
    buf_clk cell_3597 ( .C (CLK), .D (signal_5740), .Q (signal_5741) ) ;
    buf_clk cell_3603 ( .C (CLK), .D (signal_5746), .Q (signal_5747) ) ;
    buf_clk cell_3609 ( .C (CLK), .D (signal_5752), .Q (signal_5753) ) ;
    buf_clk cell_3615 ( .C (CLK), .D (signal_5758), .Q (signal_5759) ) ;
    buf_clk cell_3621 ( .C (CLK), .D (signal_5764), .Q (signal_5765) ) ;
    buf_clk cell_3627 ( .C (CLK), .D (signal_5770), .Q (signal_5771) ) ;
    buf_clk cell_3633 ( .C (CLK), .D (signal_5776), .Q (signal_5777) ) ;
    buf_clk cell_3649 ( .C (CLK), .D (signal_5792), .Q (signal_5793) ) ;
    buf_clk cell_3665 ( .C (CLK), .D (signal_5808), .Q (signal_5809) ) ;
    buf_clk cell_3681 ( .C (CLK), .D (signal_5824), .Q (signal_5825) ) ;
    buf_clk cell_3697 ( .C (CLK), .D (signal_5840), .Q (signal_5841) ) ;
    buf_clk cell_3713 ( .C (CLK), .D (signal_5856), .Q (signal_5857) ) ;
    buf_clk cell_3729 ( .C (CLK), .D (signal_5872), .Q (signal_5873) ) ;
    buf_clk cell_3745 ( .C (CLK), .D (signal_5888), .Q (signal_5889) ) ;
    buf_clk cell_3761 ( .C (CLK), .D (signal_5904), .Q (signal_5905) ) ;
    buf_clk cell_3777 ( .C (CLK), .D (signal_5920), .Q (signal_5921) ) ;
    buf_clk cell_3793 ( .C (CLK), .D (signal_5936), .Q (signal_5937) ) ;
    buf_clk cell_3797 ( .C (CLK), .D (signal_5940), .Q (signal_5941) ) ;
    buf_clk cell_3801 ( .C (CLK), .D (signal_5944), .Q (signal_5945) ) ;
    buf_clk cell_3809 ( .C (CLK), .D (signal_5952), .Q (signal_5953) ) ;
    buf_clk cell_3817 ( .C (CLK), .D (signal_5960), .Q (signal_5961) ) ;
    buf_clk cell_3823 ( .C (CLK), .D (signal_5966), .Q (signal_5967) ) ;
    buf_clk cell_3829 ( .C (CLK), .D (signal_5972), .Q (signal_5973) ) ;
    buf_clk cell_3837 ( .C (CLK), .D (signal_5980), .Q (signal_5981) ) ;
    buf_clk cell_3845 ( .C (CLK), .D (signal_5988), .Q (signal_5989) ) ;
    buf_clk cell_3853 ( .C (CLK), .D (signal_5996), .Q (signal_5997) ) ;
    buf_clk cell_3861 ( .C (CLK), .D (signal_6004), .Q (signal_6005) ) ;
    buf_clk cell_3865 ( .C (CLK), .D (signal_6008), .Q (signal_6009) ) ;
    buf_clk cell_3869 ( .C (CLK), .D (signal_6012), .Q (signal_6013) ) ;
    buf_clk cell_3877 ( .C (CLK), .D (signal_6020), .Q (signal_6021) ) ;
    buf_clk cell_3885 ( .C (CLK), .D (signal_6028), .Q (signal_6029) ) ;
    buf_clk cell_3901 ( .C (CLK), .D (signal_6044), .Q (signal_6045) ) ;
    buf_clk cell_3917 ( .C (CLK), .D (signal_6060), .Q (signal_6061) ) ;
    buf_clk cell_3933 ( .C (CLK), .D (signal_6076), .Q (signal_6077) ) ;
    buf_clk cell_3949 ( .C (CLK), .D (signal_6092), .Q (signal_6093) ) ;
    buf_clk cell_3965 ( .C (CLK), .D (signal_6108), .Q (signal_6109) ) ;
    buf_clk cell_3981 ( .C (CLK), .D (signal_6124), .Q (signal_6125) ) ;
    buf_clk cell_3997 ( .C (CLK), .D (signal_6140), .Q (signal_6141) ) ;
    buf_clk cell_4013 ( .C (CLK), .D (signal_6156), .Q (signal_6157) ) ;
    buf_clk cell_4029 ( .C (CLK), .D (signal_6172), .Q (signal_6173) ) ;
    buf_clk cell_4045 ( .C (CLK), .D (signal_6188), .Q (signal_6189) ) ;
    buf_clk cell_4061 ( .C (CLK), .D (signal_6204), .Q (signal_6205) ) ;
    buf_clk cell_4077 ( .C (CLK), .D (signal_6220), .Q (signal_6221) ) ;
    buf_clk cell_4093 ( .C (CLK), .D (signal_6236), .Q (signal_6237) ) ;
    buf_clk cell_4109 ( .C (CLK), .D (signal_6252), .Q (signal_6253) ) ;
    buf_clk cell_4119 ( .C (CLK), .D (signal_6262), .Q (signal_6263) ) ;
    buf_clk cell_4129 ( .C (CLK), .D (signal_6272), .Q (signal_6273) ) ;
    buf_clk cell_4135 ( .C (CLK), .D (signal_6278), .Q (signal_6279) ) ;
    buf_clk cell_4141 ( .C (CLK), .D (signal_6284), .Q (signal_6285) ) ;
    buf_clk cell_4149 ( .C (CLK), .D (signal_6292), .Q (signal_6293) ) ;
    buf_clk cell_4157 ( .C (CLK), .D (signal_6300), .Q (signal_6301) ) ;
    buf_clk cell_4167 ( .C (CLK), .D (signal_6310), .Q (signal_6311) ) ;
    buf_clk cell_4177 ( .C (CLK), .D (signal_6320), .Q (signal_6321) ) ;
    buf_clk cell_4193 ( .C (CLK), .D (signal_6336), .Q (signal_6337) ) ;
    buf_clk cell_4205 ( .C (CLK), .D (signal_6348), .Q (signal_6349) ) ;
    buf_clk cell_4217 ( .C (CLK), .D (signal_6360), .Q (signal_6361) ) ;
    buf_clk cell_4225 ( .C (CLK), .D (signal_6368), .Q (signal_6369) ) ;
    buf_clk cell_4233 ( .C (CLK), .D (signal_6376), .Q (signal_6377) ) ;
    buf_clk cell_4245 ( .C (CLK), .D (signal_6388), .Q (signal_6389) ) ;
    buf_clk cell_4257 ( .C (CLK), .D (signal_6400), .Q (signal_6401) ) ;
    buf_clk cell_4271 ( .C (CLK), .D (signal_6414), .Q (signal_6415) ) ;
    buf_clk cell_4285 ( .C (CLK), .D (signal_6428), .Q (signal_6429) ) ;
    buf_clk cell_4301 ( .C (CLK), .D (signal_6444), .Q (signal_6445) ) ;
    buf_clk cell_4317 ( .C (CLK), .D (signal_6460), .Q (signal_6461) ) ;
    buf_clk cell_4333 ( .C (CLK), .D (signal_6476), .Q (signal_6477) ) ;
    buf_clk cell_4349 ( .C (CLK), .D (signal_6492), .Q (signal_6493) ) ;
    buf_clk cell_4365 ( .C (CLK), .D (signal_6508), .Q (signal_6509) ) ;
    buf_clk cell_4381 ( .C (CLK), .D (signal_6524), .Q (signal_6525) ) ;
    buf_clk cell_4397 ( .C (CLK), .D (signal_6540), .Q (signal_6541) ) ;
    buf_clk cell_4413 ( .C (CLK), .D (signal_6556), .Q (signal_6557) ) ;
    buf_clk cell_4429 ( .C (CLK), .D (signal_6572), .Q (signal_6573) ) ;
    buf_clk cell_4445 ( .C (CLK), .D (signal_6588), .Q (signal_6589) ) ;
    buf_clk cell_4461 ( .C (CLK), .D (signal_6604), .Q (signal_6605) ) ;
    buf_clk cell_4477 ( .C (CLK), .D (signal_6620), .Q (signal_6621) ) ;
    buf_clk cell_4493 ( .C (CLK), .D (signal_6636), .Q (signal_6637) ) ;
    buf_clk cell_4509 ( .C (CLK), .D (signal_6652), .Q (signal_6653) ) ;
    buf_clk cell_4525 ( .C (CLK), .D (signal_6668), .Q (signal_6669) ) ;
    buf_clk cell_4541 ( .C (CLK), .D (signal_6684), .Q (signal_6685) ) ;
    buf_clk cell_4551 ( .C (CLK), .D (signal_6694), .Q (signal_6695) ) ;
    buf_clk cell_4561 ( .C (CLK), .D (signal_6704), .Q (signal_6705) ) ;
    buf_clk cell_4569 ( .C (CLK), .D (signal_6712), .Q (signal_6713) ) ;
    buf_clk cell_4577 ( .C (CLK), .D (signal_6720), .Q (signal_6721) ) ;
    buf_clk cell_4589 ( .C (CLK), .D (signal_6732), .Q (signal_6733) ) ;
    buf_clk cell_4601 ( .C (CLK), .D (signal_6744), .Q (signal_6745) ) ;
    buf_clk cell_4615 ( .C (CLK), .D (signal_6758), .Q (signal_6759) ) ;
    buf_clk cell_4629 ( .C (CLK), .D (signal_6772), .Q (signal_6773) ) ;
    buf_clk cell_4645 ( .C (CLK), .D (signal_6788), .Q (signal_6789) ) ;
    buf_clk cell_4661 ( .C (CLK), .D (signal_6804), .Q (signal_6805) ) ;
    buf_clk cell_4667 ( .C (CLK), .D (signal_6810), .Q (signal_6811) ) ;
    buf_clk cell_4673 ( .C (CLK), .D (signal_6816), .Q (signal_6817) ) ;
    buf_clk cell_4681 ( .C (CLK), .D (signal_6824), .Q (signal_6825) ) ;
    buf_clk cell_4689 ( .C (CLK), .D (signal_6832), .Q (signal_6833) ) ;
    buf_clk cell_4699 ( .C (CLK), .D (signal_6842), .Q (signal_6843) ) ;
    buf_clk cell_4709 ( .C (CLK), .D (signal_6852), .Q (signal_6853) ) ;
    buf_clk cell_4721 ( .C (CLK), .D (signal_6864), .Q (signal_6865) ) ;
    buf_clk cell_4733 ( .C (CLK), .D (signal_6876), .Q (signal_6877) ) ;
    buf_clk cell_4741 ( .C (CLK), .D (signal_6884), .Q (signal_6885) ) ;
    buf_clk cell_4757 ( .C (CLK), .D (signal_6900), .Q (signal_6901) ) ;
    buf_clk cell_4773 ( .C (CLK), .D (signal_6916), .Q (signal_6917) ) ;
    buf_clk cell_4789 ( .C (CLK), .D (signal_6932), .Q (signal_6933) ) ;
    buf_clk cell_4805 ( .C (CLK), .D (signal_6948), .Q (signal_6949) ) ;
    buf_clk cell_4821 ( .C (CLK), .D (signal_6964), .Q (signal_6965) ) ;
    buf_clk cell_4837 ( .C (CLK), .D (signal_6980), .Q (signal_6981) ) ;
    buf_clk cell_4853 ( .C (CLK), .D (signal_6996), .Q (signal_6997) ) ;
    buf_clk cell_4869 ( .C (CLK), .D (signal_7012), .Q (signal_7013) ) ;
    buf_clk cell_4885 ( .C (CLK), .D (signal_7028), .Q (signal_7029) ) ;
    buf_clk cell_4901 ( .C (CLK), .D (signal_7044), .Q (signal_7045) ) ;
    buf_clk cell_4917 ( .C (CLK), .D (signal_7060), .Q (signal_7061) ) ;
    buf_clk cell_4933 ( .C (CLK), .D (signal_7076), .Q (signal_7077) ) ;
    buf_clk cell_4949 ( .C (CLK), .D (signal_7092), .Q (signal_7093) ) ;
    buf_clk cell_4965 ( .C (CLK), .D (signal_7108), .Q (signal_7109) ) ;
    buf_clk cell_4981 ( .C (CLK), .D (signal_7124), .Q (signal_7125) ) ;
    buf_clk cell_4997 ( .C (CLK), .D (signal_7140), .Q (signal_7141) ) ;
    buf_clk cell_5013 ( .C (CLK), .D (signal_7156), .Q (signal_7157) ) ;
    buf_clk cell_5029 ( .C (CLK), .D (signal_7172), .Q (signal_7173) ) ;
    buf_clk cell_5045 ( .C (CLK), .D (signal_7188), .Q (signal_7189) ) ;
    buf_clk cell_5061 ( .C (CLK), .D (signal_7204), .Q (signal_7205) ) ;
    buf_clk cell_5077 ( .C (CLK), .D (signal_7220), .Q (signal_7221) ) ;
    buf_clk cell_5093 ( .C (CLK), .D (signal_7236), .Q (signal_7237) ) ;
    buf_clk cell_5109 ( .C (CLK), .D (signal_7252), .Q (signal_7253) ) ;
    buf_clk cell_5125 ( .C (CLK), .D (signal_7268), .Q (signal_7269) ) ;
    buf_clk cell_5141 ( .C (CLK), .D (signal_7284), .Q (signal_7285) ) ;
    buf_clk cell_5157 ( .C (CLK), .D (signal_7300), .Q (signal_7301) ) ;
    buf_clk cell_5173 ( .C (CLK), .D (signal_7316), .Q (signal_7317) ) ;
    buf_clk cell_5189 ( .C (CLK), .D (signal_7332), .Q (signal_7333) ) ;
    buf_clk cell_5205 ( .C (CLK), .D (signal_7348), .Q (signal_7349) ) ;
    buf_clk cell_5221 ( .C (CLK), .D (signal_7364), .Q (signal_7365) ) ;
    buf_clk cell_5237 ( .C (CLK), .D (signal_7380), .Q (signal_7381) ) ;
    buf_clk cell_5253 ( .C (CLK), .D (signal_7396), .Q (signal_7397) ) ;
    buf_clk cell_5269 ( .C (CLK), .D (signal_7412), .Q (signal_7413) ) ;
    buf_clk cell_5285 ( .C (CLK), .D (signal_7428), .Q (signal_7429) ) ;
    buf_clk cell_5301 ( .C (CLK), .D (signal_7444), .Q (signal_7445) ) ;
    buf_clk cell_5317 ( .C (CLK), .D (signal_7460), .Q (signal_7461) ) ;
    buf_clk cell_5333 ( .C (CLK), .D (signal_7476), .Q (signal_7477) ) ;
    buf_clk cell_5349 ( .C (CLK), .D (signal_7492), .Q (signal_7493) ) ;
    buf_clk cell_5365 ( .C (CLK), .D (signal_7508), .Q (signal_7509) ) ;
    buf_clk cell_5381 ( .C (CLK), .D (signal_7524), .Q (signal_7525) ) ;
    buf_clk cell_5397 ( .C (CLK), .D (signal_7540), .Q (signal_7541) ) ;
    buf_clk cell_5413 ( .C (CLK), .D (signal_7556), .Q (signal_7557) ) ;
    buf_clk cell_5429 ( .C (CLK), .D (signal_7572), .Q (signal_7573) ) ;
    buf_clk cell_5445 ( .C (CLK), .D (signal_7588), .Q (signal_7589) ) ;
    buf_clk cell_5461 ( .C (CLK), .D (signal_7604), .Q (signal_7605) ) ;
    buf_clk cell_5477 ( .C (CLK), .D (signal_7620), .Q (signal_7621) ) ;
    buf_clk cell_5493 ( .C (CLK), .D (signal_7636), .Q (signal_7637) ) ;
    buf_clk cell_5509 ( .C (CLK), .D (signal_7652), .Q (signal_7653) ) ;
    buf_clk cell_5525 ( .C (CLK), .D (signal_7668), .Q (signal_7669) ) ;
    buf_clk cell_5541 ( .C (CLK), .D (signal_7684), .Q (signal_7685) ) ;
    buf_clk cell_5557 ( .C (CLK), .D (signal_7700), .Q (signal_7701) ) ;
    buf_clk cell_5573 ( .C (CLK), .D (signal_7716), .Q (signal_7717) ) ;
    buf_clk cell_5589 ( .C (CLK), .D (signal_7732), .Q (signal_7733) ) ;
    buf_clk cell_5605 ( .C (CLK), .D (signal_7748), .Q (signal_7749) ) ;
    buf_clk cell_5621 ( .C (CLK), .D (signal_7764), .Q (signal_7765) ) ;
    buf_clk cell_5637 ( .C (CLK), .D (signal_7780), .Q (signal_7781) ) ;
    buf_clk cell_5653 ( .C (CLK), .D (signal_7796), .Q (signal_7797) ) ;
    buf_clk cell_5669 ( .C (CLK), .D (signal_7812), .Q (signal_7813) ) ;
    buf_clk cell_5685 ( .C (CLK), .D (signal_7828), .Q (signal_7829) ) ;
    buf_clk cell_5701 ( .C (CLK), .D (signal_7844), .Q (signal_7845) ) ;
    buf_clk cell_5717 ( .C (CLK), .D (signal_7860), .Q (signal_7861) ) ;
    buf_clk cell_5733 ( .C (CLK), .D (signal_7876), .Q (signal_7877) ) ;
    buf_clk cell_5749 ( .C (CLK), .D (signal_7892), .Q (signal_7893) ) ;
    buf_clk cell_5765 ( .C (CLK), .D (signal_7908), .Q (signal_7909) ) ;
    buf_clk cell_5781 ( .C (CLK), .D (signal_7924), .Q (signal_7925) ) ;
    buf_clk cell_5797 ( .C (CLK), .D (signal_7940), .Q (signal_7941) ) ;
    buf_clk cell_5813 ( .C (CLK), .D (signal_7956), .Q (signal_7957) ) ;
    buf_clk cell_5829 ( .C (CLK), .D (signal_7972), .Q (signal_7973) ) ;
    buf_clk cell_5845 ( .C (CLK), .D (signal_7988), .Q (signal_7989) ) ;
    buf_clk cell_5861 ( .C (CLK), .D (signal_8004), .Q (signal_8005) ) ;
    buf_clk cell_5877 ( .C (CLK), .D (signal_8020), .Q (signal_8021) ) ;
    buf_clk cell_5893 ( .C (CLK), .D (signal_8036), .Q (signal_8037) ) ;
    buf_clk cell_5909 ( .C (CLK), .D (signal_8052), .Q (signal_8053) ) ;
    buf_clk cell_5925 ( .C (CLK), .D (signal_8068), .Q (signal_8069) ) ;
    buf_clk cell_5941 ( .C (CLK), .D (signal_8084), .Q (signal_8085) ) ;
    buf_clk cell_5957 ( .C (CLK), .D (signal_8100), .Q (signal_8101) ) ;
    buf_clk cell_5973 ( .C (CLK), .D (signal_8116), .Q (signal_8117) ) ;
    buf_clk cell_5989 ( .C (CLK), .D (signal_8132), .Q (signal_8133) ) ;
    buf_clk cell_6005 ( .C (CLK), .D (signal_8148), .Q (signal_8149) ) ;
    buf_clk cell_6021 ( .C (CLK), .D (signal_8164), .Q (signal_8165) ) ;
    buf_clk cell_6037 ( .C (CLK), .D (signal_8180), .Q (signal_8181) ) ;
    buf_clk cell_6053 ( .C (CLK), .D (signal_8196), .Q (signal_8197) ) ;
    buf_clk cell_6069 ( .C (CLK), .D (signal_8212), .Q (signal_8213) ) ;
    buf_clk cell_6085 ( .C (CLK), .D (signal_8228), .Q (signal_8229) ) ;
    buf_clk cell_6101 ( .C (CLK), .D (signal_8244), .Q (signal_8245) ) ;
    buf_clk cell_6117 ( .C (CLK), .D (signal_8260), .Q (signal_8261) ) ;
    buf_clk cell_6133 ( .C (CLK), .D (signal_8276), .Q (signal_8277) ) ;
    buf_clk cell_6149 ( .C (CLK), .D (signal_8292), .Q (signal_8293) ) ;
    buf_clk cell_6165 ( .C (CLK), .D (signal_8308), .Q (signal_8309) ) ;
    buf_clk cell_6181 ( .C (CLK), .D (signal_8324), .Q (signal_8325) ) ;
    buf_clk cell_6197 ( .C (CLK), .D (signal_8340), .Q (signal_8341) ) ;
    buf_clk cell_6213 ( .C (CLK), .D (signal_8356), .Q (signal_8357) ) ;
    buf_clk cell_6229 ( .C (CLK), .D (signal_8372), .Q (signal_8373) ) ;
    buf_clk cell_6245 ( .C (CLK), .D (signal_8388), .Q (signal_8389) ) ;
    buf_clk cell_6261 ( .C (CLK), .D (signal_8404), .Q (signal_8405) ) ;
    buf_clk cell_6277 ( .C (CLK), .D (signal_8420), .Q (signal_8421) ) ;
    buf_clk cell_6293 ( .C (CLK), .D (signal_8436), .Q (signal_8437) ) ;
    buf_clk cell_6309 ( .C (CLK), .D (signal_8452), .Q (signal_8453) ) ;
    buf_clk cell_6325 ( .C (CLK), .D (signal_8468), .Q (signal_8469) ) ;
    buf_clk cell_6341 ( .C (CLK), .D (signal_8484), .Q (signal_8485) ) ;
    buf_clk cell_6357 ( .C (CLK), .D (signal_8500), .Q (signal_8501) ) ;
    buf_clk cell_6373 ( .C (CLK), .D (signal_8516), .Q (signal_8517) ) ;
    buf_clk cell_6389 ( .C (CLK), .D (signal_8532), .Q (signal_8533) ) ;
    buf_clk cell_6405 ( .C (CLK), .D (signal_8548), .Q (signal_8549) ) ;
    buf_clk cell_6413 ( .C (CLK), .D (signal_8556), .Q (signal_8557) ) ;
    buf_clk cell_6421 ( .C (CLK), .D (signal_8564), .Q (signal_8565) ) ;
    buf_clk cell_6429 ( .C (CLK), .D (signal_8572), .Q (signal_8573) ) ;
    buf_clk cell_6437 ( .C (CLK), .D (signal_8580), .Q (signal_8581) ) ;
    buf_clk cell_6445 ( .C (CLK), .D (signal_8588), .Q (signal_8589) ) ;
    buf_clk cell_6453 ( .C (CLK), .D (signal_8596), .Q (signal_8597) ) ;
    buf_clk cell_6461 ( .C (CLK), .D (signal_8604), .Q (signal_8605) ) ;
    buf_clk cell_6469 ( .C (CLK), .D (signal_8612), .Q (signal_8613) ) ;
    buf_clk cell_6477 ( .C (CLK), .D (signal_8620), .Q (signal_8621) ) ;
    buf_clk cell_6485 ( .C (CLK), .D (signal_8628), .Q (signal_8629) ) ;
    buf_clk cell_6493 ( .C (CLK), .D (signal_8636), .Q (signal_8637) ) ;
    buf_clk cell_6501 ( .C (CLK), .D (signal_8644), .Q (signal_8645) ) ;
    buf_clk cell_6509 ( .C (CLK), .D (signal_8652), .Q (signal_8653) ) ;
    buf_clk cell_6517 ( .C (CLK), .D (signal_8660), .Q (signal_8661) ) ;
    buf_clk cell_6525 ( .C (CLK), .D (signal_8668), .Q (signal_8669) ) ;
    buf_clk cell_6533 ( .C (CLK), .D (signal_8676), .Q (signal_8677) ) ;
    buf_clk cell_6541 ( .C (CLK), .D (signal_8684), .Q (signal_8685) ) ;
    buf_clk cell_6549 ( .C (CLK), .D (signal_8692), .Q (signal_8693) ) ;
    buf_clk cell_6557 ( .C (CLK), .D (signal_8700), .Q (signal_8701) ) ;
    buf_clk cell_6565 ( .C (CLK), .D (signal_8708), .Q (signal_8709) ) ;
    buf_clk cell_6573 ( .C (CLK), .D (signal_8716), .Q (signal_8717) ) ;
    buf_clk cell_6581 ( .C (CLK), .D (signal_8724), .Q (signal_8725) ) ;
    buf_clk cell_6589 ( .C (CLK), .D (signal_8732), .Q (signal_8733) ) ;
    buf_clk cell_6597 ( .C (CLK), .D (signal_8740), .Q (signal_8741) ) ;
    buf_clk cell_6605 ( .C (CLK), .D (signal_8748), .Q (signal_8749) ) ;
    buf_clk cell_6613 ( .C (CLK), .D (signal_8756), .Q (signal_8757) ) ;
    buf_clk cell_6621 ( .C (CLK), .D (signal_8764), .Q (signal_8765) ) ;
    buf_clk cell_6629 ( .C (CLK), .D (signal_8772), .Q (signal_8773) ) ;
    buf_clk cell_6637 ( .C (CLK), .D (signal_8780), .Q (signal_8781) ) ;
    buf_clk cell_6645 ( .C (CLK), .D (signal_8788), .Q (signal_8789) ) ;
    buf_clk cell_6653 ( .C (CLK), .D (signal_8796), .Q (signal_8797) ) ;
    buf_clk cell_6661 ( .C (CLK), .D (signal_8804), .Q (signal_8805) ) ;
    buf_clk cell_6669 ( .C (CLK), .D (signal_8812), .Q (signal_8813) ) ;
    buf_clk cell_6677 ( .C (CLK), .D (signal_8820), .Q (signal_8821) ) ;
    buf_clk cell_6685 ( .C (CLK), .D (signal_8828), .Q (signal_8829) ) ;
    buf_clk cell_6693 ( .C (CLK), .D (signal_8836), .Q (signal_8837) ) ;
    buf_clk cell_6701 ( .C (CLK), .D (signal_8844), .Q (signal_8845) ) ;
    buf_clk cell_6709 ( .C (CLK), .D (signal_8852), .Q (signal_8853) ) ;
    buf_clk cell_6717 ( .C (CLK), .D (signal_8860), .Q (signal_8861) ) ;
    buf_clk cell_6725 ( .C (CLK), .D (signal_8868), .Q (signal_8869) ) ;
    buf_clk cell_6733 ( .C (CLK), .D (signal_8876), .Q (signal_8877) ) ;
    buf_clk cell_6741 ( .C (CLK), .D (signal_8884), .Q (signal_8885) ) ;
    buf_clk cell_6749 ( .C (CLK), .D (signal_8892), .Q (signal_8893) ) ;
    buf_clk cell_6757 ( .C (CLK), .D (signal_8900), .Q (signal_8901) ) ;
    buf_clk cell_6765 ( .C (CLK), .D (signal_8908), .Q (signal_8909) ) ;
    buf_clk cell_6773 ( .C (CLK), .D (signal_8916), .Q (signal_8917) ) ;
    buf_clk cell_6781 ( .C (CLK), .D (signal_8924), .Q (signal_8925) ) ;
    buf_clk cell_6789 ( .C (CLK), .D (signal_8932), .Q (signal_8933) ) ;
    buf_clk cell_6797 ( .C (CLK), .D (signal_8940), .Q (signal_8941) ) ;
    buf_clk cell_6805 ( .C (CLK), .D (signal_8948), .Q (signal_8949) ) ;
    buf_clk cell_6813 ( .C (CLK), .D (signal_8956), .Q (signal_8957) ) ;
    buf_clk cell_6821 ( .C (CLK), .D (signal_8964), .Q (signal_8965) ) ;
    buf_clk cell_6829 ( .C (CLK), .D (signal_8972), .Q (signal_8973) ) ;
    buf_clk cell_6837 ( .C (CLK), .D (signal_8980), .Q (signal_8981) ) ;
    buf_clk cell_6845 ( .C (CLK), .D (signal_8988), .Q (signal_8989) ) ;
    buf_clk cell_6853 ( .C (CLK), .D (signal_8996), .Q (signal_8997) ) ;
    buf_clk cell_6861 ( .C (CLK), .D (signal_9004), .Q (signal_9005) ) ;
    buf_clk cell_6869 ( .C (CLK), .D (signal_9012), .Q (signal_9013) ) ;
    buf_clk cell_6877 ( .C (CLK), .D (signal_9020), .Q (signal_9021) ) ;
    buf_clk cell_6885 ( .C (CLK), .D (signal_9028), .Q (signal_9029) ) ;
    buf_clk cell_6893 ( .C (CLK), .D (signal_9036), .Q (signal_9037) ) ;
    buf_clk cell_6901 ( .C (CLK), .D (signal_9044), .Q (signal_9045) ) ;
    buf_clk cell_6909 ( .C (CLK), .D (signal_9052), .Q (signal_9053) ) ;
    buf_clk cell_6917 ( .C (CLK), .D (signal_9060), .Q (signal_9061) ) ;
    buf_clk cell_6925 ( .C (CLK), .D (signal_9068), .Q (signal_9069) ) ;
    buf_clk cell_6933 ( .C (CLK), .D (signal_9076), .Q (signal_9077) ) ;
    buf_clk cell_6941 ( .C (CLK), .D (signal_9084), .Q (signal_9085) ) ;
    buf_clk cell_6949 ( .C (CLK), .D (signal_9092), .Q (signal_9093) ) ;
    buf_clk cell_6957 ( .C (CLK), .D (signal_9100), .Q (signal_9101) ) ;
    buf_clk cell_6965 ( .C (CLK), .D (signal_9108), .Q (signal_9109) ) ;
    buf_clk cell_6973 ( .C (CLK), .D (signal_9116), .Q (signal_9117) ) ;
    buf_clk cell_6981 ( .C (CLK), .D (signal_9124), .Q (signal_9125) ) ;
    buf_clk cell_6989 ( .C (CLK), .D (signal_9132), .Q (signal_9133) ) ;
    buf_clk cell_6997 ( .C (CLK), .D (signal_9140), .Q (signal_9141) ) ;
    buf_clk cell_7005 ( .C (CLK), .D (signal_9148), .Q (signal_9149) ) ;
    buf_clk cell_7013 ( .C (CLK), .D (signal_9156), .Q (signal_9157) ) ;
    buf_clk cell_7021 ( .C (CLK), .D (signal_9164), .Q (signal_9165) ) ;
    buf_clk cell_7029 ( .C (CLK), .D (signal_9172), .Q (signal_9173) ) ;
    buf_clk cell_7037 ( .C (CLK), .D (signal_9180), .Q (signal_9181) ) ;
    buf_clk cell_7045 ( .C (CLK), .D (signal_9188), .Q (signal_9189) ) ;
    buf_clk cell_7053 ( .C (CLK), .D (signal_9196), .Q (signal_9197) ) ;
    buf_clk cell_7061 ( .C (CLK), .D (signal_9204), .Q (signal_9205) ) ;
    buf_clk cell_7069 ( .C (CLK), .D (signal_9212), .Q (signal_9213) ) ;
    buf_clk cell_7077 ( .C (CLK), .D (signal_9220), .Q (signal_9221) ) ;
    buf_clk cell_7085 ( .C (CLK), .D (signal_9228), .Q (signal_9229) ) ;
    buf_clk cell_7093 ( .C (CLK), .D (signal_9236), .Q (signal_9237) ) ;
    buf_clk cell_7101 ( .C (CLK), .D (signal_9244), .Q (signal_9245) ) ;
    buf_clk cell_7109 ( .C (CLK), .D (signal_9252), .Q (signal_9253) ) ;
    buf_clk cell_7117 ( .C (CLK), .D (signal_9260), .Q (signal_9261) ) ;
    buf_clk cell_7125 ( .C (CLK), .D (signal_9268), .Q (signal_9269) ) ;
    buf_clk cell_7133 ( .C (CLK), .D (signal_9276), .Q (signal_9277) ) ;
    buf_clk cell_7141 ( .C (CLK), .D (signal_9284), .Q (signal_9285) ) ;
    buf_clk cell_7149 ( .C (CLK), .D (signal_9292), .Q (signal_9293) ) ;
    buf_clk cell_7157 ( .C (CLK), .D (signal_9300), .Q (signal_9301) ) ;
    buf_clk cell_7165 ( .C (CLK), .D (signal_9308), .Q (signal_9309) ) ;
    buf_clk cell_7173 ( .C (CLK), .D (signal_9316), .Q (signal_9317) ) ;
    buf_clk cell_7181 ( .C (CLK), .D (signal_9324), .Q (signal_9325) ) ;
    buf_clk cell_7189 ( .C (CLK), .D (signal_9332), .Q (signal_9333) ) ;
    buf_clk cell_7197 ( .C (CLK), .D (signal_9340), .Q (signal_9341) ) ;
    buf_clk cell_7205 ( .C (CLK), .D (signal_9348), .Q (signal_9349) ) ;
    buf_clk cell_7213 ( .C (CLK), .D (signal_9356), .Q (signal_9357) ) ;
    buf_clk cell_7221 ( .C (CLK), .D (signal_9364), .Q (signal_9365) ) ;
    buf_clk cell_7229 ( .C (CLK), .D (signal_9372), .Q (signal_9373) ) ;
    buf_clk cell_7237 ( .C (CLK), .D (signal_9380), .Q (signal_9381) ) ;
    buf_clk cell_7245 ( .C (CLK), .D (signal_9388), .Q (signal_9389) ) ;
    buf_clk cell_7253 ( .C (CLK), .D (signal_9396), .Q (signal_9397) ) ;
    buf_clk cell_7261 ( .C (CLK), .D (signal_9404), .Q (signal_9405) ) ;
    buf_clk cell_7269 ( .C (CLK), .D (signal_9412), .Q (signal_9413) ) ;
    buf_clk cell_7277 ( .C (CLK), .D (signal_9420), .Q (signal_9421) ) ;
    buf_clk cell_7285 ( .C (CLK), .D (signal_9428), .Q (signal_9429) ) ;
    buf_clk cell_7293 ( .C (CLK), .D (signal_9436), .Q (signal_9437) ) ;
    buf_clk cell_7301 ( .C (CLK), .D (signal_9444), .Q (signal_9445) ) ;
    buf_clk cell_7309 ( .C (CLK), .D (signal_9452), .Q (signal_9453) ) ;
    buf_clk cell_7317 ( .C (CLK), .D (signal_9460), .Q (signal_9461) ) ;
    buf_clk cell_7325 ( .C (CLK), .D (signal_9468), .Q (signal_9469) ) ;
    buf_clk cell_7333 ( .C (CLK), .D (signal_9476), .Q (signal_9477) ) ;
    buf_clk cell_7341 ( .C (CLK), .D (signal_9484), .Q (signal_9485) ) ;
    buf_clk cell_7349 ( .C (CLK), .D (signal_9492), .Q (signal_9493) ) ;
    buf_clk cell_7357 ( .C (CLK), .D (signal_9500), .Q (signal_9501) ) ;
    buf_clk cell_7365 ( .C (CLK), .D (signal_9508), .Q (signal_9509) ) ;
    buf_clk cell_7373 ( .C (CLK), .D (signal_9516), .Q (signal_9517) ) ;
    buf_clk cell_7381 ( .C (CLK), .D (signal_9524), .Q (signal_9525) ) ;
    buf_clk cell_7389 ( .C (CLK), .D (signal_9532), .Q (signal_9533) ) ;
    buf_clk cell_7397 ( .C (CLK), .D (signal_9540), .Q (signal_9541) ) ;
    buf_clk cell_7405 ( .C (CLK), .D (signal_9548), .Q (signal_9549) ) ;
    buf_clk cell_7413 ( .C (CLK), .D (signal_9556), .Q (signal_9557) ) ;
    buf_clk cell_7421 ( .C (CLK), .D (signal_9564), .Q (signal_9565) ) ;
    buf_clk cell_7429 ( .C (CLK), .D (signal_9572), .Q (signal_9573) ) ;
    buf_clk cell_7437 ( .C (CLK), .D (signal_9580), .Q (signal_9581) ) ;
    buf_clk cell_7445 ( .C (CLK), .D (signal_9588), .Q (signal_9589) ) ;
    buf_clk cell_7453 ( .C (CLK), .D (signal_9596), .Q (signal_9597) ) ;
    buf_clk cell_7461 ( .C (CLK), .D (signal_9604), .Q (signal_9605) ) ;
    buf_clk cell_7469 ( .C (CLK), .D (signal_9612), .Q (signal_9613) ) ;
    buf_clk cell_7477 ( .C (CLK), .D (signal_9620), .Q (signal_9621) ) ;
    buf_clk cell_7485 ( .C (CLK), .D (signal_9628), .Q (signal_9629) ) ;
    buf_clk cell_7493 ( .C (CLK), .D (signal_9636), .Q (signal_9637) ) ;
    buf_clk cell_7501 ( .C (CLK), .D (signal_9644), .Q (signal_9645) ) ;
    buf_clk cell_7509 ( .C (CLK), .D (signal_9652), .Q (signal_9653) ) ;
    buf_clk cell_7517 ( .C (CLK), .D (signal_9660), .Q (signal_9661) ) ;
    buf_clk cell_7525 ( .C (CLK), .D (signal_9668), .Q (signal_9669) ) ;
    buf_clk cell_7533 ( .C (CLK), .D (signal_9676), .Q (signal_9677) ) ;
    buf_clk cell_7541 ( .C (CLK), .D (signal_9684), .Q (signal_9685) ) ;
    buf_clk cell_7549 ( .C (CLK), .D (signal_9692), .Q (signal_9693) ) ;
    buf_clk cell_7557 ( .C (CLK), .D (signal_9700), .Q (signal_9701) ) ;
    buf_clk cell_7605 ( .C (CLK), .D (signal_9748), .Q (signal_9749) ) ;
    buf_clk cell_7621 ( .C (CLK), .D (signal_9764), .Q (signal_9765) ) ;
    buf_clk cell_7637 ( .C (CLK), .D (signal_9780), .Q (signal_9781) ) ;
    buf_clk cell_7653 ( .C (CLK), .D (signal_9796), .Q (signal_9797) ) ;
    buf_clk cell_7669 ( .C (CLK), .D (signal_9812), .Q (signal_9813) ) ;
    buf_clk cell_7685 ( .C (CLK), .D (signal_9828), .Q (signal_9829) ) ;
    buf_clk cell_7701 ( .C (CLK), .D (signal_9844), .Q (signal_9845) ) ;
    buf_clk cell_7717 ( .C (CLK), .D (signal_9860), .Q (signal_9861) ) ;
    buf_clk cell_7733 ( .C (CLK), .D (signal_9876), .Q (signal_9877) ) ;
    buf_clk cell_7749 ( .C (CLK), .D (signal_9892), .Q (signal_9893) ) ;
    buf_clk cell_7757 ( .C (CLK), .D (signal_9900), .Q (signal_9901) ) ;
    buf_clk cell_7765 ( .C (CLK), .D (signal_9908), .Q (signal_9909) ) ;
    buf_clk cell_7773 ( .C (CLK), .D (signal_9916), .Q (signal_9917) ) ;
    buf_clk cell_7781 ( .C (CLK), .D (signal_9924), .Q (signal_9925) ) ;
    buf_clk cell_7789 ( .C (CLK), .D (signal_9932), .Q (signal_9933) ) ;
    buf_clk cell_7797 ( .C (CLK), .D (signal_9940), .Q (signal_9941) ) ;
    buf_clk cell_7805 ( .C (CLK), .D (signal_9948), .Q (signal_9949) ) ;
    buf_clk cell_7813 ( .C (CLK), .D (signal_9956), .Q (signal_9957) ) ;
    buf_clk cell_7821 ( .C (CLK), .D (signal_9964), .Q (signal_9965) ) ;
    buf_clk cell_7829 ( .C (CLK), .D (signal_9972), .Q (signal_9973) ) ;
    buf_clk cell_7837 ( .C (CLK), .D (signal_9980), .Q (signal_9981) ) ;
    buf_clk cell_7845 ( .C (CLK), .D (signal_9988), .Q (signal_9989) ) ;
    buf_clk cell_7853 ( .C (CLK), .D (signal_9996), .Q (signal_9997) ) ;
    buf_clk cell_7861 ( .C (CLK), .D (signal_10004), .Q (signal_10005) ) ;
    buf_clk cell_7869 ( .C (CLK), .D (signal_10012), .Q (signal_10013) ) ;
    buf_clk cell_7877 ( .C (CLK), .D (signal_10020), .Q (signal_10021) ) ;
    buf_clk cell_7885 ( .C (CLK), .D (signal_10028), .Q (signal_10029) ) ;
    buf_clk cell_7893 ( .C (CLK), .D (signal_10036), .Q (signal_10037) ) ;
    buf_clk cell_7901 ( .C (CLK), .D (signal_10044), .Q (signal_10045) ) ;
    buf_clk cell_7909 ( .C (CLK), .D (signal_10052), .Q (signal_10053) ) ;
    buf_clk cell_7917 ( .C (CLK), .D (signal_10060), .Q (signal_10061) ) ;
    buf_clk cell_7925 ( .C (CLK), .D (signal_10068), .Q (signal_10069) ) ;
    buf_clk cell_7933 ( .C (CLK), .D (signal_10076), .Q (signal_10077) ) ;
    buf_clk cell_7941 ( .C (CLK), .D (signal_10084), .Q (signal_10085) ) ;
    buf_clk cell_7957 ( .C (CLK), .D (signal_10100), .Q (signal_10101) ) ;

    /* register cells */
    DFF_X1 cell_979 ( .CK (CLK), .D (signal_9749), .Q (signal_808), .QN () ) ;
    DFF_X1 cell_981 ( .CK (CLK), .D (signal_9765), .Q (signal_307), .QN () ) ;
    DFF_X1 cell_983 ( .CK (CLK), .D (signal_9781), .Q (signal_304), .QN () ) ;
    DFF_X1 cell_985 ( .CK (CLK), .D (signal_9797), .Q (signal_288), .QN () ) ;
    DFF_X1 cell_987 ( .CK (CLK), .D (signal_9813), .Q (signal_879), .QN () ) ;
    DFF_X1 cell_989 ( .CK (CLK), .D (signal_9829), .Q (signal_878), .QN () ) ;
    DFF_X1 cell_991 ( .CK (CLK), .D (signal_9845), .Q (signal_877), .QN () ) ;
    DFF_X1 cell_993 ( .CK (CLK), .D (signal_9861), .Q (signal_876), .QN () ) ;
    DFF_X1 cell_995 ( .CK (CLK), .D (signal_9877), .Q (signal_875), .QN () ) ;
    DFF_X1 cell_997 ( .CK (CLK), .D (signal_9893), .Q (signal_874), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_999 ( .clk (CLK), .D ({signal_3026, signal_1199}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1001 ( .clk (CLK), .D ({signal_9909, signal_9901}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1003 ( .clk (CLK), .D ({signal_3065, signal_1197}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1005 ( .clk (CLK), .D ({signal_9925, signal_9917}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1007 ( .clk (CLK), .D ({signal_3030, signal_1195}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1009 ( .clk (CLK), .D ({signal_9941, signal_9933}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1011 ( .clk (CLK), .D ({signal_3034, signal_1193}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1013 ( .clk (CLK), .D ({signal_9957, signal_9949}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1015 ( .clk (CLK), .D ({signal_2994, signal_1191}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1017 ( .clk (CLK), .D ({signal_9973, signal_9965}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1019 ( .clk (CLK), .D ({signal_3067, signal_1189}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1021 ( .clk (CLK), .D ({signal_9989, signal_9981}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1023 ( .clk (CLK), .D ({signal_3036, signal_1187}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1025 ( .clk (CLK), .D ({signal_10005, signal_9997}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1027 ( .clk (CLK), .D ({signal_3069, signal_1185}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1029 ( .clk (CLK), .D ({signal_10021, signal_10013}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1031 ( .clk (CLK), .D ({signal_3071, signal_1183}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1033 ( .clk (CLK), .D ({signal_3143, signal_1182}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1035 ( .clk (CLK), .D ({signal_10037, signal_10029}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1037 ( .clk (CLK), .D ({signal_3145, signal_1180}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1039 ( .clk (CLK), .D ({signal_3038, signal_1179}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1041 ( .clk (CLK), .D ({signal_3147, signal_1178}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1043 ( .clk (CLK), .D ({signal_10053, signal_10045}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1045 ( .clk (CLK), .D ({signal_3116, signal_1176}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1047 ( .clk (CLK), .D ({signal_3040, signal_1175}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1049 ( .clk (CLK), .D ({signal_3118, signal_1174}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1051 ( .clk (CLK), .D ({signal_10069, signal_10061}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1053 ( .clk (CLK), .D ({signal_3149, signal_1172}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1055 ( .clk (CLK), .D ({signal_3075, signal_1171}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1057 ( .clk (CLK), .D ({signal_3151, signal_1170}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1059 ( .clk (CLK), .D ({signal_10085, signal_10077}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1061 ( .clk (CLK), .D ({signal_3153, signal_1168}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1063 ( .clk (CLK), .D ({signal_3215, signal_1167}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1065 ( .clk (CLK), .D ({signal_3217, signal_1166}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1067 ( .clk (CLK), .D ({signal_3155, signal_1165}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1069 ( .clk (CLK), .D ({signal_3189, signal_1164}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1071 ( .clk (CLK), .D ({signal_3191, signal_1163}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1073 ( .clk (CLK), .D ({signal_3193, signal_1162}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1075 ( .clk (CLK), .D ({signal_3157, signal_1161}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1077 ( .clk (CLK), .D ({signal_3195, signal_1160}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1079 ( .clk (CLK), .D ({signal_3219, signal_1159}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1081 ( .clk (CLK), .D ({signal_3221, signal_1158}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1083 ( .clk (CLK), .D ({signal_3120, signal_1157}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1085 ( .clk (CLK), .D ({signal_3159, signal_1156}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1087 ( .clk (CLK), .D ({signal_3223, signal_1155}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1089 ( .clk (CLK), .D ({signal_3225, signal_1154}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1091 ( .clk (CLK), .D ({signal_3161, signal_1153}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1093 ( .clk (CLK), .D ({signal_3163, signal_1152}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1095 ( .clk (CLK), .D ({signal_3261, signal_1151}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1097 ( .clk (CLK), .D ({signal_3265, signal_1150}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1099 ( .clk (CLK), .D ({signal_3243, signal_1149}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1101 ( .clk (CLK), .D ({signal_3227, signal_1148}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1103 ( .clk (CLK), .D ({signal_3263, signal_1147}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1105 ( .clk (CLK), .D ({signal_3267, signal_1146}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1107 ( .clk (CLK), .D ({signal_3229, signal_1145}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1109 ( .clk (CLK), .D ({signal_3231, signal_1144}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1111 ( .clk (CLK), .D ({signal_3245, signal_1143}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1113 ( .clk (CLK), .D ({signal_3269, signal_1142}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1115 ( .clk (CLK), .D ({signal_3247, signal_1141}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1117 ( .clk (CLK), .D ({signal_3197, signal_1140}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1119 ( .clk (CLK), .D ({signal_3249, signal_1139}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1121 ( .clk (CLK), .D ({signal_3271, signal_1138}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1123 ( .clk (CLK), .D ({signal_3251, signal_1137}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1125 ( .clk (CLK), .D ({signal_3233, signal_1136}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 cell_1127 ( .CK (CLK), .D (signal_10101), .Q (OUT_done), .QN () ) ;
endmodule
