/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d1 (SI_s0, clk, SI_s1, Fresh, SO_s0, SO_s1);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [878:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2393 ;
    wire signal_2395 ;
    wire signal_2397 ;
    wire signal_2399 ;
    wire signal_2401 ;
    wire signal_2403 ;
    wire signal_2405 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;
    wire signal_4813 ;
    wire signal_4814 ;
    wire signal_4815 ;
    wire signal_4816 ;
    wire signal_4817 ;
    wire signal_4818 ;
    wire signal_4819 ;
    wire signal_4820 ;
    wire signal_4821 ;
    wire signal_4822 ;
    wire signal_4823 ;
    wire signal_4824 ;
    wire signal_4825 ;
    wire signal_4826 ;
    wire signal_4827 ;
    wire signal_4828 ;
    wire signal_4829 ;
    wire signal_4830 ;
    wire signal_4831 ;
    wire signal_4832 ;
    wire signal_4833 ;
    wire signal_4834 ;
    wire signal_4835 ;
    wire signal_4836 ;
    wire signal_4837 ;
    wire signal_4838 ;
    wire signal_4839 ;
    wire signal_4840 ;
    wire signal_4841 ;
    wire signal_4842 ;
    wire signal_4843 ;
    wire signal_4844 ;
    wire signal_4845 ;
    wire signal_4846 ;
    wire signal_4847 ;
    wire signal_4848 ;
    wire signal_4849 ;
    wire signal_4850 ;
    wire signal_4851 ;
    wire signal_4852 ;
    wire signal_4853 ;
    wire signal_4854 ;
    wire signal_4855 ;
    wire signal_4856 ;
    wire signal_4857 ;
    wire signal_4858 ;
    wire signal_4859 ;
    wire signal_4860 ;
    wire signal_4861 ;
    wire signal_4862 ;
    wire signal_4863 ;
    wire signal_4864 ;
    wire signal_4865 ;
    wire signal_4866 ;
    wire signal_4867 ;
    wire signal_4868 ;
    wire signal_4869 ;
    wire signal_4870 ;
    wire signal_4871 ;
    wire signal_4872 ;
    wire signal_4873 ;
    wire signal_4874 ;
    wire signal_4875 ;
    wire signal_4876 ;
    wire signal_4877 ;
    wire signal_4878 ;
    wire signal_4879 ;
    wire signal_4880 ;
    wire signal_4881 ;
    wire signal_4882 ;
    wire signal_4883 ;
    wire signal_4884 ;
    wire signal_4885 ;
    wire signal_4886 ;
    wire signal_4887 ;
    wire signal_4888 ;
    wire signal_4889 ;
    wire signal_4890 ;
    wire signal_4891 ;
    wire signal_4892 ;
    wire signal_4893 ;
    wire signal_4894 ;
    wire signal_4895 ;
    wire signal_4896 ;
    wire signal_4897 ;
    wire signal_4898 ;
    wire signal_4899 ;
    wire signal_4900 ;
    wire signal_4901 ;
    wire signal_4902 ;
    wire signal_4903 ;
    wire signal_4904 ;
    wire signal_4905 ;
    wire signal_4906 ;
    wire signal_4907 ;
    wire signal_4908 ;
    wire signal_4909 ;
    wire signal_4910 ;
    wire signal_4911 ;
    wire signal_4912 ;
    wire signal_4913 ;
    wire signal_4914 ;
    wire signal_4915 ;
    wire signal_4916 ;
    wire signal_4917 ;
    wire signal_4918 ;
    wire signal_4919 ;
    wire signal_4920 ;
    wire signal_4921 ;
    wire signal_4922 ;
    wire signal_4923 ;
    wire signal_4924 ;
    wire signal_4925 ;
    wire signal_4926 ;
    wire signal_4927 ;
    wire signal_4928 ;
    wire signal_4929 ;
    wire signal_4930 ;
    wire signal_4931 ;
    wire signal_4932 ;
    wire signal_4933 ;
    wire signal_4934 ;
    wire signal_4935 ;
    wire signal_4936 ;
    wire signal_4937 ;
    wire signal_4938 ;
    wire signal_4939 ;
    wire signal_4940 ;
    wire signal_4941 ;
    wire signal_4942 ;
    wire signal_4943 ;
    wire signal_4944 ;
    wire signal_4945 ;
    wire signal_4946 ;
    wire signal_4947 ;
    wire signal_4948 ;
    wire signal_4949 ;
    wire signal_4950 ;
    wire signal_4951 ;
    wire signal_4952 ;
    wire signal_4953 ;
    wire signal_4954 ;
    wire signal_4955 ;
    wire signal_4956 ;
    wire signal_4957 ;
    wire signal_4958 ;
    wire signal_4959 ;
    wire signal_4960 ;
    wire signal_4961 ;
    wire signal_4962 ;
    wire signal_4963 ;
    wire signal_4964 ;
    wire signal_4965 ;
    wire signal_4966 ;
    wire signal_4967 ;
    wire signal_4968 ;
    wire signal_4969 ;
    wire signal_4970 ;
    wire signal_4971 ;
    wire signal_4972 ;
    wire signal_4973 ;
    wire signal_4974 ;
    wire signal_4975 ;
    wire signal_4976 ;
    wire signal_4977 ;
    wire signal_4978 ;
    wire signal_4979 ;
    wire signal_4980 ;
    wire signal_4981 ;
    wire signal_4982 ;
    wire signal_4983 ;
    wire signal_4984 ;
    wire signal_4985 ;
    wire signal_4986 ;
    wire signal_4987 ;
    wire signal_4988 ;
    wire signal_4989 ;
    wire signal_4990 ;
    wire signal_4991 ;
    wire signal_4992 ;
    wire signal_4993 ;
    wire signal_4994 ;
    wire signal_4995 ;
    wire signal_4996 ;
    wire signal_4997 ;
    wire signal_4998 ;
    wire signal_4999 ;
    wire signal_5000 ;
    wire signal_5001 ;
    wire signal_5002 ;
    wire signal_5003 ;
    wire signal_5004 ;
    wire signal_5005 ;
    wire signal_5006 ;
    wire signal_5007 ;
    wire signal_5008 ;
    wire signal_5009 ;
    wire signal_5010 ;
    wire signal_5011 ;
    wire signal_5012 ;
    wire signal_5013 ;
    wire signal_5014 ;
    wire signal_5015 ;
    wire signal_5016 ;
    wire signal_5017 ;
    wire signal_5018 ;
    wire signal_5019 ;
    wire signal_5020 ;
    wire signal_5021 ;
    wire signal_5022 ;
    wire signal_5023 ;
    wire signal_5024 ;
    wire signal_5025 ;
    wire signal_5026 ;
    wire signal_5027 ;
    wire signal_5028 ;
    wire signal_5029 ;
    wire signal_5030 ;
    wire signal_5031 ;
    wire signal_5032 ;
    wire signal_5033 ;
    wire signal_5034 ;
    wire signal_5035 ;
    wire signal_5036 ;
    wire signal_5037 ;
    wire signal_5038 ;
    wire signal_5039 ;
    wire signal_5040 ;
    wire signal_5041 ;
    wire signal_5042 ;
    wire signal_5043 ;
    wire signal_5044 ;
    wire signal_5045 ;
    wire signal_5046 ;
    wire signal_5047 ;
    wire signal_5048 ;
    wire signal_5049 ;
    wire signal_5050 ;
    wire signal_5051 ;
    wire signal_5052 ;
    wire signal_5053 ;
    wire signal_5054 ;
    wire signal_5055 ;
    wire signal_5056 ;
    wire signal_5057 ;
    wire signal_5058 ;
    wire signal_5059 ;
    wire signal_5060 ;
    wire signal_5061 ;
    wire signal_5062 ;
    wire signal_5063 ;
    wire signal_5064 ;
    wire signal_5065 ;
    wire signal_5066 ;
    wire signal_5067 ;
    wire signal_5068 ;
    wire signal_5069 ;
    wire signal_5070 ;
    wire signal_5071 ;
    wire signal_5072 ;
    wire signal_5073 ;
    wire signal_5074 ;
    wire signal_5075 ;
    wire signal_5076 ;
    wire signal_5077 ;
    wire signal_5078 ;
    wire signal_5079 ;
    wire signal_5080 ;
    wire signal_5081 ;
    wire signal_5082 ;
    wire signal_5083 ;
    wire signal_5084 ;
    wire signal_5085 ;
    wire signal_5086 ;
    wire signal_5087 ;
    wire signal_5088 ;
    wire signal_5089 ;
    wire signal_5090 ;
    wire signal_5091 ;
    wire signal_5092 ;
    wire signal_5093 ;
    wire signal_5094 ;
    wire signal_5095 ;
    wire signal_5096 ;
    wire signal_5097 ;
    wire signal_5098 ;
    wire signal_5099 ;
    wire signal_5100 ;
    wire signal_5101 ;
    wire signal_5102 ;
    wire signal_5103 ;
    wire signal_5104 ;
    wire signal_5105 ;
    wire signal_5106 ;
    wire signal_5107 ;
    wire signal_5108 ;
    wire signal_5109 ;
    wire signal_5110 ;
    wire signal_5111 ;
    wire signal_5112 ;
    wire signal_5113 ;
    wire signal_5114 ;
    wire signal_5115 ;
    wire signal_5116 ;
    wire signal_5117 ;
    wire signal_5118 ;
    wire signal_5119 ;
    wire signal_5120 ;
    wire signal_5121 ;
    wire signal_5122 ;
    wire signal_5123 ;
    wire signal_5124 ;
    wire signal_5125 ;
    wire signal_5126 ;
    wire signal_5127 ;
    wire signal_5128 ;
    wire signal_5129 ;
    wire signal_5130 ;
    wire signal_5131 ;
    wire signal_5132 ;
    wire signal_5133 ;
    wire signal_5134 ;
    wire signal_5135 ;
    wire signal_5136 ;
    wire signal_5137 ;
    wire signal_5138 ;
    wire signal_5139 ;
    wire signal_5140 ;
    wire signal_5141 ;
    wire signal_5142 ;
    wire signal_5143 ;
    wire signal_5144 ;
    wire signal_5145 ;
    wire signal_5146 ;
    wire signal_5147 ;
    wire signal_5148 ;
    wire signal_5149 ;
    wire signal_5150 ;
    wire signal_5151 ;
    wire signal_5152 ;
    wire signal_5153 ;
    wire signal_5154 ;
    wire signal_5155 ;
    wire signal_5156 ;
    wire signal_5157 ;
    wire signal_5158 ;
    wire signal_5159 ;
    wire signal_5160 ;
    wire signal_5161 ;
    wire signal_5162 ;
    wire signal_5163 ;
    wire signal_5164 ;
    wire signal_5165 ;
    wire signal_5166 ;
    wire signal_5167 ;
    wire signal_5168 ;
    wire signal_5169 ;
    wire signal_5170 ;
    wire signal_5171 ;
    wire signal_5172 ;
    wire signal_5173 ;
    wire signal_5174 ;
    wire signal_5175 ;
    wire signal_5176 ;
    wire signal_5177 ;
    wire signal_5178 ;
    wire signal_5179 ;
    wire signal_5180 ;
    wire signal_5181 ;
    wire signal_5182 ;
    wire signal_5183 ;
    wire signal_5184 ;
    wire signal_5185 ;
    wire signal_5186 ;
    wire signal_5187 ;
    wire signal_5188 ;
    wire signal_5189 ;
    wire signal_5190 ;
    wire signal_5191 ;
    wire signal_5192 ;
    wire signal_5193 ;
    wire signal_5194 ;
    wire signal_5195 ;
    wire signal_5196 ;
    wire signal_5197 ;
    wire signal_5198 ;
    wire signal_5199 ;
    wire signal_5200 ;
    wire signal_5201 ;
    wire signal_5202 ;
    wire signal_5203 ;
    wire signal_5204 ;
    wire signal_5205 ;
    wire signal_5206 ;
    wire signal_5207 ;
    wire signal_5208 ;
    wire signal_5209 ;
    wire signal_5210 ;
    wire signal_5211 ;
    wire signal_5212 ;
    wire signal_5213 ;
    wire signal_5214 ;
    wire signal_5215 ;
    wire signal_5216 ;
    wire signal_5217 ;
    wire signal_5218 ;
    wire signal_5219 ;
    wire signal_5220 ;
    wire signal_5221 ;
    wire signal_5222 ;
    wire signal_5223 ;
    wire signal_5224 ;
    wire signal_5225 ;
    wire signal_5226 ;
    wire signal_5227 ;
    wire signal_5228 ;
    wire signal_5229 ;
    wire signal_5230 ;
    wire signal_5231 ;
    wire signal_5232 ;
    wire signal_5233 ;
    wire signal_5234 ;
    wire signal_5235 ;
    wire signal_5236 ;
    wire signal_5237 ;
    wire signal_5238 ;
    wire signal_5239 ;
    wire signal_5240 ;
    wire signal_5241 ;
    wire signal_5242 ;
    wire signal_5243 ;
    wire signal_5244 ;
    wire signal_5245 ;
    wire signal_5246 ;
    wire signal_5247 ;
    wire signal_5248 ;
    wire signal_5249 ;
    wire signal_5250 ;
    wire signal_5251 ;
    wire signal_5252 ;
    wire signal_5253 ;
    wire signal_5254 ;
    wire signal_5255 ;
    wire signal_5256 ;
    wire signal_5257 ;
    wire signal_5258 ;
    wire signal_5259 ;
    wire signal_5260 ;
    wire signal_5261 ;
    wire signal_5262 ;
    wire signal_5263 ;
    wire signal_5264 ;
    wire signal_5265 ;
    wire signal_5266 ;
    wire signal_5267 ;
    wire signal_5268 ;
    wire signal_5269 ;
    wire signal_5270 ;
    wire signal_5271 ;
    wire signal_5272 ;
    wire signal_5273 ;
    wire signal_5274 ;
    wire signal_5275 ;
    wire signal_5276 ;
    wire signal_5277 ;
    wire signal_5278 ;
    wire signal_5279 ;
    wire signal_5280 ;
    wire signal_5281 ;
    wire signal_5282 ;
    wire signal_5283 ;
    wire signal_5284 ;
    wire signal_5285 ;
    wire signal_5286 ;
    wire signal_5287 ;
    wire signal_5288 ;
    wire signal_5289 ;
    wire signal_5290 ;
    wire signal_5291 ;
    wire signal_5292 ;
    wire signal_5293 ;
    wire signal_5294 ;
    wire signal_5295 ;
    wire signal_5296 ;
    wire signal_5297 ;
    wire signal_5298 ;
    wire signal_5299 ;
    wire signal_5300 ;
    wire signal_5301 ;
    wire signal_5302 ;
    wire signal_5303 ;
    wire signal_5304 ;
    wire signal_5305 ;
    wire signal_5306 ;
    wire signal_5307 ;
    wire signal_5308 ;
    wire signal_5309 ;
    wire signal_5310 ;
    wire signal_5311 ;
    wire signal_5312 ;
    wire signal_5313 ;
    wire signal_5314 ;
    wire signal_5315 ;
    wire signal_5316 ;
    wire signal_5317 ;
    wire signal_5318 ;
    wire signal_5319 ;
    wire signal_5320 ;
    wire signal_5321 ;
    wire signal_5322 ;
    wire signal_5323 ;
    wire signal_5324 ;
    wire signal_5325 ;
    wire signal_5326 ;
    wire signal_5327 ;
    wire signal_5328 ;
    wire signal_5329 ;
    wire signal_5330 ;
    wire signal_5331 ;
    wire signal_5332 ;
    wire signal_5333 ;
    wire signal_5334 ;
    wire signal_5335 ;
    wire signal_5336 ;
    wire signal_5337 ;
    wire signal_5338 ;
    wire signal_5339 ;
    wire signal_5340 ;
    wire signal_5341 ;
    wire signal_5342 ;
    wire signal_5343 ;
    wire signal_5344 ;
    wire signal_5345 ;
    wire signal_5346 ;
    wire signal_5347 ;
    wire signal_5348 ;
    wire signal_5349 ;
    wire signal_5350 ;
    wire signal_5351 ;
    wire signal_5352 ;
    wire signal_5353 ;
    wire signal_5354 ;
    wire signal_5355 ;
    wire signal_5356 ;
    wire signal_5357 ;
    wire signal_5358 ;
    wire signal_5359 ;
    wire signal_5360 ;
    wire signal_5361 ;
    wire signal_5362 ;
    wire signal_5363 ;
    wire signal_5364 ;
    wire signal_5365 ;
    wire signal_5366 ;
    wire signal_5367 ;
    wire signal_5368 ;
    wire signal_5369 ;
    wire signal_5370 ;
    wire signal_5371 ;
    wire signal_5372 ;
    wire signal_5373 ;
    wire signal_5374 ;
    wire signal_5375 ;
    wire signal_5376 ;
    wire signal_5377 ;
    wire signal_5378 ;
    wire signal_5379 ;
    wire signal_5380 ;
    wire signal_5381 ;
    wire signal_5382 ;
    wire signal_5383 ;
    wire signal_5384 ;
    wire signal_5385 ;
    wire signal_5386 ;
    wire signal_5387 ;
    wire signal_5388 ;
    wire signal_5389 ;
    wire signal_5390 ;
    wire signal_5391 ;
    wire signal_5392 ;
    wire signal_5393 ;
    wire signal_5394 ;
    wire signal_5395 ;
    wire signal_5396 ;
    wire signal_5397 ;
    wire signal_5398 ;
    wire signal_5399 ;
    wire signal_5400 ;
    wire signal_5401 ;
    wire signal_5402 ;
    wire signal_5403 ;
    wire signal_5404 ;
    wire signal_5405 ;
    wire signal_5406 ;
    wire signal_5407 ;
    wire signal_5408 ;
    wire signal_5409 ;
    wire signal_5410 ;
    wire signal_5411 ;
    wire signal_5412 ;
    wire signal_5413 ;
    wire signal_5414 ;
    wire signal_5415 ;
    wire signal_5416 ;
    wire signal_5417 ;
    wire signal_5418 ;
    wire signal_5419 ;
    wire signal_5420 ;
    wire signal_5421 ;
    wire signal_5422 ;
    wire signal_5423 ;
    wire signal_5424 ;
    wire signal_5425 ;
    wire signal_5426 ;
    wire signal_5427 ;
    wire signal_5428 ;
    wire signal_5429 ;
    wire signal_5430 ;
    wire signal_5431 ;
    wire signal_5432 ;
    wire signal_5433 ;
    wire signal_5434 ;
    wire signal_5435 ;
    wire signal_5436 ;
    wire signal_5437 ;
    wire signal_5438 ;
    wire signal_5439 ;
    wire signal_5440 ;
    wire signal_5441 ;
    wire signal_5442 ;
    wire signal_5443 ;
    wire signal_5444 ;
    wire signal_5445 ;
    wire signal_5446 ;
    wire signal_5447 ;
    wire signal_5448 ;
    wire signal_5449 ;
    wire signal_5450 ;
    wire signal_5451 ;
    wire signal_5452 ;
    wire signal_5453 ;
    wire signal_5454 ;
    wire signal_5455 ;
    wire signal_5456 ;
    wire signal_5457 ;
    wire signal_5458 ;
    wire signal_5459 ;
    wire signal_5460 ;
    wire signal_5461 ;
    wire signal_5462 ;
    wire signal_5463 ;
    wire signal_5464 ;
    wire signal_5465 ;
    wire signal_5466 ;
    wire signal_5467 ;
    wire signal_5468 ;
    wire signal_5469 ;
    wire signal_5470 ;
    wire signal_5471 ;
    wire signal_5472 ;
    wire signal_5473 ;
    wire signal_5474 ;
    wire signal_5475 ;
    wire signal_5476 ;
    wire signal_5477 ;
    wire signal_5478 ;
    wire signal_5479 ;
    wire signal_5480 ;
    wire signal_5481 ;
    wire signal_5482 ;
    wire signal_5483 ;
    wire signal_5484 ;
    wire signal_5485 ;
    wire signal_5486 ;
    wire signal_5487 ;
    wire signal_5488 ;
    wire signal_5489 ;
    wire signal_5490 ;
    wire signal_5491 ;
    wire signal_5492 ;
    wire signal_5493 ;
    wire signal_5494 ;
    wire signal_5495 ;
    wire signal_5496 ;
    wire signal_5497 ;
    wire signal_5498 ;
    wire signal_5499 ;
    wire signal_5500 ;
    wire signal_5501 ;
    wire signal_5502 ;
    wire signal_5503 ;
    wire signal_5504 ;
    wire signal_5505 ;
    wire signal_5506 ;
    wire signal_5507 ;
    wire signal_5508 ;
    wire signal_5509 ;
    wire signal_5510 ;
    wire signal_5511 ;
    wire signal_5512 ;
    wire signal_5513 ;
    wire signal_5514 ;
    wire signal_5515 ;
    wire signal_5516 ;
    wire signal_5517 ;
    wire signal_5518 ;
    wire signal_5519 ;
    wire signal_5520 ;
    wire signal_5521 ;
    wire signal_5522 ;
    wire signal_5523 ;
    wire signal_5524 ;
    wire signal_5525 ;
    wire signal_5526 ;
    wire signal_5527 ;
    wire signal_5528 ;
    wire signal_5529 ;
    wire signal_5530 ;
    wire signal_5531 ;
    wire signal_5532 ;
    wire signal_5533 ;
    wire signal_5534 ;
    wire signal_5535 ;
    wire signal_5536 ;
    wire signal_5537 ;
    wire signal_5538 ;
    wire signal_5539 ;
    wire signal_5540 ;
    wire signal_5541 ;
    wire signal_5542 ;
    wire signal_5543 ;
    wire signal_5544 ;
    wire signal_5545 ;
    wire signal_5546 ;
    wire signal_5547 ;
    wire signal_5548 ;
    wire signal_5549 ;
    wire signal_5550 ;
    wire signal_5551 ;
    wire signal_5552 ;
    wire signal_5553 ;
    wire signal_5554 ;
    wire signal_5555 ;
    wire signal_5556 ;
    wire signal_5557 ;
    wire signal_5558 ;
    wire signal_5559 ;
    wire signal_5560 ;
    wire signal_5561 ;
    wire signal_5562 ;
    wire signal_5563 ;
    wire signal_5564 ;
    wire signal_5565 ;
    wire signal_5566 ;
    wire signal_5567 ;
    wire signal_5568 ;
    wire signal_5569 ;
    wire signal_5570 ;
    wire signal_5571 ;
    wire signal_5572 ;
    wire signal_5573 ;
    wire signal_5574 ;
    wire signal_5575 ;
    wire signal_5576 ;
    wire signal_5577 ;
    wire signal_5578 ;
    wire signal_5579 ;
    wire signal_5580 ;
    wire signal_5581 ;
    wire signal_5582 ;
    wire signal_5583 ;
    wire signal_5584 ;
    wire signal_5585 ;
    wire signal_5586 ;
    wire signal_5587 ;
    wire signal_5588 ;
    wire signal_5589 ;
    wire signal_5590 ;
    wire signal_5591 ;
    wire signal_5592 ;
    wire signal_5593 ;
    wire signal_5594 ;
    wire signal_5595 ;
    wire signal_5596 ;
    wire signal_5597 ;
    wire signal_5598 ;
    wire signal_5599 ;
    wire signal_5600 ;
    wire signal_5601 ;
    wire signal_5602 ;
    wire signal_5603 ;
    wire signal_5604 ;
    wire signal_5605 ;
    wire signal_5606 ;
    wire signal_5607 ;
    wire signal_5608 ;
    wire signal_5609 ;
    wire signal_5610 ;
    wire signal_5611 ;
    wire signal_5612 ;
    wire signal_5613 ;
    wire signal_5614 ;
    wire signal_5615 ;
    wire signal_5616 ;
    wire signal_5617 ;
    wire signal_5618 ;
    wire signal_5619 ;
    wire signal_5620 ;
    wire signal_5621 ;
    wire signal_5622 ;
    wire signal_5623 ;
    wire signal_5624 ;
    wire signal_5625 ;
    wire signal_5626 ;
    wire signal_5627 ;
    wire signal_5628 ;
    wire signal_5629 ;
    wire signal_5630 ;
    wire signal_5631 ;
    wire signal_5632 ;
    wire signal_5633 ;
    wire signal_5634 ;
    wire signal_5635 ;
    wire signal_5636 ;
    wire signal_5637 ;
    wire signal_5638 ;
    wire signal_5639 ;
    wire signal_5640 ;
    wire signal_5641 ;
    wire signal_5642 ;
    wire signal_5643 ;
    wire signal_5644 ;
    wire signal_5645 ;
    wire signal_5646 ;
    wire signal_5647 ;
    wire signal_5648 ;
    wire signal_5649 ;
    wire signal_5650 ;
    wire signal_5651 ;
    wire signal_5652 ;
    wire signal_5653 ;
    wire signal_5654 ;
    wire signal_5655 ;
    wire signal_5656 ;
    wire signal_5657 ;
    wire signal_5658 ;
    wire signal_5659 ;
    wire signal_5660 ;
    wire signal_5661 ;
    wire signal_5662 ;
    wire signal_5663 ;
    wire signal_5664 ;
    wire signal_5665 ;
    wire signal_5666 ;
    wire signal_5667 ;
    wire signal_5668 ;
    wire signal_5669 ;
    wire signal_5670 ;
    wire signal_5671 ;
    wire signal_5672 ;
    wire signal_5673 ;
    wire signal_5674 ;
    wire signal_5675 ;
    wire signal_5676 ;
    wire signal_5677 ;
    wire signal_5678 ;
    wire signal_5679 ;
    wire signal_5680 ;
    wire signal_5681 ;
    wire signal_5682 ;
    wire signal_5683 ;
    wire signal_5684 ;
    wire signal_5685 ;
    wire signal_5686 ;
    wire signal_5687 ;
    wire signal_5688 ;
    wire signal_5689 ;
    wire signal_5690 ;
    wire signal_5691 ;
    wire signal_5692 ;
    wire signal_5693 ;
    wire signal_5694 ;
    wire signal_5695 ;
    wire signal_5696 ;
    wire signal_5697 ;
    wire signal_5698 ;
    wire signal_5699 ;
    wire signal_5700 ;
    wire signal_5701 ;
    wire signal_5702 ;
    wire signal_5703 ;
    wire signal_5704 ;
    wire signal_5705 ;
    wire signal_5706 ;
    wire signal_5707 ;
    wire signal_5708 ;
    wire signal_5709 ;
    wire signal_5710 ;
    wire signal_5711 ;
    wire signal_5712 ;
    wire signal_5713 ;
    wire signal_5714 ;
    wire signal_5715 ;
    wire signal_5716 ;
    wire signal_5717 ;
    wire signal_5718 ;
    wire signal_5719 ;
    wire signal_5720 ;
    wire signal_5721 ;
    wire signal_5722 ;
    wire signal_5723 ;
    wire signal_5724 ;
    wire signal_5725 ;
    wire signal_5726 ;
    wire signal_5727 ;
    wire signal_5728 ;
    wire signal_5729 ;
    wire signal_5730 ;
    wire signal_5731 ;
    wire signal_5732 ;
    wire signal_5733 ;
    wire signal_5734 ;
    wire signal_5735 ;
    wire signal_5736 ;
    wire signal_5737 ;
    wire signal_5738 ;
    wire signal_5739 ;
    wire signal_5740 ;
    wire signal_5741 ;
    wire signal_5742 ;
    wire signal_5743 ;
    wire signal_5744 ;
    wire signal_5745 ;
    wire signal_5746 ;
    wire signal_5747 ;
    wire signal_5748 ;
    wire signal_5749 ;
    wire signal_5750 ;
    wire signal_5751 ;
    wire signal_5752 ;
    wire signal_5753 ;
    wire signal_5754 ;
    wire signal_5755 ;
    wire signal_5756 ;
    wire signal_5757 ;
    wire signal_5758 ;
    wire signal_5759 ;
    wire signal_5760 ;
    wire signal_5761 ;
    wire signal_5762 ;
    wire signal_5763 ;
    wire signal_5764 ;
    wire signal_5765 ;
    wire signal_5766 ;
    wire signal_5767 ;
    wire signal_5768 ;
    wire signal_5769 ;
    wire signal_5770 ;
    wire signal_5771 ;
    wire signal_5772 ;
    wire signal_5773 ;
    wire signal_5774 ;
    wire signal_5775 ;
    wire signal_5776 ;
    wire signal_5777 ;
    wire signal_5778 ;
    wire signal_5779 ;
    wire signal_5780 ;
    wire signal_5781 ;
    wire signal_5782 ;
    wire signal_5783 ;
    wire signal_5784 ;
    wire signal_5785 ;
    wire signal_5786 ;
    wire signal_5787 ;
    wire signal_5788 ;
    wire signal_5789 ;
    wire signal_5790 ;
    wire signal_5791 ;
    wire signal_5792 ;
    wire signal_5793 ;
    wire signal_5794 ;
    wire signal_5795 ;
    wire signal_5796 ;
    wire signal_5797 ;
    wire signal_5798 ;
    wire signal_5799 ;
    wire signal_5800 ;
    wire signal_5801 ;
    wire signal_5802 ;
    wire signal_5803 ;
    wire signal_5804 ;
    wire signal_5805 ;
    wire signal_5806 ;
    wire signal_5807 ;
    wire signal_5808 ;
    wire signal_5809 ;
    wire signal_5810 ;
    wire signal_5811 ;
    wire signal_5812 ;
    wire signal_5813 ;
    wire signal_5814 ;
    wire signal_5815 ;
    wire signal_5816 ;
    wire signal_5817 ;
    wire signal_5818 ;
    wire signal_5819 ;
    wire signal_5820 ;
    wire signal_5821 ;
    wire signal_5822 ;
    wire signal_5823 ;
    wire signal_5824 ;
    wire signal_5825 ;
    wire signal_5826 ;
    wire signal_5827 ;
    wire signal_5828 ;
    wire signal_5829 ;
    wire signal_5830 ;
    wire signal_5831 ;
    wire signal_5832 ;
    wire signal_5833 ;
    wire signal_5834 ;
    wire signal_5835 ;
    wire signal_5836 ;
    wire signal_5837 ;
    wire signal_5838 ;
    wire signal_5839 ;
    wire signal_5840 ;
    wire signal_5841 ;
    wire signal_5842 ;
    wire signal_5843 ;
    wire signal_5844 ;
    wire signal_5845 ;
    wire signal_5846 ;
    wire signal_5847 ;
    wire signal_5848 ;
    wire signal_5849 ;
    wire signal_5850 ;
    wire signal_5851 ;
    wire signal_5852 ;
    wire signal_5853 ;
    wire signal_5854 ;
    wire signal_5855 ;
    wire signal_5856 ;
    wire signal_5857 ;
    wire signal_5858 ;
    wire signal_5859 ;
    wire signal_5860 ;
    wire signal_5861 ;
    wire signal_5862 ;
    wire signal_5863 ;
    wire signal_5864 ;
    wire signal_5865 ;
    wire signal_5866 ;
    wire signal_5867 ;
    wire signal_5868 ;
    wire signal_5869 ;
    wire signal_5870 ;
    wire signal_5871 ;
    wire signal_5872 ;
    wire signal_5873 ;
    wire signal_5874 ;
    wire signal_5875 ;
    wire signal_5876 ;
    wire signal_5877 ;
    wire signal_5878 ;
    wire signal_5879 ;
    wire signal_5880 ;
    wire signal_5881 ;
    wire signal_5882 ;
    wire signal_5883 ;
    wire signal_5884 ;
    wire signal_5885 ;
    wire signal_5886 ;
    wire signal_5887 ;
    wire signal_5888 ;
    wire signal_5889 ;
    wire signal_5890 ;
    wire signal_5891 ;
    wire signal_5892 ;
    wire signal_5893 ;
    wire signal_5894 ;
    wire signal_5895 ;
    wire signal_5896 ;
    wire signal_5897 ;
    wire signal_5898 ;
    wire signal_5899 ;
    wire signal_5900 ;
    wire signal_5901 ;
    wire signal_5902 ;
    wire signal_5903 ;
    wire signal_5904 ;
    wire signal_5905 ;
    wire signal_5906 ;
    wire signal_5907 ;
    wire signal_5908 ;
    wire signal_5909 ;
    wire signal_5910 ;
    wire signal_5911 ;
    wire signal_5912 ;
    wire signal_5913 ;
    wire signal_5914 ;
    wire signal_5915 ;
    wire signal_5916 ;
    wire signal_5917 ;
    wire signal_5918 ;
    wire signal_5919 ;
    wire signal_5920 ;
    wire signal_5921 ;
    wire signal_5922 ;
    wire signal_5923 ;
    wire signal_5924 ;
    wire signal_5925 ;
    wire signal_5926 ;
    wire signal_5927 ;
    wire signal_5928 ;
    wire signal_5929 ;
    wire signal_5930 ;
    wire signal_5931 ;
    wire signal_5932 ;
    wire signal_5933 ;
    wire signal_5934 ;
    wire signal_5935 ;
    wire signal_5936 ;
    wire signal_5937 ;
    wire signal_5938 ;
    wire signal_5939 ;
    wire signal_5940 ;
    wire signal_5941 ;
    wire signal_5942 ;
    wire signal_5943 ;
    wire signal_5944 ;
    wire signal_5945 ;
    wire signal_5946 ;
    wire signal_5947 ;
    wire signal_5948 ;
    wire signal_5949 ;
    wire signal_5950 ;
    wire signal_5951 ;
    wire signal_5952 ;
    wire signal_5953 ;
    wire signal_5954 ;
    wire signal_5955 ;
    wire signal_5956 ;
    wire signal_5957 ;
    wire signal_5958 ;
    wire signal_5959 ;
    wire signal_5960 ;
    wire signal_5961 ;
    wire signal_5962 ;
    wire signal_5963 ;
    wire signal_5964 ;
    wire signal_5965 ;
    wire signal_5966 ;
    wire signal_5967 ;
    wire signal_5968 ;
    wire signal_5969 ;
    wire signal_5970 ;
    wire signal_5971 ;
    wire signal_5972 ;
    wire signal_5973 ;
    wire signal_5974 ;
    wire signal_5975 ;
    wire signal_5976 ;
    wire signal_5977 ;
    wire signal_5978 ;
    wire signal_5979 ;
    wire signal_5980 ;
    wire signal_5981 ;
    wire signal_5982 ;
    wire signal_5983 ;
    wire signal_5984 ;
    wire signal_5985 ;
    wire signal_5986 ;
    wire signal_5987 ;
    wire signal_5988 ;
    wire signal_5989 ;
    wire signal_5990 ;
    wire signal_5991 ;
    wire signal_5992 ;
    wire signal_5993 ;
    wire signal_5994 ;
    wire signal_5995 ;
    wire signal_5996 ;
    wire signal_5997 ;
    wire signal_5998 ;
    wire signal_5999 ;
    wire signal_6000 ;
    wire signal_6001 ;
    wire signal_6002 ;
    wire signal_6003 ;
    wire signal_6004 ;
    wire signal_6005 ;
    wire signal_6006 ;
    wire signal_6007 ;
    wire signal_6008 ;
    wire signal_6009 ;
    wire signal_6010 ;
    wire signal_6011 ;
    wire signal_6012 ;
    wire signal_6013 ;
    wire signal_6014 ;
    wire signal_6015 ;
    wire signal_6016 ;
    wire signal_6017 ;
    wire signal_6018 ;
    wire signal_6019 ;
    wire signal_6020 ;
    wire signal_6021 ;
    wire signal_6022 ;
    wire signal_6023 ;
    wire signal_6024 ;
    wire signal_6025 ;
    wire signal_6026 ;
    wire signal_6027 ;
    wire signal_6028 ;
    wire signal_6029 ;
    wire signal_6030 ;
    wire signal_6031 ;
    wire signal_6032 ;
    wire signal_6033 ;
    wire signal_6034 ;
    wire signal_6035 ;
    wire signal_6036 ;
    wire signal_6037 ;
    wire signal_6038 ;
    wire signal_6039 ;
    wire signal_6040 ;
    wire signal_6041 ;
    wire signal_6042 ;
    wire signal_6043 ;
    wire signal_6044 ;
    wire signal_6045 ;
    wire signal_6046 ;
    wire signal_6047 ;
    wire signal_6048 ;
    wire signal_6049 ;
    wire signal_6050 ;
    wire signal_6051 ;
    wire signal_6052 ;
    wire signal_6053 ;
    wire signal_6054 ;
    wire signal_6055 ;
    wire signal_6056 ;
    wire signal_6057 ;
    wire signal_6058 ;
    wire signal_6059 ;
    wire signal_6060 ;
    wire signal_6061 ;
    wire signal_6062 ;
    wire signal_6063 ;
    wire signal_6064 ;
    wire signal_6065 ;
    wire signal_6066 ;
    wire signal_6067 ;
    wire signal_6068 ;
    wire signal_6069 ;
    wire signal_6070 ;
    wire signal_6071 ;
    wire signal_6072 ;
    wire signal_6073 ;
    wire signal_6074 ;
    wire signal_6075 ;
    wire signal_6076 ;
    wire signal_6077 ;
    wire signal_6078 ;
    wire signal_6079 ;
    wire signal_6080 ;
    wire signal_6081 ;
    wire signal_6082 ;
    wire signal_6083 ;
    wire signal_6084 ;
    wire signal_6085 ;
    wire signal_6086 ;
    wire signal_6087 ;
    wire signal_6088 ;
    wire signal_6089 ;
    wire signal_6090 ;
    wire signal_6091 ;
    wire signal_6092 ;
    wire signal_6093 ;
    wire signal_6094 ;
    wire signal_6095 ;
    wire signal_6096 ;
    wire signal_6097 ;
    wire signal_6098 ;
    wire signal_6099 ;
    wire signal_6100 ;
    wire signal_6101 ;
    wire signal_6102 ;
    wire signal_6103 ;
    wire signal_6104 ;
    wire signal_6105 ;
    wire signal_6106 ;
    wire signal_6107 ;
    wire signal_6108 ;
    wire signal_6109 ;
    wire signal_6110 ;
    wire signal_6111 ;
    wire signal_6112 ;
    wire signal_6113 ;
    wire signal_6114 ;
    wire signal_6115 ;
    wire signal_6116 ;
    wire signal_6117 ;
    wire signal_6118 ;
    wire signal_6119 ;
    wire signal_6120 ;
    wire signal_6121 ;
    wire signal_6122 ;
    wire signal_6123 ;
    wire signal_6124 ;
    wire signal_6125 ;
    wire signal_6126 ;
    wire signal_6127 ;
    wire signal_6128 ;
    wire signal_6129 ;
    wire signal_6130 ;
    wire signal_6131 ;
    wire signal_6132 ;
    wire signal_6133 ;
    wire signal_6134 ;
    wire signal_6135 ;
    wire signal_6136 ;
    wire signal_6137 ;
    wire signal_6138 ;
    wire signal_6139 ;
    wire signal_6140 ;
    wire signal_6141 ;
    wire signal_6142 ;
    wire signal_6143 ;
    wire signal_6144 ;
    wire signal_6145 ;
    wire signal_6146 ;
    wire signal_6147 ;
    wire signal_6148 ;
    wire signal_6149 ;
    wire signal_6150 ;
    wire signal_6151 ;
    wire signal_6152 ;
    wire signal_6153 ;
    wire signal_6154 ;
    wire signal_6155 ;
    wire signal_6156 ;
    wire signal_6157 ;
    wire signal_6158 ;
    wire signal_6159 ;
    wire signal_6160 ;
    wire signal_6161 ;
    wire signal_6162 ;
    wire signal_6163 ;
    wire signal_6164 ;
    wire signal_6165 ;
    wire signal_6166 ;
    wire signal_6167 ;
    wire signal_6168 ;
    wire signal_6169 ;
    wire signal_6170 ;
    wire signal_6171 ;
    wire signal_6172 ;
    wire signal_6173 ;
    wire signal_6174 ;
    wire signal_6175 ;
    wire signal_6176 ;
    wire signal_6177 ;
    wire signal_6178 ;
    wire signal_6179 ;
    wire signal_6180 ;
    wire signal_6181 ;
    wire signal_6182 ;
    wire signal_6183 ;
    wire signal_6184 ;
    wire signal_6185 ;
    wire signal_6186 ;
    wire signal_6187 ;
    wire signal_6188 ;
    wire signal_6189 ;
    wire signal_6190 ;
    wire signal_6191 ;
    wire signal_6192 ;
    wire signal_6193 ;
    wire signal_6194 ;
    wire signal_6195 ;
    wire signal_6196 ;
    wire signal_6197 ;
    wire signal_6198 ;
    wire signal_6199 ;
    wire signal_6200 ;
    wire signal_6201 ;
    wire signal_6202 ;
    wire signal_6203 ;
    wire signal_6204 ;
    wire signal_6205 ;
    wire signal_6206 ;
    wire signal_6207 ;
    wire signal_6208 ;
    wire signal_6209 ;
    wire signal_6210 ;
    wire signal_6211 ;
    wire signal_6212 ;
    wire signal_6213 ;
    wire signal_6214 ;
    wire signal_6215 ;
    wire signal_6216 ;
    wire signal_6217 ;
    wire signal_6218 ;
    wire signal_6219 ;
    wire signal_6220 ;
    wire signal_6221 ;
    wire signal_6222 ;
    wire signal_6223 ;
    wire signal_6224 ;
    wire signal_6225 ;
    wire signal_6226 ;
    wire signal_6227 ;
    wire signal_6228 ;
    wire signal_6229 ;
    wire signal_6230 ;
    wire signal_6231 ;
    wire signal_6232 ;
    wire signal_6233 ;
    wire signal_6234 ;
    wire signal_6235 ;
    wire signal_6236 ;
    wire signal_6237 ;
    wire signal_6238 ;
    wire signal_6239 ;
    wire signal_6240 ;
    wire signal_6241 ;
    wire signal_6242 ;
    wire signal_6243 ;
    wire signal_6244 ;
    wire signal_6245 ;
    wire signal_6246 ;
    wire signal_6247 ;
    wire signal_6248 ;
    wire signal_6249 ;
    wire signal_6250 ;
    wire signal_6251 ;
    wire signal_6252 ;
    wire signal_6253 ;
    wire signal_6254 ;
    wire signal_6255 ;
    wire signal_6256 ;
    wire signal_6257 ;
    wire signal_6258 ;
    wire signal_6259 ;
    wire signal_6260 ;
    wire signal_6261 ;
    wire signal_6262 ;
    wire signal_6263 ;
    wire signal_6264 ;
    wire signal_6265 ;
    wire signal_6266 ;
    wire signal_6267 ;
    wire signal_6268 ;
    wire signal_6269 ;
    wire signal_6270 ;
    wire signal_6271 ;
    wire signal_6272 ;
    wire signal_6273 ;
    wire signal_6274 ;
    wire signal_6275 ;
    wire signal_6276 ;
    wire signal_6277 ;
    wire signal_6278 ;
    wire signal_6279 ;
    wire signal_6280 ;
    wire signal_6281 ;
    wire signal_6282 ;
    wire signal_6283 ;
    wire signal_6284 ;
    wire signal_6285 ;
    wire signal_6286 ;
    wire signal_6287 ;
    wire signal_6288 ;
    wire signal_6289 ;
    wire signal_6290 ;
    wire signal_6291 ;
    wire signal_6292 ;
    wire signal_6293 ;
    wire signal_6294 ;
    wire signal_6295 ;
    wire signal_6296 ;
    wire signal_6297 ;
    wire signal_6298 ;
    wire signal_6299 ;
    wire signal_6300 ;
    wire signal_6301 ;
    wire signal_6302 ;
    wire signal_6303 ;
    wire signal_6304 ;
    wire signal_6305 ;
    wire signal_6306 ;
    wire signal_6307 ;
    wire signal_6308 ;
    wire signal_6309 ;
    wire signal_6310 ;
    wire signal_6311 ;
    wire signal_6312 ;
    wire signal_6313 ;
    wire signal_6314 ;
    wire signal_6315 ;
    wire signal_6316 ;
    wire signal_6317 ;
    wire signal_6318 ;
    wire signal_6319 ;
    wire signal_6320 ;
    wire signal_6321 ;
    wire signal_6322 ;
    wire signal_6323 ;
    wire signal_6324 ;
    wire signal_6325 ;
    wire signal_6326 ;
    wire signal_6327 ;
    wire signal_6328 ;
    wire signal_6329 ;
    wire signal_6330 ;
    wire signal_6331 ;
    wire signal_6332 ;
    wire signal_6333 ;
    wire signal_6334 ;
    wire signal_6335 ;
    wire signal_6336 ;
    wire signal_6337 ;
    wire signal_6338 ;
    wire signal_6339 ;
    wire signal_6340 ;
    wire signal_6341 ;
    wire signal_6342 ;
    wire signal_6343 ;
    wire signal_6344 ;
    wire signal_6345 ;
    wire signal_6346 ;
    wire signal_6347 ;
    wire signal_6348 ;
    wire signal_6349 ;
    wire signal_6350 ;
    wire signal_6351 ;
    wire signal_6352 ;
    wire signal_6353 ;
    wire signal_6354 ;
    wire signal_6355 ;
    wire signal_6356 ;
    wire signal_6357 ;
    wire signal_6358 ;
    wire signal_6359 ;
    wire signal_6360 ;
    wire signal_6361 ;
    wire signal_6362 ;
    wire signal_6363 ;
    wire signal_6364 ;
    wire signal_6365 ;
    wire signal_6366 ;
    wire signal_6367 ;
    wire signal_6368 ;
    wire signal_6369 ;
    wire signal_6370 ;
    wire signal_6371 ;
    wire signal_6372 ;
    wire signal_6373 ;
    wire signal_6374 ;
    wire signal_6375 ;
    wire signal_6376 ;
    wire signal_6377 ;
    wire signal_6378 ;
    wire signal_6379 ;
    wire signal_6380 ;
    wire signal_6381 ;
    wire signal_6382 ;
    wire signal_6383 ;
    wire signal_6384 ;
    wire signal_6385 ;
    wire signal_6386 ;
    wire signal_6387 ;
    wire signal_6388 ;
    wire signal_6389 ;
    wire signal_6390 ;
    wire signal_6391 ;
    wire signal_6392 ;
    wire signal_6393 ;
    wire signal_6394 ;
    wire signal_6395 ;
    wire signal_6396 ;
    wire signal_6397 ;
    wire signal_6398 ;
    wire signal_6399 ;
    wire signal_6400 ;
    wire signal_6401 ;
    wire signal_6402 ;
    wire signal_6403 ;
    wire signal_6404 ;
    wire signal_6405 ;
    wire signal_6406 ;
    wire signal_6407 ;
    wire signal_6408 ;
    wire signal_6409 ;
    wire signal_6410 ;
    wire signal_6411 ;
    wire signal_6412 ;
    wire signal_6413 ;
    wire signal_6414 ;
    wire signal_6415 ;
    wire signal_6416 ;
    wire signal_6417 ;
    wire signal_6418 ;
    wire signal_6419 ;
    wire signal_6420 ;
    wire signal_6421 ;
    wire signal_6422 ;
    wire signal_6423 ;
    wire signal_6424 ;
    wire signal_6425 ;
    wire signal_6426 ;
    wire signal_6427 ;
    wire signal_6428 ;
    wire signal_6429 ;
    wire signal_6430 ;
    wire signal_6431 ;
    wire signal_6432 ;
    wire signal_6433 ;
    wire signal_6434 ;
    wire signal_6435 ;
    wire signal_6436 ;
    wire signal_6437 ;
    wire signal_6438 ;
    wire signal_6439 ;
    wire signal_6440 ;
    wire signal_6441 ;
    wire signal_6442 ;
    wire signal_6443 ;
    wire signal_6444 ;
    wire signal_6445 ;
    wire signal_6446 ;
    wire signal_6447 ;
    wire signal_6448 ;
    wire signal_6449 ;
    wire signal_6450 ;
    wire signal_6451 ;
    wire signal_6452 ;
    wire signal_6453 ;
    wire signal_6454 ;
    wire signal_6455 ;
    wire signal_6456 ;
    wire signal_6457 ;
    wire signal_6458 ;
    wire signal_6459 ;
    wire signal_6460 ;
    wire signal_6461 ;
    wire signal_6462 ;
    wire signal_6463 ;
    wire signal_6464 ;
    wire signal_6465 ;
    wire signal_6466 ;
    wire signal_6467 ;
    wire signal_6468 ;
    wire signal_6469 ;
    wire signal_6470 ;
    wire signal_6471 ;
    wire signal_6472 ;
    wire signal_6473 ;
    wire signal_6474 ;
    wire signal_6475 ;
    wire signal_6476 ;
    wire signal_6477 ;
    wire signal_6478 ;
    wire signal_6479 ;
    wire signal_6480 ;
    wire signal_6481 ;
    wire signal_6482 ;
    wire signal_6483 ;
    wire signal_6484 ;
    wire signal_6485 ;
    wire signal_6486 ;
    wire signal_6487 ;
    wire signal_6488 ;
    wire signal_6489 ;
    wire signal_6490 ;
    wire signal_6491 ;
    wire signal_6492 ;
    wire signal_6493 ;
    wire signal_6494 ;
    wire signal_6495 ;
    wire signal_6496 ;
    wire signal_6497 ;
    wire signal_6498 ;
    wire signal_6499 ;
    wire signal_6500 ;
    wire signal_6501 ;
    wire signal_6502 ;
    wire signal_6503 ;
    wire signal_6504 ;
    wire signal_6505 ;
    wire signal_6506 ;
    wire signal_6507 ;
    wire signal_6508 ;
    wire signal_6509 ;
    wire signal_6510 ;
    wire signal_6511 ;
    wire signal_6512 ;
    wire signal_6513 ;
    wire signal_6514 ;
    wire signal_6515 ;
    wire signal_6516 ;
    wire signal_6517 ;
    wire signal_6518 ;
    wire signal_6519 ;
    wire signal_6520 ;
    wire signal_6521 ;
    wire signal_6522 ;
    wire signal_6523 ;
    wire signal_6524 ;
    wire signal_6525 ;
    wire signal_6526 ;
    wire signal_6527 ;
    wire signal_6528 ;
    wire signal_6529 ;
    wire signal_6530 ;
    wire signal_6531 ;
    wire signal_6532 ;
    wire signal_6533 ;
    wire signal_6534 ;
    wire signal_6535 ;
    wire signal_6536 ;
    wire signal_6537 ;
    wire signal_6538 ;
    wire signal_6539 ;
    wire signal_6540 ;
    wire signal_6541 ;
    wire signal_6542 ;
    wire signal_6543 ;
    wire signal_6544 ;
    wire signal_6545 ;
    wire signal_6546 ;
    wire signal_6547 ;
    wire signal_6548 ;
    wire signal_6549 ;
    wire signal_6550 ;
    wire signal_6551 ;
    wire signal_6552 ;
    wire signal_6553 ;
    wire signal_6554 ;
    wire signal_6555 ;
    wire signal_6556 ;
    wire signal_6557 ;
    wire signal_6558 ;
    wire signal_6559 ;
    wire signal_6560 ;
    wire signal_6561 ;
    wire signal_6562 ;
    wire signal_6563 ;
    wire signal_6564 ;
    wire signal_6565 ;
    wire signal_6566 ;
    wire signal_6567 ;
    wire signal_6568 ;
    wire signal_6569 ;
    wire signal_6570 ;
    wire signal_6571 ;
    wire signal_6572 ;
    wire signal_6573 ;
    wire signal_6574 ;
    wire signal_6575 ;
    wire signal_6576 ;
    wire signal_6577 ;
    wire signal_6578 ;
    wire signal_6579 ;
    wire signal_6580 ;
    wire signal_6581 ;
    wire signal_6582 ;
    wire signal_6583 ;
    wire signal_6584 ;
    wire signal_6585 ;
    wire signal_6586 ;
    wire signal_6587 ;
    wire signal_6588 ;
    wire signal_6589 ;
    wire signal_6590 ;
    wire signal_6591 ;
    wire signal_6592 ;
    wire signal_6593 ;
    wire signal_6594 ;
    wire signal_6595 ;
    wire signal_6596 ;
    wire signal_6597 ;
    wire signal_6598 ;
    wire signal_6599 ;
    wire signal_6600 ;
    wire signal_6601 ;
    wire signal_6602 ;
    wire signal_6603 ;
    wire signal_6604 ;
    wire signal_6605 ;
    wire signal_6606 ;
    wire signal_6607 ;
    wire signal_6608 ;
    wire signal_6609 ;
    wire signal_6610 ;
    wire signal_6611 ;
    wire signal_6612 ;
    wire signal_6613 ;
    wire signal_6614 ;
    wire signal_6615 ;
    wire signal_6616 ;
    wire signal_6617 ;
    wire signal_6618 ;
    wire signal_6619 ;
    wire signal_6620 ;
    wire signal_6621 ;
    wire signal_6622 ;
    wire signal_6623 ;
    wire signal_6624 ;
    wire signal_6625 ;
    wire signal_6626 ;
    wire signal_6627 ;
    wire signal_6628 ;
    wire signal_6629 ;
    wire signal_6630 ;
    wire signal_6631 ;
    wire signal_6632 ;
    wire signal_6633 ;
    wire signal_6634 ;
    wire signal_6635 ;
    wire signal_6636 ;
    wire signal_6637 ;
    wire signal_6638 ;
    wire signal_6639 ;
    wire signal_6640 ;
    wire signal_6641 ;
    wire signal_6642 ;
    wire signal_6643 ;
    wire signal_6644 ;
    wire signal_6645 ;
    wire signal_6646 ;
    wire signal_6647 ;
    wire signal_6648 ;
    wire signal_6649 ;
    wire signal_6650 ;
    wire signal_6651 ;
    wire signal_6652 ;
    wire signal_6653 ;
    wire signal_6654 ;
    wire signal_6655 ;
    wire signal_6656 ;
    wire signal_6657 ;
    wire signal_6658 ;
    wire signal_6659 ;
    wire signal_6660 ;
    wire signal_6661 ;
    wire signal_6662 ;
    wire signal_6663 ;
    wire signal_6664 ;
    wire signal_6665 ;
    wire signal_6666 ;
    wire signal_6667 ;
    wire signal_6668 ;
    wire signal_6669 ;
    wire signal_6670 ;
    wire signal_6671 ;
    wire signal_6672 ;
    wire signal_6673 ;
    wire signal_6674 ;
    wire signal_6675 ;
    wire signal_6676 ;
    wire signal_6677 ;
    wire signal_6678 ;
    wire signal_6679 ;
    wire signal_6680 ;
    wire signal_6681 ;
    wire signal_6682 ;
    wire signal_6683 ;
    wire signal_6684 ;
    wire signal_6685 ;
    wire signal_6686 ;
    wire signal_6687 ;
    wire signal_6688 ;
    wire signal_6689 ;
    wire signal_6690 ;
    wire signal_6691 ;
    wire signal_6692 ;
    wire signal_6693 ;
    wire signal_6694 ;
    wire signal_6695 ;
    wire signal_6696 ;
    wire signal_6697 ;
    wire signal_6698 ;
    wire signal_6699 ;
    wire signal_6700 ;
    wire signal_6701 ;
    wire signal_6702 ;
    wire signal_6703 ;
    wire signal_6704 ;
    wire signal_6705 ;
    wire signal_6706 ;
    wire signal_6707 ;
    wire signal_6708 ;
    wire signal_6709 ;
    wire signal_6710 ;
    wire signal_6711 ;
    wire signal_6712 ;
    wire signal_6713 ;
    wire signal_6714 ;
    wire signal_6715 ;
    wire signal_6716 ;
    wire signal_6717 ;
    wire signal_6718 ;
    wire signal_6719 ;
    wire signal_6720 ;
    wire signal_6721 ;
    wire signal_6722 ;
    wire signal_6723 ;
    wire signal_6724 ;
    wire signal_6725 ;
    wire signal_6726 ;
    wire signal_6727 ;
    wire signal_6728 ;
    wire signal_6729 ;
    wire signal_6730 ;
    wire signal_6731 ;
    wire signal_6732 ;
    wire signal_6733 ;
    wire signal_6734 ;
    wire signal_6735 ;
    wire signal_6736 ;
    wire signal_6737 ;
    wire signal_6738 ;
    wire signal_6739 ;
    wire signal_6740 ;
    wire signal_6741 ;
    wire signal_6742 ;
    wire signal_6743 ;
    wire signal_6744 ;
    wire signal_6745 ;
    wire signal_6746 ;
    wire signal_6747 ;
    wire signal_6748 ;
    wire signal_6749 ;
    wire signal_6750 ;
    wire signal_6751 ;
    wire signal_6752 ;
    wire signal_6753 ;
    wire signal_6754 ;
    wire signal_6755 ;
    wire signal_6756 ;
    wire signal_6757 ;
    wire signal_6758 ;
    wire signal_6759 ;
    wire signal_6760 ;
    wire signal_6761 ;
    wire signal_6762 ;
    wire signal_6763 ;
    wire signal_6764 ;
    wire signal_6765 ;
    wire signal_6766 ;
    wire signal_6767 ;
    wire signal_6768 ;
    wire signal_6769 ;
    wire signal_6770 ;
    wire signal_6771 ;
    wire signal_6772 ;
    wire signal_6773 ;
    wire signal_6774 ;
    wire signal_6775 ;
    wire signal_6776 ;
    wire signal_6777 ;
    wire signal_6778 ;
    wire signal_6779 ;
    wire signal_6780 ;
    wire signal_6781 ;
    wire signal_6782 ;
    wire signal_6783 ;
    wire signal_6784 ;
    wire signal_6785 ;
    wire signal_6786 ;
    wire signal_6787 ;
    wire signal_6788 ;
    wire signal_6789 ;
    wire signal_6790 ;
    wire signal_6791 ;
    wire signal_6792 ;
    wire signal_6793 ;
    wire signal_6794 ;
    wire signal_6795 ;
    wire signal_6796 ;
    wire signal_6797 ;
    wire signal_6798 ;
    wire signal_6799 ;
    wire signal_6800 ;
    wire signal_6801 ;
    wire signal_6802 ;
    wire signal_6803 ;
    wire signal_6804 ;
    wire signal_6805 ;
    wire signal_6806 ;
    wire signal_6807 ;
    wire signal_6808 ;
    wire signal_6809 ;
    wire signal_6810 ;
    wire signal_6811 ;
    wire signal_6812 ;
    wire signal_6813 ;
    wire signal_6814 ;
    wire signal_6815 ;
    wire signal_6816 ;
    wire signal_6817 ;
    wire signal_6818 ;
    wire signal_6819 ;
    wire signal_6820 ;
    wire signal_6821 ;
    wire signal_6822 ;
    wire signal_6823 ;
    wire signal_6824 ;
    wire signal_6825 ;
    wire signal_6826 ;
    wire signal_6827 ;
    wire signal_6828 ;
    wire signal_6829 ;
    wire signal_6830 ;
    wire signal_6831 ;
    wire signal_6832 ;
    wire signal_6833 ;
    wire signal_6834 ;
    wire signal_6835 ;
    wire signal_6836 ;
    wire signal_6837 ;
    wire signal_6838 ;
    wire signal_6839 ;
    wire signal_6840 ;
    wire signal_6841 ;
    wire signal_6842 ;
    wire signal_6843 ;
    wire signal_6844 ;
    wire signal_6845 ;
    wire signal_6846 ;
    wire signal_6847 ;
    wire signal_6848 ;
    wire signal_6849 ;
    wire signal_6850 ;
    wire signal_6851 ;
    wire signal_6852 ;
    wire signal_6853 ;
    wire signal_6854 ;
    wire signal_6855 ;
    wire signal_6856 ;
    wire signal_6857 ;
    wire signal_6858 ;
    wire signal_6859 ;
    wire signal_6860 ;
    wire signal_6861 ;
    wire signal_6862 ;
    wire signal_6863 ;
    wire signal_6864 ;
    wire signal_6865 ;
    wire signal_6866 ;
    wire signal_6867 ;
    wire signal_6868 ;
    wire signal_6869 ;
    wire signal_6870 ;
    wire signal_6871 ;
    wire signal_6872 ;
    wire signal_6873 ;
    wire signal_6874 ;
    wire signal_6875 ;
    wire signal_6876 ;
    wire signal_6877 ;
    wire signal_6878 ;
    wire signal_6879 ;
    wire signal_6880 ;
    wire signal_6881 ;
    wire signal_6882 ;
    wire signal_6883 ;
    wire signal_6884 ;
    wire signal_6885 ;
    wire signal_6886 ;
    wire signal_6887 ;
    wire signal_6888 ;
    wire signal_6889 ;
    wire signal_6890 ;
    wire signal_6891 ;
    wire signal_6892 ;
    wire signal_6893 ;
    wire signal_6894 ;
    wire signal_6895 ;
    wire signal_6896 ;
    wire signal_6897 ;
    wire signal_6898 ;
    wire signal_6899 ;
    wire signal_6900 ;
    wire signal_6901 ;
    wire signal_6902 ;
    wire signal_6903 ;
    wire signal_6904 ;
    wire signal_6905 ;
    wire signal_6906 ;
    wire signal_6907 ;
    wire signal_6908 ;
    wire signal_6909 ;
    wire signal_6910 ;
    wire signal_6911 ;
    wire signal_6912 ;
    wire signal_6913 ;
    wire signal_6914 ;
    wire signal_6915 ;
    wire signal_6916 ;
    wire signal_6917 ;
    wire signal_6918 ;
    wire signal_6919 ;
    wire signal_6920 ;
    wire signal_6921 ;
    wire signal_6922 ;
    wire signal_6923 ;
    wire signal_6924 ;
    wire signal_6925 ;
    wire signal_6926 ;
    wire signal_6927 ;
    wire signal_6928 ;
    wire signal_6929 ;
    wire signal_6930 ;
    wire signal_6931 ;
    wire signal_6932 ;
    wire signal_6933 ;
    wire signal_6934 ;
    wire signal_6935 ;
    wire signal_6936 ;
    wire signal_6937 ;
    wire signal_6938 ;
    wire signal_6939 ;
    wire signal_6940 ;
    wire signal_6941 ;
    wire signal_6942 ;
    wire signal_6943 ;
    wire signal_6944 ;
    wire signal_6945 ;
    wire signal_6946 ;
    wire signal_6947 ;
    wire signal_6948 ;
    wire signal_6949 ;
    wire signal_6950 ;
    wire signal_6951 ;
    wire signal_6952 ;
    wire signal_6953 ;
    wire signal_6954 ;
    wire signal_6955 ;
    wire signal_6956 ;
    wire signal_6957 ;
    wire signal_6958 ;
    wire signal_6959 ;
    wire signal_6960 ;
    wire signal_6961 ;
    wire signal_6962 ;
    wire signal_6963 ;
    wire signal_6964 ;
    wire signal_6965 ;
    wire signal_6966 ;
    wire signal_6967 ;
    wire signal_6968 ;
    wire signal_6969 ;
    wire signal_6970 ;
    wire signal_6971 ;
    wire signal_6972 ;
    wire signal_6973 ;
    wire signal_6974 ;
    wire signal_6975 ;
    wire signal_6976 ;
    wire signal_6977 ;
    wire signal_6978 ;
    wire signal_6979 ;
    wire signal_6980 ;
    wire signal_6981 ;
    wire signal_6982 ;
    wire signal_6983 ;
    wire signal_6984 ;
    wire signal_6985 ;
    wire signal_6986 ;
    wire signal_6987 ;
    wire signal_6988 ;
    wire signal_6989 ;
    wire signal_6990 ;
    wire signal_6991 ;
    wire signal_6992 ;
    wire signal_6993 ;
    wire signal_6994 ;
    wire signal_6995 ;
    wire signal_6996 ;
    wire signal_6997 ;
    wire signal_6998 ;
    wire signal_6999 ;
    wire signal_7000 ;
    wire signal_7001 ;
    wire signal_7002 ;
    wire signal_7003 ;
    wire signal_7004 ;
    wire signal_7005 ;
    wire signal_7006 ;
    wire signal_7007 ;
    wire signal_7008 ;
    wire signal_7009 ;
    wire signal_7010 ;
    wire signal_7011 ;
    wire signal_7012 ;
    wire signal_7013 ;
    wire signal_7014 ;
    wire signal_7015 ;
    wire signal_7016 ;
    wire signal_7017 ;
    wire signal_7018 ;
    wire signal_7019 ;
    wire signal_7020 ;
    wire signal_7021 ;
    wire signal_7022 ;
    wire signal_7023 ;
    wire signal_7024 ;
    wire signal_7025 ;
    wire signal_7026 ;
    wire signal_7027 ;
    wire signal_7028 ;
    wire signal_7029 ;
    wire signal_7030 ;
    wire signal_7031 ;
    wire signal_7032 ;
    wire signal_7033 ;
    wire signal_7034 ;
    wire signal_7035 ;
    wire signal_7036 ;
    wire signal_7037 ;
    wire signal_7038 ;
    wire signal_7039 ;
    wire signal_7040 ;
    wire signal_7041 ;
    wire signal_7042 ;
    wire signal_7043 ;
    wire signal_7044 ;
    wire signal_7045 ;
    wire signal_7046 ;
    wire signal_7047 ;
    wire signal_7048 ;
    wire signal_7049 ;
    wire signal_7050 ;
    wire signal_7051 ;
    wire signal_7052 ;
    wire signal_7053 ;
    wire signal_7054 ;
    wire signal_7055 ;
    wire signal_7056 ;
    wire signal_7057 ;
    wire signal_7058 ;
    wire signal_7059 ;
    wire signal_7060 ;
    wire signal_7061 ;
    wire signal_7062 ;
    wire signal_7063 ;
    wire signal_7064 ;
    wire signal_7065 ;
    wire signal_7066 ;
    wire signal_7067 ;
    wire signal_7068 ;
    wire signal_7069 ;
    wire signal_7070 ;
    wire signal_7071 ;
    wire signal_7072 ;
    wire signal_7073 ;
    wire signal_7074 ;
    wire signal_7075 ;
    wire signal_7076 ;
    wire signal_7077 ;
    wire signal_7078 ;
    wire signal_7079 ;
    wire signal_7080 ;
    wire signal_7081 ;
    wire signal_7082 ;
    wire signal_7083 ;
    wire signal_7084 ;
    wire signal_7085 ;
    wire signal_7086 ;
    wire signal_7087 ;
    wire signal_7088 ;
    wire signal_7089 ;
    wire signal_7090 ;
    wire signal_7091 ;
    wire signal_7092 ;
    wire signal_7093 ;
    wire signal_7094 ;
    wire signal_7095 ;
    wire signal_7096 ;
    wire signal_7097 ;
    wire signal_7098 ;
    wire signal_7099 ;
    wire signal_7100 ;
    wire signal_7101 ;
    wire signal_7102 ;
    wire signal_7103 ;
    wire signal_7104 ;
    wire signal_7105 ;
    wire signal_7106 ;
    wire signal_7107 ;
    wire signal_7108 ;
    wire signal_7109 ;
    wire signal_7110 ;
    wire signal_7111 ;
    wire signal_7112 ;
    wire signal_7113 ;
    wire signal_7114 ;
    wire signal_7115 ;
    wire signal_7116 ;
    wire signal_7117 ;
    wire signal_7118 ;
    wire signal_7119 ;
    wire signal_7120 ;
    wire signal_7121 ;
    wire signal_7122 ;
    wire signal_7123 ;
    wire signal_7124 ;
    wire signal_7125 ;
    wire signal_7126 ;
    wire signal_7127 ;
    wire signal_7128 ;
    wire signal_7129 ;
    wire signal_7130 ;
    wire signal_7131 ;
    wire signal_7132 ;
    wire signal_7133 ;
    wire signal_7134 ;
    wire signal_7135 ;
    wire signal_7136 ;
    wire signal_7137 ;
    wire signal_7138 ;
    wire signal_7139 ;
    wire signal_7140 ;
    wire signal_7141 ;
    wire signal_7142 ;
    wire signal_7143 ;
    wire signal_7144 ;
    wire signal_7145 ;
    wire signal_7146 ;
    wire signal_7147 ;
    wire signal_7148 ;
    wire signal_7149 ;
    wire signal_7150 ;
    wire signal_7151 ;
    wire signal_7152 ;
    wire signal_7153 ;
    wire signal_7154 ;
    wire signal_7155 ;
    wire signal_7156 ;
    wire signal_7157 ;
    wire signal_7158 ;
    wire signal_7159 ;
    wire signal_7160 ;
    wire signal_7161 ;
    wire signal_7162 ;
    wire signal_7163 ;
    wire signal_7164 ;
    wire signal_7165 ;
    wire signal_7166 ;
    wire signal_7167 ;
    wire signal_7168 ;
    wire signal_7169 ;
    wire signal_7170 ;
    wire signal_7171 ;
    wire signal_7172 ;
    wire signal_7173 ;
    wire signal_7174 ;
    wire signal_7175 ;
    wire signal_7176 ;
    wire signal_7177 ;
    wire signal_7178 ;
    wire signal_7179 ;
    wire signal_7180 ;
    wire signal_7181 ;
    wire signal_7182 ;
    wire signal_7183 ;
    wire signal_7184 ;
    wire signal_7185 ;
    wire signal_7186 ;
    wire signal_7187 ;
    wire signal_7188 ;
    wire signal_7189 ;
    wire signal_7190 ;
    wire signal_7191 ;
    wire signal_7192 ;
    wire signal_7193 ;
    wire signal_7194 ;
    wire signal_7195 ;
    wire signal_7196 ;
    wire signal_7197 ;
    wire signal_7198 ;
    wire signal_7199 ;
    wire signal_7200 ;
    wire signal_7201 ;
    wire signal_7202 ;
    wire signal_7203 ;
    wire signal_7204 ;
    wire signal_7205 ;
    wire signal_7206 ;
    wire signal_7207 ;
    wire signal_7208 ;
    wire signal_7209 ;
    wire signal_7210 ;
    wire signal_7211 ;
    wire signal_7212 ;
    wire signal_7213 ;
    wire signal_7214 ;
    wire signal_7215 ;
    wire signal_7216 ;
    wire signal_7217 ;
    wire signal_7218 ;
    wire signal_7219 ;
    wire signal_7220 ;
    wire signal_7221 ;
    wire signal_7222 ;
    wire signal_7223 ;
    wire signal_7224 ;
    wire signal_7225 ;
    wire signal_7226 ;
    wire signal_7227 ;
    wire signal_7228 ;
    wire signal_7229 ;
    wire signal_7230 ;
    wire signal_7231 ;
    wire signal_7232 ;
    wire signal_7233 ;
    wire signal_7234 ;
    wire signal_7235 ;
    wire signal_7236 ;
    wire signal_7237 ;
    wire signal_7238 ;
    wire signal_7239 ;
    wire signal_7240 ;
    wire signal_7241 ;
    wire signal_7242 ;
    wire signal_7243 ;
    wire signal_7244 ;
    wire signal_7245 ;
    wire signal_7246 ;
    wire signal_7247 ;
    wire signal_7248 ;
    wire signal_7249 ;
    wire signal_7250 ;
    wire signal_7251 ;
    wire signal_7252 ;
    wire signal_7253 ;
    wire signal_7254 ;
    wire signal_7255 ;
    wire signal_7256 ;
    wire signal_7257 ;
    wire signal_7258 ;
    wire signal_7259 ;
    wire signal_7260 ;
    wire signal_7261 ;
    wire signal_7262 ;
    wire signal_7263 ;
    wire signal_7264 ;
    wire signal_7265 ;
    wire signal_7266 ;
    wire signal_7267 ;
    wire signal_7268 ;
    wire signal_7269 ;
    wire signal_7270 ;
    wire signal_7271 ;
    wire signal_7272 ;
    wire signal_7273 ;
    wire signal_7274 ;
    wire signal_7275 ;
    wire signal_7276 ;
    wire signal_7277 ;
    wire signal_7278 ;
    wire signal_7279 ;
    wire signal_7280 ;
    wire signal_7281 ;
    wire signal_7282 ;
    wire signal_7283 ;
    wire signal_7284 ;
    wire signal_7285 ;
    wire signal_7286 ;
    wire signal_7287 ;
    wire signal_7288 ;
    wire signal_7289 ;
    wire signal_7290 ;
    wire signal_7291 ;
    wire signal_7292 ;
    wire signal_7293 ;
    wire signal_7294 ;
    wire signal_7295 ;
    wire signal_7296 ;
    wire signal_7297 ;
    wire signal_7298 ;
    wire signal_7299 ;
    wire signal_7300 ;
    wire signal_7301 ;
    wire signal_7302 ;
    wire signal_7303 ;
    wire signal_7304 ;
    wire signal_7305 ;
    wire signal_7306 ;
    wire signal_7307 ;
    wire signal_7308 ;
    wire signal_7309 ;
    wire signal_7310 ;
    wire signal_7311 ;
    wire signal_7312 ;
    wire signal_7313 ;
    wire signal_7314 ;
    wire signal_7315 ;
    wire signal_7316 ;
    wire signal_7317 ;
    wire signal_7318 ;
    wire signal_7319 ;
    wire signal_7320 ;
    wire signal_7321 ;
    wire signal_7322 ;
    wire signal_7323 ;
    wire signal_7324 ;
    wire signal_7325 ;
    wire signal_7326 ;
    wire signal_7327 ;
    wire signal_7328 ;
    wire signal_7329 ;
    wire signal_7330 ;
    wire signal_7331 ;
    wire signal_7332 ;
    wire signal_7333 ;
    wire signal_7334 ;
    wire signal_7335 ;
    wire signal_7336 ;
    wire signal_7337 ;
    wire signal_7338 ;
    wire signal_7339 ;
    wire signal_7340 ;
    wire signal_7341 ;
    wire signal_7342 ;
    wire signal_7343 ;
    wire signal_7344 ;
    wire signal_7345 ;
    wire signal_7346 ;
    wire signal_7347 ;
    wire signal_7348 ;
    wire signal_7349 ;
    wire signal_7350 ;
    wire signal_7351 ;
    wire signal_7352 ;
    wire signal_7353 ;
    wire signal_7354 ;
    wire signal_7355 ;
    wire signal_7356 ;
    wire signal_7357 ;
    wire signal_7358 ;
    wire signal_7359 ;
    wire signal_7360 ;
    wire signal_7361 ;
    wire signal_7362 ;
    wire signal_7363 ;
    wire signal_7364 ;
    wire signal_7365 ;
    wire signal_7366 ;
    wire signal_7367 ;
    wire signal_7368 ;
    wire signal_7369 ;
    wire signal_7370 ;
    wire signal_7371 ;
    wire signal_7372 ;
    wire signal_7373 ;
    wire signal_7374 ;
    wire signal_7375 ;
    wire signal_7376 ;
    wire signal_7377 ;
    wire signal_7378 ;
    wire signal_7379 ;
    wire signal_7380 ;
    wire signal_7381 ;
    wire signal_7382 ;
    wire signal_7383 ;
    wire signal_7384 ;
    wire signal_7385 ;
    wire signal_7386 ;
    wire signal_7387 ;
    wire signal_7388 ;
    wire signal_7389 ;
    wire signal_7390 ;
    wire signal_7391 ;
    wire signal_7392 ;
    wire signal_7393 ;
    wire signal_7394 ;
    wire signal_7395 ;
    wire signal_7396 ;
    wire signal_7397 ;
    wire signal_7398 ;
    wire signal_7399 ;
    wire signal_7400 ;
    wire signal_7401 ;
    wire signal_7402 ;
    wire signal_7403 ;
    wire signal_7404 ;
    wire signal_7405 ;
    wire signal_7406 ;
    wire signal_7407 ;
    wire signal_7408 ;
    wire signal_7409 ;
    wire signal_7410 ;
    wire signal_7411 ;
    wire signal_7412 ;
    wire signal_7413 ;
    wire signal_7414 ;
    wire signal_7415 ;
    wire signal_7416 ;
    wire signal_7417 ;
    wire signal_7418 ;
    wire signal_7419 ;
    wire signal_7420 ;
    wire signal_7421 ;
    wire signal_7422 ;
    wire signal_7423 ;
    wire signal_7424 ;
    wire signal_7425 ;
    wire signal_7426 ;
    wire signal_7427 ;
    wire signal_7428 ;
    wire signal_7429 ;
    wire signal_7430 ;
    wire signal_7431 ;
    wire signal_7432 ;
    wire signal_7433 ;
    wire signal_7434 ;
    wire signal_7435 ;
    wire signal_7436 ;
    wire signal_7437 ;
    wire signal_7438 ;
    wire signal_7439 ;
    wire signal_7440 ;
    wire signal_7441 ;
    wire signal_7442 ;
    wire signal_7443 ;
    wire signal_7444 ;
    wire signal_7445 ;
    wire signal_7446 ;
    wire signal_7447 ;
    wire signal_7448 ;
    wire signal_7449 ;
    wire signal_7450 ;
    wire signal_7451 ;
    wire signal_7452 ;
    wire signal_7453 ;
    wire signal_7454 ;
    wire signal_7455 ;
    wire signal_7456 ;
    wire signal_7457 ;
    wire signal_7458 ;
    wire signal_7459 ;
    wire signal_7460 ;
    wire signal_7461 ;
    wire signal_7462 ;
    wire signal_7463 ;
    wire signal_7464 ;
    wire signal_7465 ;
    wire signal_7466 ;
    wire signal_7467 ;
    wire signal_7468 ;
    wire signal_7469 ;
    wire signal_7470 ;
    wire signal_7471 ;
    wire signal_7472 ;
    wire signal_7473 ;
    wire signal_7474 ;
    wire signal_7475 ;
    wire signal_7476 ;
    wire signal_7477 ;
    wire signal_7478 ;
    wire signal_7479 ;
    wire signal_7480 ;
    wire signal_7481 ;
    wire signal_7482 ;
    wire signal_7483 ;
    wire signal_7484 ;
    wire signal_7485 ;
    wire signal_7486 ;
    wire signal_7487 ;
    wire signal_7488 ;
    wire signal_7489 ;
    wire signal_7490 ;
    wire signal_7491 ;
    wire signal_7492 ;
    wire signal_7493 ;
    wire signal_7494 ;
    wire signal_7495 ;
    wire signal_7496 ;
    wire signal_7497 ;
    wire signal_7498 ;
    wire signal_7499 ;
    wire signal_7500 ;
    wire signal_7501 ;
    wire signal_7502 ;
    wire signal_7503 ;
    wire signal_7504 ;
    wire signal_7505 ;
    wire signal_7506 ;
    wire signal_7507 ;
    wire signal_7508 ;
    wire signal_7509 ;
    wire signal_7510 ;
    wire signal_7511 ;
    wire signal_7512 ;
    wire signal_7513 ;
    wire signal_7514 ;
    wire signal_7515 ;
    wire signal_7516 ;
    wire signal_7517 ;
    wire signal_7518 ;
    wire signal_7519 ;
    wire signal_7520 ;
    wire signal_7521 ;
    wire signal_7522 ;
    wire signal_7523 ;
    wire signal_7524 ;
    wire signal_7525 ;
    wire signal_7526 ;
    wire signal_7527 ;
    wire signal_7528 ;
    wire signal_7529 ;
    wire signal_7530 ;
    wire signal_7531 ;
    wire signal_7532 ;
    wire signal_7533 ;
    wire signal_7534 ;
    wire signal_7535 ;
    wire signal_7536 ;
    wire signal_7537 ;
    wire signal_7538 ;
    wire signal_7539 ;
    wire signal_7540 ;
    wire signal_7541 ;
    wire signal_7542 ;
    wire signal_7543 ;
    wire signal_7544 ;
    wire signal_7545 ;
    wire signal_7546 ;
    wire signal_7547 ;
    wire signal_7548 ;
    wire signal_7549 ;
    wire signal_7550 ;
    wire signal_7551 ;
    wire signal_7552 ;
    wire signal_7553 ;
    wire signal_7554 ;
    wire signal_7555 ;
    wire signal_7556 ;
    wire signal_7557 ;
    wire signal_7558 ;
    wire signal_7559 ;
    wire signal_7560 ;
    wire signal_7561 ;
    wire signal_7562 ;
    wire signal_7563 ;
    wire signal_7564 ;
    wire signal_7565 ;
    wire signal_7566 ;
    wire signal_7567 ;
    wire signal_7568 ;
    wire signal_7569 ;
    wire signal_7570 ;
    wire signal_7571 ;
    wire signal_7572 ;
    wire signal_7573 ;
    wire signal_7574 ;
    wire signal_7575 ;
    wire signal_7576 ;
    wire signal_7577 ;
    wire signal_7578 ;
    wire signal_7579 ;
    wire signal_7580 ;
    wire signal_7581 ;
    wire signal_7582 ;
    wire signal_7583 ;
    wire signal_7584 ;
    wire signal_7585 ;
    wire signal_7586 ;
    wire signal_7587 ;
    wire signal_7588 ;
    wire signal_7589 ;
    wire signal_7590 ;
    wire signal_7591 ;
    wire signal_7592 ;
    wire signal_7593 ;
    wire signal_7594 ;
    wire signal_7595 ;
    wire signal_7596 ;
    wire signal_7597 ;
    wire signal_7598 ;
    wire signal_7599 ;
    wire signal_7600 ;
    wire signal_7601 ;
    wire signal_7602 ;
    wire signal_7603 ;
    wire signal_7604 ;
    wire signal_7605 ;
    wire signal_7606 ;
    wire signal_7607 ;
    wire signal_7608 ;
    wire signal_7609 ;
    wire signal_7610 ;
    wire signal_7611 ;
    wire signal_7612 ;
    wire signal_7613 ;
    wire signal_7614 ;
    wire signal_7615 ;
    wire signal_7616 ;
    wire signal_7617 ;
    wire signal_7618 ;
    wire signal_7619 ;
    wire signal_7620 ;
    wire signal_7621 ;
    wire signal_7622 ;
    wire signal_7623 ;
    wire signal_7624 ;
    wire signal_7625 ;
    wire signal_7626 ;
    wire signal_7627 ;
    wire signal_7628 ;
    wire signal_7629 ;
    wire signal_7630 ;
    wire signal_7631 ;
    wire signal_7632 ;
    wire signal_7633 ;
    wire signal_7634 ;
    wire signal_7635 ;
    wire signal_7636 ;
    wire signal_7637 ;
    wire signal_7638 ;
    wire signal_7639 ;
    wire signal_7640 ;
    wire signal_7641 ;
    wire signal_7642 ;
    wire signal_7643 ;
    wire signal_7644 ;
    wire signal_7645 ;
    wire signal_7646 ;
    wire signal_7647 ;
    wire signal_7648 ;
    wire signal_7649 ;
    wire signal_7650 ;
    wire signal_7651 ;
    wire signal_7652 ;
    wire signal_7653 ;
    wire signal_7654 ;
    wire signal_7655 ;
    wire signal_7656 ;
    wire signal_7657 ;
    wire signal_7658 ;
    wire signal_7659 ;
    wire signal_7660 ;
    wire signal_7661 ;
    wire signal_7662 ;
    wire signal_7663 ;
    wire signal_7664 ;
    wire signal_7665 ;
    wire signal_7666 ;
    wire signal_7667 ;
    wire signal_7668 ;
    wire signal_7669 ;
    wire signal_7670 ;
    wire signal_7671 ;
    wire signal_7672 ;
    wire signal_7673 ;
    wire signal_7674 ;
    wire signal_7675 ;
    wire signal_7676 ;
    wire signal_7677 ;
    wire signal_7678 ;
    wire signal_7679 ;
    wire signal_7680 ;
    wire signal_7681 ;
    wire signal_7682 ;
    wire signal_7683 ;
    wire signal_7684 ;
    wire signal_7685 ;
    wire signal_7686 ;
    wire signal_7687 ;
    wire signal_7688 ;
    wire signal_7689 ;
    wire signal_7690 ;
    wire signal_7691 ;
    wire signal_7692 ;
    wire signal_7693 ;
    wire signal_7694 ;
    wire signal_7695 ;
    wire signal_7696 ;
    wire signal_7697 ;
    wire signal_7698 ;
    wire signal_7699 ;
    wire signal_7700 ;
    wire signal_7701 ;
    wire signal_7702 ;
    wire signal_7703 ;
    wire signal_7704 ;
    wire signal_7705 ;
    wire signal_7706 ;
    wire signal_7707 ;
    wire signal_7708 ;
    wire signal_7709 ;
    wire signal_7710 ;
    wire signal_7711 ;
    wire signal_7712 ;
    wire signal_7713 ;
    wire signal_7714 ;
    wire signal_7715 ;
    wire signal_7716 ;
    wire signal_7717 ;
    wire signal_7718 ;
    wire signal_7719 ;
    wire signal_7720 ;
    wire signal_7721 ;
    wire signal_7722 ;
    wire signal_7723 ;
    wire signal_7724 ;
    wire signal_7725 ;
    wire signal_7726 ;
    wire signal_7727 ;
    wire signal_7728 ;
    wire signal_7729 ;
    wire signal_7730 ;
    wire signal_7731 ;
    wire signal_7732 ;
    wire signal_7733 ;
    wire signal_7734 ;
    wire signal_7735 ;
    wire signal_7736 ;
    wire signal_7737 ;
    wire signal_7738 ;
    wire signal_7739 ;
    wire signal_7740 ;
    wire signal_7741 ;
    wire signal_7742 ;
    wire signal_7743 ;
    wire signal_7744 ;
    wire signal_7745 ;
    wire signal_7746 ;
    wire signal_7747 ;
    wire signal_7748 ;
    wire signal_7749 ;
    wire signal_7750 ;
    wire signal_7751 ;
    wire signal_7752 ;
    wire signal_7753 ;
    wire signal_7754 ;
    wire signal_7755 ;
    wire signal_7756 ;
    wire signal_7757 ;
    wire signal_7758 ;
    wire signal_7759 ;
    wire signal_7760 ;
    wire signal_7761 ;
    wire signal_7762 ;
    wire signal_7763 ;
    wire signal_7764 ;
    wire signal_7765 ;
    wire signal_7766 ;
    wire signal_7767 ;
    wire signal_7768 ;
    wire signal_7769 ;
    wire signal_7770 ;
    wire signal_7771 ;
    wire signal_7772 ;
    wire signal_7773 ;
    wire signal_7774 ;
    wire signal_7775 ;
    wire signal_7776 ;
    wire signal_7777 ;
    wire signal_7778 ;
    wire signal_7779 ;
    wire signal_7780 ;
    wire signal_7781 ;
    wire signal_7782 ;
    wire signal_7783 ;
    wire signal_7784 ;
    wire signal_7785 ;
    wire signal_7786 ;
    wire signal_7787 ;
    wire signal_7788 ;
    wire signal_7789 ;
    wire signal_7790 ;
    wire signal_7791 ;
    wire signal_7792 ;
    wire signal_7793 ;
    wire signal_7794 ;
    wire signal_7795 ;
    wire signal_7796 ;
    wire signal_7797 ;
    wire signal_7798 ;
    wire signal_7799 ;
    wire signal_7800 ;
    wire signal_7801 ;
    wire signal_7802 ;
    wire signal_7803 ;
    wire signal_7804 ;
    wire signal_7805 ;
    wire signal_7806 ;
    wire signal_7807 ;
    wire signal_7808 ;
    wire signal_7809 ;
    wire signal_7810 ;
    wire signal_7811 ;
    wire signal_7812 ;
    wire signal_7813 ;
    wire signal_7814 ;
    wire signal_7815 ;
    wire signal_7816 ;
    wire signal_7817 ;
    wire signal_7818 ;
    wire signal_7819 ;
    wire signal_7820 ;
    wire signal_7821 ;
    wire signal_7822 ;
    wire signal_7823 ;
    wire signal_7824 ;
    wire signal_7825 ;
    wire signal_7826 ;
    wire signal_7827 ;
    wire signal_7828 ;
    wire signal_7829 ;
    wire signal_7830 ;
    wire signal_7831 ;
    wire signal_7832 ;
    wire signal_7833 ;
    wire signal_7834 ;
    wire signal_7835 ;
    wire signal_7836 ;
    wire signal_7837 ;
    wire signal_7838 ;
    wire signal_7839 ;
    wire signal_7840 ;
    wire signal_7841 ;
    wire signal_7842 ;
    wire signal_7843 ;
    wire signal_7844 ;
    wire signal_7845 ;
    wire signal_7846 ;
    wire signal_7847 ;
    wire signal_7848 ;
    wire signal_7849 ;
    wire signal_7850 ;
    wire signal_7851 ;
    wire signal_7852 ;
    wire signal_7853 ;
    wire signal_7854 ;
    wire signal_7855 ;
    wire signal_7856 ;
    wire signal_7857 ;
    wire signal_7858 ;
    wire signal_7859 ;
    wire signal_7860 ;
    wire signal_7861 ;
    wire signal_7862 ;
    wire signal_7863 ;
    wire signal_7864 ;
    wire signal_7865 ;
    wire signal_7866 ;
    wire signal_7867 ;
    wire signal_7868 ;
    wire signal_7869 ;
    wire signal_7870 ;
    wire signal_7871 ;
    wire signal_7872 ;
    wire signal_7873 ;
    wire signal_7874 ;
    wire signal_7875 ;
    wire signal_7876 ;
    wire signal_7877 ;
    wire signal_7878 ;
    wire signal_7879 ;
    wire signal_7880 ;
    wire signal_7881 ;
    wire signal_7882 ;
    wire signal_7883 ;
    wire signal_7884 ;
    wire signal_7885 ;
    wire signal_7886 ;
    wire signal_7887 ;
    wire signal_7888 ;
    wire signal_7889 ;
    wire signal_7890 ;
    wire signal_7891 ;
    wire signal_7892 ;
    wire signal_7893 ;
    wire signal_7894 ;
    wire signal_7895 ;
    wire signal_7896 ;
    wire signal_7897 ;
    wire signal_7898 ;
    wire signal_7899 ;
    wire signal_7900 ;
    wire signal_7901 ;
    wire signal_7902 ;
    wire signal_7903 ;
    wire signal_7904 ;
    wire signal_7905 ;
    wire signal_7906 ;
    wire signal_7907 ;
    wire signal_7908 ;
    wire signal_7909 ;
    wire signal_7910 ;
    wire signal_7911 ;
    wire signal_7912 ;
    wire signal_7913 ;
    wire signal_7914 ;
    wire signal_7915 ;
    wire signal_7916 ;
    wire signal_7917 ;
    wire signal_7918 ;
    wire signal_7919 ;
    wire signal_7920 ;
    wire signal_7921 ;
    wire signal_7922 ;
    wire signal_7923 ;
    wire signal_7924 ;
    wire signal_7925 ;
    wire signal_7926 ;
    wire signal_7927 ;
    wire signal_7928 ;
    wire signal_7929 ;
    wire signal_7930 ;
    wire signal_7931 ;
    wire signal_7932 ;
    wire signal_7933 ;
    wire signal_7934 ;
    wire signal_7935 ;
    wire signal_7936 ;
    wire signal_7937 ;
    wire signal_7938 ;
    wire signal_7939 ;
    wire signal_7940 ;
    wire signal_7941 ;
    wire signal_7942 ;
    wire signal_7943 ;
    wire signal_7944 ;
    wire signal_7945 ;
    wire signal_7946 ;
    wire signal_7947 ;
    wire signal_7948 ;
    wire signal_7949 ;
    wire signal_7950 ;
    wire signal_7951 ;
    wire signal_7952 ;
    wire signal_7953 ;
    wire signal_7954 ;
    wire signal_7955 ;
    wire signal_7956 ;
    wire signal_7957 ;
    wire signal_7958 ;
    wire signal_7959 ;
    wire signal_7960 ;
    wire signal_7961 ;
    wire signal_7962 ;
    wire signal_7963 ;
    wire signal_7964 ;
    wire signal_7965 ;
    wire signal_7966 ;
    wire signal_7967 ;
    wire signal_7968 ;
    wire signal_7969 ;
    wire signal_7970 ;
    wire signal_7971 ;
    wire signal_7972 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(1)) cell_927 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2393, signal_942}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_928 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2395, signal_943}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_929 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2397, signal_944}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_930 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2399, signal_945}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_931 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2401, signal_946}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_932 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2403, signal_947}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_933 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2405, signal_948}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_934 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2407, signal_949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_949 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .c ({signal_2422, signal_964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_950 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[0], SI_s0[0]}), .c ({signal_2423, signal_965}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_962 ( .a ({signal_2422, signal_964}), .b ({signal_2435, signal_977}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_963 ( .a ({signal_2423, signal_965}), .b ({signal_2436, signal_978}) ) ;

    /* cells in depth 1 */
    buf_clk cell_2385 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( signal_4745 ) ) ;
    buf_clk cell_2387 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( signal_4747 ) ) ;
    buf_clk cell_2389 ( .C ( clk ), .D ( signal_949 ), .Q ( signal_4749 ) ) ;
    buf_clk cell_2391 ( .C ( clk ), .D ( signal_2407 ), .Q ( signal_4751 ) ) ;
    buf_clk cell_2393 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_4753 ) ) ;
    buf_clk cell_2395 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_4755 ) ) ;
    buf_clk cell_2397 ( .C ( clk ), .D ( signal_944 ), .Q ( signal_4757 ) ) ;
    buf_clk cell_2399 ( .C ( clk ), .D ( signal_2397 ), .Q ( signal_4759 ) ) ;
    buf_clk cell_2401 ( .C ( clk ), .D ( signal_942 ), .Q ( signal_4761 ) ) ;
    buf_clk cell_2403 ( .C ( clk ), .D ( signal_2393 ), .Q ( signal_4763 ) ) ;
    buf_clk cell_2405 ( .C ( clk ), .D ( signal_946 ), .Q ( signal_4765 ) ) ;
    buf_clk cell_2407 ( .C ( clk ), .D ( signal_2401 ), .Q ( signal_4767 ) ) ;
    buf_clk cell_2409 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_4769 ) ) ;
    buf_clk cell_2411 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_4771 ) ) ;
    buf_clk cell_2413 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( signal_4773 ) ) ;
    buf_clk cell_2415 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( signal_4775 ) ) ;
    buf_clk cell_2417 ( .C ( clk ), .D ( signal_945 ), .Q ( signal_4777 ) ) ;
    buf_clk cell_2419 ( .C ( clk ), .D ( signal_2399 ), .Q ( signal_4779 ) ) ;
    buf_clk cell_2421 ( .C ( clk ), .D ( signal_948 ), .Q ( signal_4781 ) ) ;
    buf_clk cell_2423 ( .C ( clk ), .D ( signal_2405 ), .Q ( signal_4783 ) ) ;
    buf_clk cell_2425 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( signal_4785 ) ) ;
    buf_clk cell_2427 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( signal_4787 ) ) ;
    buf_clk cell_2429 ( .C ( clk ), .D ( signal_978 ), .Q ( signal_4789 ) ) ;
    buf_clk cell_2431 ( .C ( clk ), .D ( signal_2436 ), .Q ( signal_4791 ) ) ;
    buf_clk cell_2433 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_4793 ) ) ;
    buf_clk cell_2435 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_4795 ) ) ;
    buf_clk cell_2437 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_4797 ) ) ;
    buf_clk cell_2441 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_4801 ) ) ;
    buf_clk cell_2581 ( .C ( clk ), .D ( signal_943 ), .Q ( signal_4941 ) ) ;
    buf_clk cell_2585 ( .C ( clk ), .D ( signal_2395 ), .Q ( signal_4945 ) ) ;
    buf_clk cell_2721 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( signal_5081 ) ) ;
    buf_clk cell_2727 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( signal_5087 ) ) ;
    buf_clk cell_2913 ( .C ( clk ), .D ( signal_947 ), .Q ( signal_5273 ) ) ;
    buf_clk cell_2919 ( .C ( clk ), .D ( signal_2403 ), .Q ( signal_5279 ) ) ;
    buf_clk cell_3061 ( .C ( clk ), .D ( signal_977 ), .Q ( signal_5421 ) ) ;
    buf_clk cell_3069 ( .C ( clk ), .D ( signal_2435 ), .Q ( signal_5429 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_935 ( .a ({SI_s1[3], SI_s0[3]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_2408, signal_950}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_936 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_2409, signal_951}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_937 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_2410, signal_952}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_938 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_2411, signal_953}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_939 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_2412, signal_954}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_940 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_2413, signal_955}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_941 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_2414, signal_956}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_942 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_2415, signal_957}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_943 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_2416, signal_958}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_944 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_2417, signal_959}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_945 ( .a ({SI_s1[3], SI_s0[3]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_2418, signal_960}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_946 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_2419, signal_961}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_947 ( .a ({SI_s1[1], SI_s0[1]}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_2420, signal_962}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_948 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_2421, signal_963}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_951 ( .a ({signal_2408, signal_950}), .b ({signal_2424, signal_966}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_952 ( .a ({signal_2409, signal_951}), .b ({signal_2425, signal_967}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_953 ( .a ({signal_2410, signal_952}), .b ({signal_2426, signal_968}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_954 ( .a ({signal_2411, signal_953}), .b ({signal_2427, signal_969}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_955 ( .a ({signal_2412, signal_954}), .b ({signal_2428, signal_970}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_956 ( .a ({signal_2414, signal_956}), .b ({signal_2429, signal_971}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_957 ( .a ({signal_2415, signal_957}), .b ({signal_2430, signal_972}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_958 ( .a ({signal_2417, signal_959}), .b ({signal_2431, signal_973}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_959 ( .a ({signal_2418, signal_960}), .b ({signal_2432, signal_974}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_960 ( .a ({signal_2419, signal_961}), .b ({signal_2433, signal_975}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_961 ( .a ({signal_2420, signal_962}), .b ({signal_2434, signal_976}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_964 ( .a ({signal_2395, signal_943}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_2437, signal_979}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_965 ( .a ({signal_2405, signal_948}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_2438, signal_980}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_966 ( .a ({signal_2399, signal_945}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_2439, signal_981}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_967 ( .a ({signal_2397, signal_944}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[17] ), .c ({signal_2440, signal_982}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_968 ( .a ({signal_2397, signal_944}), .b ({signal_2399, signal_945}), .clk ( clk ), .r ( Fresh[18] ), .c ({signal_2441, signal_983}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_969 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2395, signal_943}), .clk ( clk ), .r ( Fresh[19] ), .c ({signal_2442, signal_984}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_970 ( .a ({signal_2393, signal_942}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[20] ), .c ({signal_2443, signal_985}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_971 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[21] ), .c ({signal_2444, signal_986}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_972 ( .a ({signal_2403, signal_947}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[22] ), .c ({signal_2445, signal_987}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_973 ( .a ({signal_2403, signal_947}), .b ({signal_2405, signal_948}), .clk ( clk ), .r ( Fresh[23] ), .c ({signal_2446, signal_988}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_974 ( .a ({signal_2403, signal_947}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[24] ), .c ({signal_2447, signal_989}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_975 ( .a ({signal_2395, signal_943}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[25] ), .c ({signal_2448, signal_990}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_976 ( .a ({signal_2399, signal_945}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[26] ), .c ({signal_2449, signal_991}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_977 ( .a ({signal_2405, signal_948}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[27] ), .c ({signal_2450, signal_992}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_978 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[28] ), .c ({signal_2451, signal_993}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_979 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[29] ), .c ({signal_2452, signal_994}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_980 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[30] ), .c ({signal_2453, signal_995}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_981 ( .a ({signal_2397, signal_944}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[31] ), .c ({signal_2454, signal_996}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_982 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[32] ), .c ({signal_2455, signal_997}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_983 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[33] ), .c ({signal_2456, signal_998}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_984 ( .a ({signal_2393, signal_942}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[34] ), .c ({signal_2457, signal_999}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_985 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2405, signal_948}), .clk ( clk ), .r ( Fresh[35] ), .c ({signal_2458, signal_1000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_986 ( .a ({signal_2393, signal_942}), .b ({signal_2395, signal_943}), .clk ( clk ), .r ( Fresh[36] ), .c ({signal_2459, signal_1001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_987 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2399, signal_945}), .clk ( clk ), .r ( Fresh[37] ), .c ({signal_2460, signal_1002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_989 ( .a ({signal_2401, signal_946}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[38] ), .c ({signal_2462, signal_1004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_990 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2399, signal_945}), .clk ( clk ), .r ( Fresh[39] ), .c ({signal_2463, signal_1005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_991 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[40] ), .c ({signal_2464, signal_1006}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_992 ( .a ({signal_2397, signal_944}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[41] ), .c ({signal_2465, signal_1007}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_993 ( .a ({signal_2403, signal_947}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[42] ), .c ({signal_2466, signal_1008}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_994 ( .a ({signal_2401, signal_946}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[43] ), .c ({signal_2467, signal_1009}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_995 ( .a ({signal_2393, signal_942}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[44] ), .c ({signal_2468, signal_1010}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_996 ( .a ({signal_2397, signal_944}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[45] ), .c ({signal_2469, signal_1011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_997 ( .a ({signal_2399, signal_945}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[46] ), .c ({signal_2470, signal_1012}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_998 ( .a ({signal_2399, signal_945}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[47] ), .c ({signal_2471, signal_1013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1000 ( .a ({signal_2399, signal_945}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[48] ), .c ({signal_2473, signal_1015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1001 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2405, signal_948}), .clk ( clk ), .r ( Fresh[49] ), .c ({signal_2474, signal_1016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1002 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[50] ), .c ({signal_2475, signal_1017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1003 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[51] ), .c ({signal_2476, signal_1018}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1016 ( .a ({signal_2437, signal_979}), .b ({signal_2489, signal_1031}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1017 ( .a ({signal_2438, signal_980}), .b ({signal_2490, signal_1032}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1018 ( .a ({signal_2441, signal_983}), .b ({signal_2491, signal_1033}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1019 ( .a ({signal_2442, signal_984}), .b ({signal_2492, signal_1034}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1020 ( .a ({signal_2444, signal_986}), .b ({signal_2493, signal_1035}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1021 ( .a ({signal_2445, signal_987}), .b ({signal_2494, signal_1036}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1022 ( .a ({signal_2446, signal_988}), .b ({signal_2495, signal_1037}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1023 ( .a ({signal_2447, signal_989}), .b ({signal_2496, signal_1038}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1024 ( .a ({signal_2448, signal_990}), .b ({signal_2497, signal_1039}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1025 ( .a ({signal_2449, signal_991}), .b ({signal_2498, signal_1040}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1026 ( .a ({signal_2450, signal_992}), .b ({signal_2499, signal_1041}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1027 ( .a ({signal_2451, signal_993}), .b ({signal_2500, signal_1042}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1028 ( .a ({signal_2453, signal_995}), .b ({signal_2501, signal_1043}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1029 ( .a ({signal_2454, signal_996}), .b ({signal_2502, signal_1044}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1030 ( .a ({signal_2455, signal_997}), .b ({signal_2503, signal_1045}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1031 ( .a ({signal_2456, signal_998}), .b ({signal_2504, signal_1046}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1032 ( .a ({signal_2458, signal_1000}), .b ({signal_2505, signal_1047}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1034 ( .a ({signal_2462, signal_1004}), .b ({signal_2507, signal_1049}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1035 ( .a ({signal_2463, signal_1005}), .b ({signal_2508, signal_1050}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1036 ( .a ({signal_2464, signal_1006}), .b ({signal_2509, signal_1051}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1037 ( .a ({signal_2466, signal_1008}), .b ({signal_2510, signal_1052}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1038 ( .a ({signal_2467, signal_1009}), .b ({signal_2511, signal_1053}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1039 ( .a ({signal_2471, signal_1013}), .b ({signal_2512, signal_1054}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1041 ( .a ({signal_2473, signal_1015}), .b ({signal_2514, signal_1056}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1042 ( .a ({signal_2474, signal_1016}), .b ({signal_2515, signal_1057}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1043 ( .a ({signal_2475, signal_1017}), .b ({signal_2516, signal_1058}) ) ;
    buf_clk cell_2386 ( .C ( clk ), .D ( signal_4745 ), .Q ( signal_4746 ) ) ;
    buf_clk cell_2388 ( .C ( clk ), .D ( signal_4747 ), .Q ( signal_4748 ) ) ;
    buf_clk cell_2390 ( .C ( clk ), .D ( signal_4749 ), .Q ( signal_4750 ) ) ;
    buf_clk cell_2392 ( .C ( clk ), .D ( signal_4751 ), .Q ( signal_4752 ) ) ;
    buf_clk cell_2394 ( .C ( clk ), .D ( signal_4753 ), .Q ( signal_4754 ) ) ;
    buf_clk cell_2396 ( .C ( clk ), .D ( signal_4755 ), .Q ( signal_4756 ) ) ;
    buf_clk cell_2398 ( .C ( clk ), .D ( signal_4757 ), .Q ( signal_4758 ) ) ;
    buf_clk cell_2400 ( .C ( clk ), .D ( signal_4759 ), .Q ( signal_4760 ) ) ;
    buf_clk cell_2402 ( .C ( clk ), .D ( signal_4761 ), .Q ( signal_4762 ) ) ;
    buf_clk cell_2404 ( .C ( clk ), .D ( signal_4763 ), .Q ( signal_4764 ) ) ;
    buf_clk cell_2406 ( .C ( clk ), .D ( signal_4765 ), .Q ( signal_4766 ) ) ;
    buf_clk cell_2408 ( .C ( clk ), .D ( signal_4767 ), .Q ( signal_4768 ) ) ;
    buf_clk cell_2410 ( .C ( clk ), .D ( signal_4769 ), .Q ( signal_4770 ) ) ;
    buf_clk cell_2412 ( .C ( clk ), .D ( signal_4771 ), .Q ( signal_4772 ) ) ;
    buf_clk cell_2414 ( .C ( clk ), .D ( signal_4773 ), .Q ( signal_4774 ) ) ;
    buf_clk cell_2416 ( .C ( clk ), .D ( signal_4775 ), .Q ( signal_4776 ) ) ;
    buf_clk cell_2418 ( .C ( clk ), .D ( signal_4777 ), .Q ( signal_4778 ) ) ;
    buf_clk cell_2420 ( .C ( clk ), .D ( signal_4779 ), .Q ( signal_4780 ) ) ;
    buf_clk cell_2422 ( .C ( clk ), .D ( signal_4781 ), .Q ( signal_4782 ) ) ;
    buf_clk cell_2424 ( .C ( clk ), .D ( signal_4783 ), .Q ( signal_4784 ) ) ;
    buf_clk cell_2426 ( .C ( clk ), .D ( signal_4785 ), .Q ( signal_4786 ) ) ;
    buf_clk cell_2428 ( .C ( clk ), .D ( signal_4787 ), .Q ( signal_4788 ) ) ;
    buf_clk cell_2430 ( .C ( clk ), .D ( signal_4789 ), .Q ( signal_4790 ) ) ;
    buf_clk cell_2432 ( .C ( clk ), .D ( signal_4791 ), .Q ( signal_4792 ) ) ;
    buf_clk cell_2434 ( .C ( clk ), .D ( signal_4793 ), .Q ( signal_4794 ) ) ;
    buf_clk cell_2436 ( .C ( clk ), .D ( signal_4795 ), .Q ( signal_4796 ) ) ;
    buf_clk cell_2438 ( .C ( clk ), .D ( signal_4797 ), .Q ( signal_4798 ) ) ;
    buf_clk cell_2442 ( .C ( clk ), .D ( signal_4801 ), .Q ( signal_4802 ) ) ;
    buf_clk cell_2582 ( .C ( clk ), .D ( signal_4941 ), .Q ( signal_4942 ) ) ;
    buf_clk cell_2586 ( .C ( clk ), .D ( signal_4945 ), .Q ( signal_4946 ) ) ;
    buf_clk cell_2722 ( .C ( clk ), .D ( signal_5081 ), .Q ( signal_5082 ) ) ;
    buf_clk cell_2728 ( .C ( clk ), .D ( signal_5087 ), .Q ( signal_5088 ) ) ;
    buf_clk cell_2914 ( .C ( clk ), .D ( signal_5273 ), .Q ( signal_5274 ) ) ;
    buf_clk cell_2920 ( .C ( clk ), .D ( signal_5279 ), .Q ( signal_5280 ) ) ;
    buf_clk cell_3062 ( .C ( clk ), .D ( signal_5421 ), .Q ( signal_5422 ) ) ;
    buf_clk cell_3070 ( .C ( clk ), .D ( signal_5429 ), .Q ( signal_5430 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_2439 ( .C ( clk ), .D ( signal_4798 ), .Q ( signal_4799 ) ) ;
    buf_clk cell_2443 ( .C ( clk ), .D ( signal_4802 ), .Q ( signal_4803 ) ) ;
    buf_clk cell_2445 ( .C ( clk ), .D ( signal_4778 ), .Q ( signal_4805 ) ) ;
    buf_clk cell_2447 ( .C ( clk ), .D ( signal_4780 ), .Q ( signal_4807 ) ) ;
    buf_clk cell_2449 ( .C ( clk ), .D ( signal_995 ), .Q ( signal_4809 ) ) ;
    buf_clk cell_2451 ( .C ( clk ), .D ( signal_2453 ), .Q ( signal_4811 ) ) ;
    buf_clk cell_2453 ( .C ( clk ), .D ( signal_1010 ), .Q ( signal_4813 ) ) ;
    buf_clk cell_2455 ( .C ( clk ), .D ( signal_2468 ), .Q ( signal_4815 ) ) ;
    buf_clk cell_2457 ( .C ( clk ), .D ( signal_992 ), .Q ( signal_4817 ) ) ;
    buf_clk cell_2459 ( .C ( clk ), .D ( signal_2450 ), .Q ( signal_4819 ) ) ;
    buf_clk cell_2461 ( .C ( clk ), .D ( signal_993 ), .Q ( signal_4821 ) ) ;
    buf_clk cell_2463 ( .C ( clk ), .D ( signal_2451 ), .Q ( signal_4823 ) ) ;
    buf_clk cell_2465 ( .C ( clk ), .D ( signal_1008 ), .Q ( signal_4825 ) ) ;
    buf_clk cell_2467 ( .C ( clk ), .D ( signal_2466 ), .Q ( signal_4827 ) ) ;
    buf_clk cell_2469 ( .C ( clk ), .D ( signal_991 ), .Q ( signal_4829 ) ) ;
    buf_clk cell_2471 ( .C ( clk ), .D ( signal_2449 ), .Q ( signal_4831 ) ) ;
    buf_clk cell_2473 ( .C ( clk ), .D ( signal_959 ), .Q ( signal_4833 ) ) ;
    buf_clk cell_2475 ( .C ( clk ), .D ( signal_2417 ), .Q ( signal_4835 ) ) ;
    buf_clk cell_2477 ( .C ( clk ), .D ( signal_987 ), .Q ( signal_4837 ) ) ;
    buf_clk cell_2479 ( .C ( clk ), .D ( signal_2445 ), .Q ( signal_4839 ) ) ;
    buf_clk cell_2481 ( .C ( clk ), .D ( signal_961 ), .Q ( signal_4841 ) ) ;
    buf_clk cell_2483 ( .C ( clk ), .D ( signal_2419 ), .Q ( signal_4843 ) ) ;
    buf_clk cell_2485 ( .C ( clk ), .D ( signal_979 ), .Q ( signal_4845 ) ) ;
    buf_clk cell_2487 ( .C ( clk ), .D ( signal_2437 ), .Q ( signal_4847 ) ) ;
    buf_clk cell_2489 ( .C ( clk ), .D ( signal_4770 ), .Q ( signal_4849 ) ) ;
    buf_clk cell_2491 ( .C ( clk ), .D ( signal_4772 ), .Q ( signal_4851 ) ) ;
    buf_clk cell_2493 ( .C ( clk ), .D ( signal_960 ), .Q ( signal_4853 ) ) ;
    buf_clk cell_2495 ( .C ( clk ), .D ( signal_2418 ), .Q ( signal_4855 ) ) ;
    buf_clk cell_2497 ( .C ( clk ), .D ( signal_4794 ), .Q ( signal_4857 ) ) ;
    buf_clk cell_2499 ( .C ( clk ), .D ( signal_4796 ), .Q ( signal_4859 ) ) ;
    buf_clk cell_2501 ( .C ( clk ), .D ( signal_950 ), .Q ( signal_4861 ) ) ;
    buf_clk cell_2503 ( .C ( clk ), .D ( signal_2408 ), .Q ( signal_4863 ) ) ;
    buf_clk cell_2505 ( .C ( clk ), .D ( signal_1000 ), .Q ( signal_4865 ) ) ;
    buf_clk cell_2507 ( .C ( clk ), .D ( signal_2458 ), .Q ( signal_4867 ) ) ;
    buf_clk cell_2509 ( .C ( clk ), .D ( signal_4750 ), .Q ( signal_4869 ) ) ;
    buf_clk cell_2511 ( .C ( clk ), .D ( signal_4752 ), .Q ( signal_4871 ) ) ;
    buf_clk cell_2513 ( .C ( clk ), .D ( signal_4766 ), .Q ( signal_4873 ) ) ;
    buf_clk cell_2515 ( .C ( clk ), .D ( signal_4768 ), .Q ( signal_4875 ) ) ;
    buf_clk cell_2517 ( .C ( clk ), .D ( signal_989 ), .Q ( signal_4877 ) ) ;
    buf_clk cell_2519 ( .C ( clk ), .D ( signal_2447 ), .Q ( signal_4879 ) ) ;
    buf_clk cell_2521 ( .C ( clk ), .D ( signal_4782 ), .Q ( signal_4881 ) ) ;
    buf_clk cell_2523 ( .C ( clk ), .D ( signal_4784 ), .Q ( signal_4883 ) ) ;
    buf_clk cell_2525 ( .C ( clk ), .D ( signal_986 ), .Q ( signal_4885 ) ) ;
    buf_clk cell_2527 ( .C ( clk ), .D ( signal_2444 ), .Q ( signal_4887 ) ) ;
    buf_clk cell_2529 ( .C ( clk ), .D ( signal_1032 ), .Q ( signal_4889 ) ) ;
    buf_clk cell_2531 ( .C ( clk ), .D ( signal_2490 ), .Q ( signal_4891 ) ) ;
    buf_clk cell_2533 ( .C ( clk ), .D ( signal_1016 ), .Q ( signal_4893 ) ) ;
    buf_clk cell_2535 ( .C ( clk ), .D ( signal_2474 ), .Q ( signal_4895 ) ) ;
    buf_clk cell_2537 ( .C ( clk ), .D ( signal_4774 ), .Q ( signal_4897 ) ) ;
    buf_clk cell_2539 ( .C ( clk ), .D ( signal_4776 ), .Q ( signal_4899 ) ) ;
    buf_clk cell_2541 ( .C ( clk ), .D ( signal_4786 ), .Q ( signal_4901 ) ) ;
    buf_clk cell_2543 ( .C ( clk ), .D ( signal_4788 ), .Q ( signal_4903 ) ) ;
    buf_clk cell_2545 ( .C ( clk ), .D ( signal_962 ), .Q ( signal_4905 ) ) ;
    buf_clk cell_2547 ( .C ( clk ), .D ( signal_2420 ), .Q ( signal_4907 ) ) ;
    buf_clk cell_2549 ( .C ( clk ), .D ( signal_998 ), .Q ( signal_4909 ) ) ;
    buf_clk cell_2551 ( .C ( clk ), .D ( signal_2456 ), .Q ( signal_4911 ) ) ;
    buf_clk cell_2553 ( .C ( clk ), .D ( signal_1001 ), .Q ( signal_4913 ) ) ;
    buf_clk cell_2555 ( .C ( clk ), .D ( signal_2459 ), .Q ( signal_4915 ) ) ;
    buf_clk cell_2557 ( .C ( clk ), .D ( signal_1009 ), .Q ( signal_4917 ) ) ;
    buf_clk cell_2559 ( .C ( clk ), .D ( signal_2467 ), .Q ( signal_4919 ) ) ;
    buf_clk cell_2561 ( .C ( clk ), .D ( signal_953 ), .Q ( signal_4921 ) ) ;
    buf_clk cell_2563 ( .C ( clk ), .D ( signal_2411 ), .Q ( signal_4923 ) ) ;
    buf_clk cell_2565 ( .C ( clk ), .D ( signal_988 ), .Q ( signal_4925 ) ) ;
    buf_clk cell_2567 ( .C ( clk ), .D ( signal_2446 ), .Q ( signal_4927 ) ) ;
    buf_clk cell_2569 ( .C ( clk ), .D ( signal_4754 ), .Q ( signal_4929 ) ) ;
    buf_clk cell_2571 ( .C ( clk ), .D ( signal_4756 ), .Q ( signal_4931 ) ) ;
    buf_clk cell_2573 ( .C ( clk ), .D ( signal_1004 ), .Q ( signal_4933 ) ) ;
    buf_clk cell_2575 ( .C ( clk ), .D ( signal_2462 ), .Q ( signal_4935 ) ) ;
    buf_clk cell_2577 ( .C ( clk ), .D ( signal_957 ), .Q ( signal_4937 ) ) ;
    buf_clk cell_2579 ( .C ( clk ), .D ( signal_2415 ), .Q ( signal_4939 ) ) ;
    buf_clk cell_2583 ( .C ( clk ), .D ( signal_4942 ), .Q ( signal_4943 ) ) ;
    buf_clk cell_2587 ( .C ( clk ), .D ( signal_4946 ), .Q ( signal_4947 ) ) ;
    buf_clk cell_2589 ( .C ( clk ), .D ( signal_984 ), .Q ( signal_4949 ) ) ;
    buf_clk cell_2591 ( .C ( clk ), .D ( signal_2442 ), .Q ( signal_4951 ) ) ;
    buf_clk cell_2593 ( .C ( clk ), .D ( signal_997 ), .Q ( signal_4953 ) ) ;
    buf_clk cell_2595 ( .C ( clk ), .D ( signal_2455 ), .Q ( signal_4955 ) ) ;
    buf_clk cell_2597 ( .C ( clk ), .D ( signal_1007 ), .Q ( signal_4957 ) ) ;
    buf_clk cell_2599 ( .C ( clk ), .D ( signal_2465 ), .Q ( signal_4959 ) ) ;
    buf_clk cell_2601 ( .C ( clk ), .D ( signal_951 ), .Q ( signal_4961 ) ) ;
    buf_clk cell_2603 ( .C ( clk ), .D ( signal_2409 ), .Q ( signal_4963 ) ) ;
    buf_clk cell_2605 ( .C ( clk ), .D ( signal_981 ), .Q ( signal_4965 ) ) ;
    buf_clk cell_2607 ( .C ( clk ), .D ( signal_2439 ), .Q ( signal_4967 ) ) ;
    buf_clk cell_2609 ( .C ( clk ), .D ( signal_4746 ), .Q ( signal_4969 ) ) ;
    buf_clk cell_2611 ( .C ( clk ), .D ( signal_4748 ), .Q ( signal_4971 ) ) ;
    buf_clk cell_2613 ( .C ( clk ), .D ( signal_990 ), .Q ( signal_4973 ) ) ;
    buf_clk cell_2615 ( .C ( clk ), .D ( signal_2448 ), .Q ( signal_4975 ) ) ;
    buf_clk cell_2617 ( .C ( clk ), .D ( signal_1006 ), .Q ( signal_4977 ) ) ;
    buf_clk cell_2619 ( .C ( clk ), .D ( signal_2464 ), .Q ( signal_4979 ) ) ;
    buf_clk cell_2621 ( .C ( clk ), .D ( signal_983 ), .Q ( signal_4981 ) ) ;
    buf_clk cell_2623 ( .C ( clk ), .D ( signal_2441 ), .Q ( signal_4983 ) ) ;
    buf_clk cell_2625 ( .C ( clk ), .D ( signal_980 ), .Q ( signal_4985 ) ) ;
    buf_clk cell_2627 ( .C ( clk ), .D ( signal_2438 ), .Q ( signal_4987 ) ) ;
    buf_clk cell_2629 ( .C ( clk ), .D ( signal_999 ), .Q ( signal_4989 ) ) ;
    buf_clk cell_2631 ( .C ( clk ), .D ( signal_2457 ), .Q ( signal_4991 ) ) ;
    buf_clk cell_2633 ( .C ( clk ), .D ( signal_972 ), .Q ( signal_4993 ) ) ;
    buf_clk cell_2635 ( .C ( clk ), .D ( signal_2430 ), .Q ( signal_4995 ) ) ;
    buf_clk cell_2637 ( .C ( clk ), .D ( signal_976 ), .Q ( signal_4997 ) ) ;
    buf_clk cell_2639 ( .C ( clk ), .D ( signal_2434 ), .Q ( signal_4999 ) ) ;
    buf_clk cell_2641 ( .C ( clk ), .D ( signal_1057 ), .Q ( signal_5001 ) ) ;
    buf_clk cell_2643 ( .C ( clk ), .D ( signal_2515 ), .Q ( signal_5003 ) ) ;
    buf_clk cell_2645 ( .C ( clk ), .D ( signal_1039 ), .Q ( signal_5005 ) ) ;
    buf_clk cell_2647 ( .C ( clk ), .D ( signal_2497 ), .Q ( signal_5007 ) ) ;
    buf_clk cell_2649 ( .C ( clk ), .D ( signal_1046 ), .Q ( signal_5009 ) ) ;
    buf_clk cell_2651 ( .C ( clk ), .D ( signal_2504 ), .Q ( signal_5011 ) ) ;
    buf_clk cell_2653 ( .C ( clk ), .D ( signal_1005 ), .Q ( signal_5013 ) ) ;
    buf_clk cell_2655 ( .C ( clk ), .D ( signal_2463 ), .Q ( signal_5015 ) ) ;
    buf_clk cell_2657 ( .C ( clk ), .D ( signal_1041 ), .Q ( signal_5017 ) ) ;
    buf_clk cell_2659 ( .C ( clk ), .D ( signal_2499 ), .Q ( signal_5019 ) ) ;
    buf_clk cell_2661 ( .C ( clk ), .D ( signal_1034 ), .Q ( signal_5021 ) ) ;
    buf_clk cell_2663 ( .C ( clk ), .D ( signal_2492 ), .Q ( signal_5023 ) ) ;
    buf_clk cell_2665 ( .C ( clk ), .D ( signal_996 ), .Q ( signal_5025 ) ) ;
    buf_clk cell_2667 ( .C ( clk ), .D ( signal_2454 ), .Q ( signal_5027 ) ) ;
    buf_clk cell_2669 ( .C ( clk ), .D ( signal_994 ), .Q ( signal_5029 ) ) ;
    buf_clk cell_2671 ( .C ( clk ), .D ( signal_2452 ), .Q ( signal_5031 ) ) ;
    buf_clk cell_2673 ( .C ( clk ), .D ( signal_985 ), .Q ( signal_5033 ) ) ;
    buf_clk cell_2675 ( .C ( clk ), .D ( signal_2443 ), .Q ( signal_5035 ) ) ;
    buf_clk cell_2723 ( .C ( clk ), .D ( signal_5082 ), .Q ( signal_5083 ) ) ;
    buf_clk cell_2729 ( .C ( clk ), .D ( signal_5088 ), .Q ( signal_5089 ) ) ;
    buf_clk cell_2813 ( .C ( clk ), .D ( signal_1054 ), .Q ( signal_5173 ) ) ;
    buf_clk cell_2817 ( .C ( clk ), .D ( signal_2512 ), .Q ( signal_5177 ) ) ;
    buf_clk cell_2829 ( .C ( clk ), .D ( signal_952 ), .Q ( signal_5189 ) ) ;
    buf_clk cell_2833 ( .C ( clk ), .D ( signal_2410 ), .Q ( signal_5193 ) ) ;
    buf_clk cell_2881 ( .C ( clk ), .D ( signal_958 ), .Q ( signal_5241 ) ) ;
    buf_clk cell_2885 ( .C ( clk ), .D ( signal_2416 ), .Q ( signal_5245 ) ) ;
    buf_clk cell_2893 ( .C ( clk ), .D ( signal_954 ), .Q ( signal_5253 ) ) ;
    buf_clk cell_2897 ( .C ( clk ), .D ( signal_2412 ), .Q ( signal_5257 ) ) ;
    buf_clk cell_2915 ( .C ( clk ), .D ( signal_5274 ), .Q ( signal_5275 ) ) ;
    buf_clk cell_2921 ( .C ( clk ), .D ( signal_5280 ), .Q ( signal_5281 ) ) ;
    buf_clk cell_2941 ( .C ( clk ), .D ( signal_963 ), .Q ( signal_5301 ) ) ;
    buf_clk cell_2945 ( .C ( clk ), .D ( signal_2421 ), .Q ( signal_5305 ) ) ;
    buf_clk cell_2985 ( .C ( clk ), .D ( signal_4762 ), .Q ( signal_5345 ) ) ;
    buf_clk cell_2989 ( .C ( clk ), .D ( signal_4764 ), .Q ( signal_5349 ) ) ;
    buf_clk cell_3063 ( .C ( clk ), .D ( signal_5422 ), .Q ( signal_5423 ) ) ;
    buf_clk cell_3071 ( .C ( clk ), .D ( signal_5430 ), .Q ( signal_5431 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_988 ( .a ({signal_2409, signal_951}), .b ({signal_2411, signal_953}), .clk ( clk ), .r ( Fresh[52] ), .c ({signal_2461, signal_1003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_999 ( .a ({signal_2410, signal_952}), .b ({signal_2413, signal_955}), .clk ( clk ), .r ( Fresh[53] ), .c ({signal_2472, signal_1014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1004 ( .a ({signal_4748, signal_4746}), .b ({signal_2411, signal_953}), .clk ( clk ), .r ( Fresh[54] ), .c ({signal_2477, signal_1019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1005 ( .a ({signal_2409, signal_951}), .b ({signal_2416, signal_958}), .clk ( clk ), .r ( Fresh[55] ), .c ({signal_2478, signal_1020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1006 ( .a ({signal_4752, signal_4750}), .b ({signal_2411, signal_953}), .clk ( clk ), .r ( Fresh[56] ), .c ({signal_2479, signal_1021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1007 ( .a ({signal_4756, signal_4754}), .b ({signal_2418, signal_960}), .clk ( clk ), .r ( Fresh[57] ), .c ({signal_2480, signal_1022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1008 ( .a ({signal_2415, signal_957}), .b ({signal_2417, signal_959}), .clk ( clk ), .r ( Fresh[58] ), .c ({signal_2481, signal_1023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1009 ( .a ({signal_2409, signal_951}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[59] ), .c ({signal_2482, signal_1024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1010 ( .a ({signal_2409, signal_951}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[60] ), .c ({signal_2483, signal_1025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1011 ( .a ({signal_2413, signal_955}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[61] ), .c ({signal_2484, signal_1026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1012 ( .a ({signal_2411, signal_953}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[62] ), .c ({signal_2485, signal_1027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1013 ( .a ({signal_2408, signal_950}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[63] ), .c ({signal_2486, signal_1028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1014 ( .a ({signal_4760, signal_4758}), .b ({signal_2418, signal_960}), .clk ( clk ), .r ( Fresh[64] ), .c ({signal_2487, signal_1029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1015 ( .a ({signal_2414, signal_956}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[65] ), .c ({signal_2488, signal_1030}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1033 ( .a ({signal_2461, signal_1003}), .b ({signal_2506, signal_1048}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1040 ( .a ({signal_2472, signal_1014}), .b ({signal_2513, signal_1055}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1044 ( .a ({signal_2478, signal_1020}), .b ({signal_2517, signal_1059}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1045 ( .a ({signal_2481, signal_1023}), .b ({signal_2518, signal_1060}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1046 ( .a ({signal_2483, signal_1025}), .b ({signal_2519, signal_1061}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1047 ( .a ({signal_2484, signal_1026}), .b ({signal_2520, signal_1062}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1048 ( .a ({signal_2485, signal_1027}), .b ({signal_2521, signal_1063}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1049 ( .a ({signal_2486, signal_1028}), .b ({signal_2522, signal_1064}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1050 ( .a ({signal_2487, signal_1029}), .b ({signal_2523, signal_1065}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1051 ( .a ({signal_2488, signal_1030}), .b ({signal_2524, signal_1066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1052 ( .a ({signal_4752, signal_4750}), .b ({signal_2437, signal_979}), .clk ( clk ), .r ( Fresh[66] ), .c ({signal_2525, signal_1067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1053 ( .a ({signal_4764, signal_4762}), .b ({signal_2441, signal_983}), .clk ( clk ), .r ( Fresh[67] ), .c ({signal_2526, signal_1068}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1054 ( .a ({signal_2425, signal_967}), .b ({signal_2426, signal_968}), .clk ( clk ), .r ( Fresh[68] ), .c ({signal_2527, signal_1069}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1055 ( .a ({signal_4756, signal_4754}), .b ({signal_2424, signal_966}), .clk ( clk ), .r ( Fresh[69] ), .c ({signal_2528, signal_1070}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1056 ( .a ({signal_4768, signal_4766}), .b ({signal_2438, signal_980}), .clk ( clk ), .r ( Fresh[70] ), .c ({signal_2529, signal_1071}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1057 ( .a ({signal_2410, signal_952}), .b ({signal_2438, signal_980}), .clk ( clk ), .r ( Fresh[71] ), .c ({signal_2530, signal_1072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1058 ( .a ({signal_2443, signal_985}), .b ({signal_2416, signal_958}), .clk ( clk ), .r ( Fresh[72] ), .c ({signal_2531, signal_1073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1059 ( .a ({signal_2409, signal_951}), .b ({signal_2439, signal_981}), .clk ( clk ), .r ( Fresh[73] ), .c ({signal_2532, signal_1074}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1060 ( .a ({signal_2409, signal_951}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[74] ), .c ({signal_2533, signal_1075}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1061 ( .a ({signal_2452, signal_994}), .b ({signal_2457, signal_999}), .clk ( clk ), .r ( Fresh[75] ), .c ({signal_2534, signal_1076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1062 ( .a ({signal_4764, signal_4762}), .b ({signal_2437, signal_979}), .clk ( clk ), .r ( Fresh[76] ), .c ({signal_2535, signal_1077}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1063 ( .a ({signal_2441, signal_983}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[77] ), .c ({signal_2536, signal_1078}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1064 ( .a ({signal_2446, signal_988}), .b ({signal_2460, signal_1002}), .clk ( clk ), .r ( Fresh[78] ), .c ({signal_2537, signal_1079}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1065 ( .a ({signal_4756, signal_4754}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[79] ), .c ({signal_2538, signal_1080}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1066 ( .a ({signal_4772, signal_4770}), .b ({signal_2462, signal_1004}), .clk ( clk ), .r ( Fresh[80] ), .c ({signal_2539, signal_1081}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1067 ( .a ({signal_2441, signal_983}), .b ({signal_2443, signal_985}), .clk ( clk ), .r ( Fresh[81] ), .c ({signal_2540, signal_1082}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1068 ( .a ({signal_2409, signal_951}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[82] ), .c ({signal_2541, signal_1083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1069 ( .a ({signal_2409, signal_951}), .b ({signal_2441, signal_983}), .clk ( clk ), .r ( Fresh[83] ), .c ({signal_2542, signal_1084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1070 ( .a ({signal_2442, signal_984}), .b ({signal_2456, signal_998}), .clk ( clk ), .r ( Fresh[84] ), .c ({signal_2543, signal_1085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1071 ( .a ({signal_2410, signal_952}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[85] ), .c ({signal_2544, signal_1086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1072 ( .a ({signal_2458, signal_1000}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[86] ), .c ({signal_2545, signal_1087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1073 ( .a ({signal_2438, signal_980}), .b ({signal_2442, signal_984}), .clk ( clk ), .r ( Fresh[87] ), .c ({signal_2546, signal_1088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1074 ( .a ({signal_4748, signal_4746}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[88] ), .c ({signal_2547, signal_1089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1075 ( .a ({signal_2411, signal_953}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[89] ), .c ({signal_2548, signal_1090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1076 ( .a ({signal_2442, signal_984}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[90] ), .c ({signal_2549, signal_1091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1077 ( .a ({signal_2409, signal_951}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[91] ), .c ({signal_2550, signal_1092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1078 ( .a ({signal_2437, signal_979}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[92] ), .c ({signal_2551, signal_1093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1079 ( .a ({signal_2408, signal_950}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[93] ), .c ({signal_2552, signal_1094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1080 ( .a ({signal_2442, signal_984}), .b ({signal_2416, signal_958}), .clk ( clk ), .r ( Fresh[94] ), .c ({signal_2553, signal_1095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1081 ( .a ({signal_2437, signal_979}), .b ({signal_2470, signal_1012}), .clk ( clk ), .r ( Fresh[95] ), .c ({signal_2554, signal_1096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1082 ( .a ({signal_2439, signal_981}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[96] ), .c ({signal_2555, signal_1097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1083 ( .a ({signal_2410, signal_952}), .b ({signal_2439, signal_981}), .clk ( clk ), .r ( Fresh[97] ), .c ({signal_2556, signal_1098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1084 ( .a ({signal_4756, signal_4754}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[98] ), .c ({signal_2557, signal_1099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1086 ( .a ({signal_2440, signal_982}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[99] ), .c ({signal_2559, signal_1101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1087 ( .a ({signal_2409, signal_951}), .b ({signal_2440, signal_982}), .clk ( clk ), .r ( Fresh[100] ), .c ({signal_2560, signal_1102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1088 ( .a ({signal_2411, signal_953}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[101] ), .c ({signal_2561, signal_1103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1089 ( .a ({signal_4752, signal_4750}), .b ({signal_2446, signal_988}), .clk ( clk ), .r ( Fresh[102] ), .c ({signal_2562, signal_1104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1090 ( .a ({signal_2441, signal_983}), .b ({signal_2418, signal_960}), .clk ( clk ), .r ( Fresh[103] ), .c ({signal_2563, signal_1105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1091 ( .a ({signal_2410, signal_952}), .b ({signal_2474, signal_1016}), .clk ( clk ), .r ( Fresh[104] ), .c ({signal_2564, signal_1106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1092 ( .a ({signal_4764, signal_4762}), .b ({signal_2462, signal_1004}), .clk ( clk ), .r ( Fresh[105] ), .c ({signal_2565, signal_1107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1093 ( .a ({signal_4776, signal_4774}), .b ({signal_2438, signal_980}), .clk ( clk ), .r ( Fresh[106] ), .c ({signal_2566, signal_1108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1094 ( .a ({signal_2410, signal_952}), .b ({signal_2470, signal_1012}), .clk ( clk ), .r ( Fresh[107] ), .c ({signal_2567, signal_1109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1095 ( .a ({signal_2448, signal_990}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[108] ), .c ({signal_2568, signal_1110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1096 ( .a ({signal_2439, signal_981}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[109] ), .c ({signal_2569, signal_1111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1097 ( .a ({signal_2419, signal_961}), .b ({signal_2471, signal_1013}), .clk ( clk ), .r ( Fresh[110] ), .c ({signal_2570, signal_1112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1098 ( .a ({signal_2439, signal_981}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[111] ), .c ({signal_2571, signal_1113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1099 ( .a ({signal_4780, signal_4778}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[112] ), .c ({signal_2572, signal_1114}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1100 ( .a ({signal_4768, signal_4766}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[113] ), .c ({signal_2573, signal_1115}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1101 ( .a ({signal_4756, signal_4754}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[114] ), .c ({signal_2574, signal_1116}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1102 ( .a ({signal_2444, signal_986}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[115] ), .c ({signal_2575, signal_1117}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1103 ( .a ({signal_4772, signal_4770}), .b ({signal_2460, signal_1002}), .clk ( clk ), .r ( Fresh[116] ), .c ({signal_2576, signal_1118}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1104 ( .a ({signal_2439, signal_981}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[117] ), .c ({signal_2577, signal_1119}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1105 ( .a ({signal_4784, signal_4782}), .b ({signal_2441, signal_983}), .clk ( clk ), .r ( Fresh[118] ), .c ({signal_2578, signal_1120}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1106 ( .a ({signal_2447, signal_989}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[119] ), .c ({signal_2579, signal_1121}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1107 ( .a ({signal_2418, signal_960}), .b ({signal_2476, signal_1018}), .clk ( clk ), .r ( Fresh[120] ), .c ({signal_2580, signal_1122}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1108 ( .a ({signal_2463, signal_1005}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[121] ), .c ({signal_2581, signal_1123}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1109 ( .a ({signal_2438, signal_980}), .b ({signal_2457, signal_999}), .clk ( clk ), .r ( Fresh[122] ), .c ({signal_2582, signal_1124}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1110 ( .a ({signal_2439, signal_981}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[123] ), .c ({signal_2583, signal_1125}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1111 ( .a ({signal_2444, signal_986}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[124] ), .c ({signal_2584, signal_1126}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1112 ( .a ({signal_2438, signal_980}), .b ({signal_2414, signal_956}), .clk ( clk ), .r ( Fresh[125] ), .c ({signal_2585, signal_1127}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1113 ( .a ({signal_2437, signal_979}), .b ({signal_2421, signal_963}), .clk ( clk ), .r ( Fresh[126] ), .c ({signal_2586, signal_1128}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1114 ( .a ({signal_2441, signal_983}), .b ({signal_2474, signal_1016}), .clk ( clk ), .r ( Fresh[127] ), .c ({signal_2587, signal_1129}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1115 ( .a ({signal_2412, signal_954}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[128] ), .c ({signal_2588, signal_1130}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1116 ( .a ({signal_2446, signal_988}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[129] ), .c ({signal_2589, signal_1131}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1117 ( .a ({signal_2409, signal_951}), .b ({signal_2444, signal_986}), .clk ( clk ), .r ( Fresh[130] ), .c ({signal_2590, signal_1132}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1118 ( .a ({signal_2447, signal_989}), .b ({signal_2448, signal_990}), .clk ( clk ), .r ( Fresh[131] ), .c ({signal_2591, signal_1133}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1119 ( .a ({signal_2448, signal_990}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[132] ), .c ({signal_2592, signal_1134}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1120 ( .a ({signal_2446, signal_988}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[133] ), .c ({signal_2593, signal_1135}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1121 ( .a ({signal_2448, signal_990}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[134] ), .c ({signal_2594, signal_1136}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1122 ( .a ({signal_2449, signal_991}), .b ({signal_2453, signal_995}), .clk ( clk ), .r ( Fresh[135] ), .c ({signal_2595, signal_1137}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1123 ( .a ({signal_4776, signal_4774}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[136] ), .c ({signal_2596, signal_1138}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1125 ( .a ({signal_2440, signal_982}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[137] ), .c ({signal_2598, signal_1140}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1126 ( .a ({signal_2415, signal_957}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[138] ), .c ({signal_2599, signal_1141}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1127 ( .a ({signal_2416, signal_958}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[139] ), .c ({signal_2600, signal_1142}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1128 ( .a ({signal_2459, signal_1001}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[140] ), .c ({signal_2601, signal_1143}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1129 ( .a ({signal_2442, signal_984}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[141] ), .c ({signal_2602, signal_1144}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1130 ( .a ({signal_4772, signal_4770}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[142] ), .c ({signal_2603, signal_1145}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1131 ( .a ({signal_2450, signal_992}), .b ({signal_2464, signal_1006}), .clk ( clk ), .r ( Fresh[143] ), .c ({signal_2604, signal_1146}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1133 ( .a ({signal_2412, signal_954}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[144] ), .c ({signal_2606, signal_1148}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1134 ( .a ({signal_2447, signal_989}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[145] ), .c ({signal_2607, signal_1149}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1135 ( .a ({signal_2462, signal_1004}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[146] ), .c ({signal_2608, signal_1150}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1136 ( .a ({signal_4788, signal_4786}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[147] ), .c ({signal_2609, signal_1151}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1137 ( .a ({signal_2463, signal_1005}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[148] ), .c ({signal_2610, signal_1152}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1138 ( .a ({signal_4752, signal_4750}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[149] ), .c ({signal_2611, signal_1153}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1139 ( .a ({signal_2411, signal_953}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[150] ), .c ({signal_2612, signal_1154}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1141 ( .a ({signal_2458, signal_1000}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[151] ), .c ({signal_2614, signal_1156}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1142 ( .a ({signal_2449, signal_991}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[152] ), .c ({signal_2615, signal_1157}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1143 ( .a ({signal_4756, signal_4754}), .b ({signal_2446, signal_988}), .clk ( clk ), .r ( Fresh[153] ), .c ({signal_2616, signal_1158}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1144 ( .a ({signal_2443, signal_985}), .b ({signal_2415, signal_957}), .clk ( clk ), .r ( Fresh[154] ), .c ({signal_2617, signal_1159}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1145 ( .a ({signal_2449, signal_991}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[155] ), .c ({signal_2618, signal_1160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1146 ( .a ({signal_2410, signal_952}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[156] ), .c ({signal_2619, signal_1161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1147 ( .a ({signal_2443, signal_985}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[157] ), .c ({signal_2620, signal_1162}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1148 ( .a ({signal_2424, signal_966}), .b ({signal_2431, signal_973}), .clk ( clk ), .r ( Fresh[158] ), .c ({signal_2621, signal_1163}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1149 ( .a ({signal_2446, signal_988}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[159] ), .c ({signal_2622, signal_1164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1150 ( .a ({signal_2450, signal_992}), .b ({signal_2469, signal_1011}), .clk ( clk ), .r ( Fresh[160] ), .c ({signal_2623, signal_1165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1151 ( .a ({signal_2440, signal_982}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[161] ), .c ({signal_2624, signal_1166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1152 ( .a ({signal_2438, signal_980}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[162] ), .c ({signal_2625, signal_1167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1153 ( .a ({signal_4788, signal_4786}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[163] ), .c ({signal_2626, signal_1168}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1154 ( .a ({signal_2415, signal_957}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[164] ), .c ({signal_2627, signal_1169}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1156 ( .a ({signal_2464, signal_1006}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[165] ), .c ({signal_2629, signal_1171}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1157 ( .a ({signal_2442, signal_984}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[166] ), .c ({signal_2630, signal_1172}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1158 ( .a ({signal_2455, signal_997}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[167] ), .c ({signal_2631, signal_1173}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1159 ( .a ({signal_2449, signal_991}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[168] ), .c ({signal_2632, signal_1174}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1160 ( .a ({signal_4776, signal_4774}), .b ({signal_2446, signal_988}), .clk ( clk ), .r ( Fresh[169] ), .c ({signal_2633, signal_1175}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1161 ( .a ({signal_4768, signal_4766}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[170] ), .c ({signal_2634, signal_1176}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1162 ( .a ({signal_4764, signal_4762}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[171] ), .c ({signal_2635, signal_1177}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1163 ( .a ({signal_2453, signal_995}), .b ({signal_2473, signal_1015}), .clk ( clk ), .r ( Fresh[172] ), .c ({signal_2636, signal_1178}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1164 ( .a ({signal_2424, signal_966}), .b ({signal_2430, signal_972}), .clk ( clk ), .r ( Fresh[173] ), .c ({signal_2637, signal_1179}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1165 ( .a ({signal_2429, signal_971}), .b ({signal_2430, signal_972}), .clk ( clk ), .r ( Fresh[174] ), .c ({signal_2638, signal_1180}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1166 ( .a ({signal_2420, signal_962}), .b ({signal_2470, signal_1012}), .clk ( clk ), .r ( Fresh[175] ), .c ({signal_2639, signal_1181}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1167 ( .a ({signal_2438, signal_980}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[176] ), .c ({signal_2640, signal_1182}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1168 ( .a ({signal_2413, signal_955}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[177] ), .c ({signal_2641, signal_1183}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1169 ( .a ({signal_4760, signal_4758}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[178] ), .c ({signal_2642, signal_1184}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1170 ( .a ({signal_2444, signal_986}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[179] ), .c ({signal_2643, signal_1185}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1171 ( .a ({signal_2420, signal_962}), .b ({signal_2473, signal_1015}), .clk ( clk ), .r ( Fresh[180] ), .c ({signal_2644, signal_1186}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1172 ( .a ({signal_2446, signal_988}), .b ({signal_2453, signal_995}), .clk ( clk ), .r ( Fresh[181] ), .c ({signal_2645, signal_1187}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1174 ( .a ({signal_2441, signal_983}), .b ({signal_2442, signal_984}), .clk ( clk ), .r ( Fresh[182] ), .c ({signal_2647, signal_1189}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1175 ( .a ({signal_2441, signal_983}), .b ({signal_2462, signal_1004}), .clk ( clk ), .r ( Fresh[183] ), .c ({signal_2648, signal_1190}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1176 ( .a ({signal_2409, signal_951}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[184] ), .c ({signal_2649, signal_1191}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1177 ( .a ({signal_2454, signal_996}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[185] ), .c ({signal_2650, signal_1192}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1178 ( .a ({signal_2427, signal_969}), .b ({signal_2434, signal_976}), .clk ( clk ), .r ( Fresh[186] ), .c ({signal_2651, signal_1193}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1179 ( .a ({signal_2411, signal_953}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[187] ), .c ({signal_2652, signal_1194}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1180 ( .a ({signal_2445, signal_987}), .b ({signal_2415, signal_957}), .clk ( clk ), .r ( Fresh[188] ), .c ({signal_2653, signal_1195}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1181 ( .a ({signal_2420, signal_962}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[189] ), .c ({signal_2654, signal_1196}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1182 ( .a ({signal_4772, signal_4770}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[190] ), .c ({signal_2655, signal_1197}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1183 ( .a ({signal_2438, signal_980}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[191] ), .c ({signal_2656, signal_1198}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1185 ( .a ({signal_2442, signal_984}), .b ({signal_2473, signal_1015}), .clk ( clk ), .r ( Fresh[192] ), .c ({signal_2658, signal_1200}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1186 ( .a ({signal_2456, signal_998}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[193] ), .c ({signal_2659, signal_1201}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1187 ( .a ({signal_4788, signal_4786}), .b ({signal_2443, signal_985}), .clk ( clk ), .r ( Fresh[194] ), .c ({signal_2660, signal_1202}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1188 ( .a ({signal_2444, signal_986}), .b ({signal_2417, signal_959}), .clk ( clk ), .r ( Fresh[195] ), .c ({signal_2661, signal_1203}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1191 ( .a ({signal_2439, signal_981}), .b ({signal_2445, signal_987}), .clk ( clk ), .r ( Fresh[196] ), .c ({signal_2664, signal_1206}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1192 ( .a ({signal_2456, signal_998}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[197] ), .c ({signal_2665, signal_1207}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1193 ( .a ({signal_2415, signal_957}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[198] ), .c ({signal_2666, signal_1208}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1194 ( .a ({signal_2444, signal_986}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[199] ), .c ({signal_2667, signal_1209}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1195 ( .a ({signal_2446, signal_988}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[200] ), .c ({signal_2668, signal_1210}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1196 ( .a ({signal_2447, signal_989}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[201] ), .c ({signal_2669, signal_1211}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1197 ( .a ({signal_2443, signal_985}), .b ({signal_2444, signal_986}), .clk ( clk ), .r ( Fresh[202] ), .c ({signal_2670, signal_1212}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1199 ( .a ({signal_2449, signal_991}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[203] ), .c ({signal_2672, signal_1214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1200 ( .a ({signal_2411, signal_953}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[204] ), .c ({signal_2673, signal_1215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1201 ( .a ({signal_2451, signal_993}), .b ({signal_2456, signal_998}), .clk ( clk ), .r ( Fresh[205] ), .c ({signal_2674, signal_1216}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1202 ( .a ({signal_2446, signal_988}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[206] ), .c ({signal_2675, signal_1217}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1203 ( .a ({signal_2453, signal_995}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[207] ), .c ({signal_2676, signal_1218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1204 ( .a ({signal_2437, signal_979}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[208] ), .c ({signal_2677, signal_1219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1205 ( .a ({signal_4780, signal_4778}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[209] ), .c ({signal_2678, signal_1220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1206 ( .a ({signal_4760, signal_4758}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[210] ), .c ({signal_2679, signal_1221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1208 ( .a ({signal_2462, signal_1004}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[211] ), .c ({signal_2681, signal_1223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1210 ( .a ({signal_4784, signal_4782}), .b ({signal_2428, signal_970}), .clk ( clk ), .r ( Fresh[212] ), .c ({signal_2683, signal_1225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1213 ( .a ({signal_2437, signal_979}), .b ({signal_4792, signal_4790}), .clk ( clk ), .r ( Fresh[213] ), .c ({signal_2686, signal_1228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1214 ( .a ({signal_4784, signal_4782}), .b ({signal_2430, signal_972}), .clk ( clk ), .r ( Fresh[214] ), .c ({signal_2687, signal_1229}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1215 ( .a ({signal_2527, signal_1069}), .b ({signal_2688, signal_1230}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1216 ( .a ({signal_2528, signal_1070}), .b ({signal_2689, signal_1231}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1217 ( .a ({signal_2530, signal_1072}), .b ({signal_2690, signal_1232}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1218 ( .a ({signal_2531, signal_1073}), .b ({signal_2691, signal_1233}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1219 ( .a ({signal_2532, signal_1074}), .b ({signal_2692, signal_1234}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1220 ( .a ({signal_2533, signal_1075}), .b ({signal_2693, signal_1235}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1221 ( .a ({signal_2534, signal_1076}), .b ({signal_2694, signal_1236}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1222 ( .a ({signal_2535, signal_1077}), .b ({signal_2695, signal_1237}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1223 ( .a ({signal_2536, signal_1078}), .b ({signal_2696, signal_1238}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1224 ( .a ({signal_2537, signal_1079}), .b ({signal_2697, signal_1239}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1225 ( .a ({signal_2538, signal_1080}), .b ({signal_2698, signal_1240}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1226 ( .a ({signal_2539, signal_1081}), .b ({signal_2699, signal_1241}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1227 ( .a ({signal_2540, signal_1082}), .b ({signal_2700, signal_1242}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1228 ( .a ({signal_2541, signal_1083}), .b ({signal_2701, signal_1243}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1229 ( .a ({signal_2542, signal_1084}), .b ({signal_2702, signal_1244}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1230 ( .a ({signal_2544, signal_1086}), .b ({signal_2703, signal_1245}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1231 ( .a ({signal_2545, signal_1087}), .b ({signal_2704, signal_1246}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1232 ( .a ({signal_2546, signal_1088}), .b ({signal_2705, signal_1247}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1233 ( .a ({signal_2548, signal_1090}), .b ({signal_2706, signal_1248}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1234 ( .a ({signal_2549, signal_1091}), .b ({signal_2707, signal_1249}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1235 ( .a ({signal_2550, signal_1092}), .b ({signal_2708, signal_1250}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1236 ( .a ({signal_2551, signal_1093}), .b ({signal_2709, signal_1251}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1237 ( .a ({signal_2552, signal_1094}), .b ({signal_2710, signal_1252}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1238 ( .a ({signal_2553, signal_1095}), .b ({signal_2711, signal_1253}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1239 ( .a ({signal_2554, signal_1096}), .b ({signal_2712, signal_1254}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1240 ( .a ({signal_2555, signal_1097}), .b ({signal_2713, signal_1255}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1241 ( .a ({signal_2556, signal_1098}), .b ({signal_2714, signal_1256}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1242 ( .a ({signal_2557, signal_1099}), .b ({signal_2715, signal_1257}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1244 ( .a ({signal_2559, signal_1101}), .b ({signal_2717, signal_1259}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1245 ( .a ({signal_2561, signal_1103}), .b ({signal_2718, signal_1260}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1246 ( .a ({signal_2563, signal_1105}), .b ({signal_2719, signal_1261}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1247 ( .a ({signal_2564, signal_1106}), .b ({signal_2720, signal_1262}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1248 ( .a ({signal_2566, signal_1108}), .b ({signal_2721, signal_1263}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1249 ( .a ({signal_2567, signal_1109}), .b ({signal_2722, signal_1264}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1250 ( .a ({signal_2568, signal_1110}), .b ({signal_2723, signal_1265}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1251 ( .a ({signal_2569, signal_1111}), .b ({signal_2724, signal_1266}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1252 ( .a ({signal_2570, signal_1112}), .b ({signal_2725, signal_1267}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1253 ( .a ({signal_2571, signal_1113}), .b ({signal_2726, signal_1268}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1254 ( .a ({signal_2573, signal_1115}), .b ({signal_2727, signal_1269}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1255 ( .a ({signal_2574, signal_1116}), .b ({signal_2728, signal_1270}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1256 ( .a ({signal_2575, signal_1117}), .b ({signal_2729, signal_1271}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1257 ( .a ({signal_2576, signal_1118}), .b ({signal_2730, signal_1272}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1258 ( .a ({signal_2578, signal_1120}), .b ({signal_2731, signal_1273}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1259 ( .a ({signal_2579, signal_1121}), .b ({signal_2732, signal_1274}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1260 ( .a ({signal_2580, signal_1122}), .b ({signal_2733, signal_1275}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1261 ( .a ({signal_2582, signal_1124}), .b ({signal_2734, signal_1276}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1262 ( .a ({signal_2583, signal_1125}), .b ({signal_2735, signal_1277}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1263 ( .a ({signal_2584, signal_1126}), .b ({signal_2736, signal_1278}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1264 ( .a ({signal_2585, signal_1127}), .b ({signal_2737, signal_1279}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1265 ( .a ({signal_2587, signal_1129}), .b ({signal_2738, signal_1280}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1266 ( .a ({signal_2588, signal_1130}), .b ({signal_2739, signal_1281}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1267 ( .a ({signal_2589, signal_1131}), .b ({signal_2740, signal_1282}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1268 ( .a ({signal_2592, signal_1134}), .b ({signal_2741, signal_1283}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1269 ( .a ({signal_2593, signal_1135}), .b ({signal_2742, signal_1284}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1270 ( .a ({signal_2594, signal_1136}), .b ({signal_2743, signal_1285}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1271 ( .a ({signal_2595, signal_1137}), .b ({signal_2744, signal_1286}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1273 ( .a ({signal_2599, signal_1141}), .b ({signal_2746, signal_1288}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1274 ( .a ({signal_2601, signal_1143}), .b ({signal_2747, signal_1289}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1275 ( .a ({signal_2602, signal_1144}), .b ({signal_2748, signal_1290}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1276 ( .a ({signal_2604, signal_1146}), .b ({signal_2749, signal_1291}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1278 ( .a ({signal_2606, signal_1148}), .b ({signal_2751, signal_1293}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1279 ( .a ({signal_2607, signal_1149}), .b ({signal_2752, signal_1294}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1280 ( .a ({signal_2608, signal_1150}), .b ({signal_2753, signal_1295}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1281 ( .a ({signal_2610, signal_1152}), .b ({signal_2754, signal_1296}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1282 ( .a ({signal_2611, signal_1153}), .b ({signal_2755, signal_1297}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1283 ( .a ({signal_2612, signal_1154}), .b ({signal_2756, signal_1298}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1285 ( .a ({signal_2614, signal_1156}), .b ({signal_2758, signal_1300}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1286 ( .a ({signal_2615, signal_1157}), .b ({signal_2759, signal_1301}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1287 ( .a ({signal_2617, signal_1159}), .b ({signal_2760, signal_1302}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1288 ( .a ({signal_2618, signal_1160}), .b ({signal_2761, signal_1303}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1289 ( .a ({signal_2619, signal_1161}), .b ({signal_2762, signal_1304}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1290 ( .a ({signal_2620, signal_1162}), .b ({signal_2763, signal_1305}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1291 ( .a ({signal_2621, signal_1163}), .b ({signal_2764, signal_1306}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1292 ( .a ({signal_2622, signal_1164}), .b ({signal_2765, signal_1307}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1293 ( .a ({signal_2623, signal_1165}), .b ({signal_2766, signal_1308}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1294 ( .a ({signal_2624, signal_1166}), .b ({signal_2767, signal_1309}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1295 ( .a ({signal_2625, signal_1167}), .b ({signal_2768, signal_1310}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1296 ( .a ({signal_2627, signal_1169}), .b ({signal_2769, signal_1311}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1298 ( .a ({signal_2629, signal_1171}), .b ({signal_2771, signal_1313}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1299 ( .a ({signal_2630, signal_1172}), .b ({signal_2772, signal_1314}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1300 ( .a ({signal_2631, signal_1173}), .b ({signal_2773, signal_1315}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1301 ( .a ({signal_2632, signal_1174}), .b ({signal_2774, signal_1316}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1302 ( .a ({signal_2633, signal_1175}), .b ({signal_2775, signal_1317}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1303 ( .a ({signal_2634, signal_1176}), .b ({signal_2776, signal_1318}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1304 ( .a ({signal_2635, signal_1177}), .b ({signal_2777, signal_1319}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1305 ( .a ({signal_2637, signal_1179}), .b ({signal_2778, signal_1320}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1306 ( .a ({signal_2638, signal_1180}), .b ({signal_2779, signal_1321}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1307 ( .a ({signal_2639, signal_1181}), .b ({signal_2780, signal_1322}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1308 ( .a ({signal_2640, signal_1182}), .b ({signal_2781, signal_1323}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1309 ( .a ({signal_2641, signal_1183}), .b ({signal_2782, signal_1324}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1310 ( .a ({signal_2642, signal_1184}), .b ({signal_2783, signal_1325}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1311 ( .a ({signal_2643, signal_1185}), .b ({signal_2784, signal_1326}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1312 ( .a ({signal_2644, signal_1186}), .b ({signal_2785, signal_1327}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1313 ( .a ({signal_2645, signal_1187}), .b ({signal_2786, signal_1328}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1315 ( .a ({signal_2647, signal_1189}), .b ({signal_2788, signal_1330}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1316 ( .a ({signal_2649, signal_1191}), .b ({signal_2789, signal_1331}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1317 ( .a ({signal_2650, signal_1192}), .b ({signal_2790, signal_1332}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1318 ( .a ({signal_2651, signal_1193}), .b ({signal_2791, signal_1333}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1319 ( .a ({signal_2652, signal_1194}), .b ({signal_2792, signal_1334}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1320 ( .a ({signal_2653, signal_1195}), .b ({signal_2793, signal_1335}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1321 ( .a ({signal_2654, signal_1196}), .b ({signal_2794, signal_1336}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1322 ( .a ({signal_2655, signal_1197}), .b ({signal_2795, signal_1337}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1324 ( .a ({signal_2658, signal_1200}), .b ({signal_2797, signal_1339}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1325 ( .a ({signal_2659, signal_1201}), .b ({signal_2798, signal_1340}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1326 ( .a ({signal_2660, signal_1202}), .b ({signal_2799, signal_1341}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1327 ( .a ({signal_2661, signal_1203}), .b ({signal_2800, signal_1342}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1330 ( .a ({signal_2665, signal_1207}), .b ({signal_2803, signal_1345}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1331 ( .a ({signal_2667, signal_1209}), .b ({signal_2804, signal_1346}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1332 ( .a ({signal_2668, signal_1210}), .b ({signal_2805, signal_1347}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1333 ( .a ({signal_2669, signal_1211}), .b ({signal_2806, signal_1348}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1334 ( .a ({signal_2670, signal_1212}), .b ({signal_2807, signal_1349}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1336 ( .a ({signal_2672, signal_1214}), .b ({signal_2809, signal_1351}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1337 ( .a ({signal_2673, signal_1215}), .b ({signal_2810, signal_1352}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1338 ( .a ({signal_2674, signal_1216}), .b ({signal_2811, signal_1353}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1339 ( .a ({signal_2676, signal_1218}), .b ({signal_2812, signal_1354}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1340 ( .a ({signal_2677, signal_1219}), .b ({signal_2813, signal_1355}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1341 ( .a ({signal_2678, signal_1220}), .b ({signal_2814, signal_1356}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1342 ( .a ({signal_2679, signal_1221}), .b ({signal_2815, signal_1357}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1344 ( .a ({signal_2681, signal_1223}), .b ({signal_2817, signal_1359}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1346 ( .a ({signal_2683, signal_1225}), .b ({signal_2819, signal_1361}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1349 ( .a ({signal_2686, signal_1228}), .b ({signal_2822, signal_1364}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1350 ( .a ({signal_2687, signal_1229}), .b ({signal_2823, signal_1365}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1353 ( .a ({signal_4796, signal_4794}), .b ({signal_2504, signal_1046}), .clk ( clk ), .r ( Fresh[215] ), .c ({signal_2826, signal_1368}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1354 ( .a ({signal_4776, signal_4774}), .b ({signal_2500, signal_1042}), .clk ( clk ), .r ( Fresh[216] ), .c ({signal_2827, signal_1369}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1355 ( .a ({signal_2489, signal_1031}), .b ({signal_2516, signal_1058}), .clk ( clk ), .r ( Fresh[217] ), .c ({signal_2828, signal_1370}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1356 ( .a ({signal_2503, signal_1045}), .b ({signal_2515, signal_1057}), .clk ( clk ), .r ( Fresh[218] ), .c ({signal_2829, signal_1371}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1357 ( .a ({signal_2494, signal_1036}), .b ({signal_2495, signal_1037}), .clk ( clk ), .r ( Fresh[219] ), .c ({signal_2830, signal_1372}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1360 ( .a ({signal_2494, signal_1036}), .b ({signal_2503, signal_1045}), .clk ( clk ), .r ( Fresh[220] ), .c ({signal_2833, signal_1375}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1361 ( .a ({signal_2499, signal_1041}), .b ({signal_2510, signal_1052}), .clk ( clk ), .r ( Fresh[221] ), .c ({signal_2834, signal_1376}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1362 ( .a ({signal_2509, signal_1051}), .b ({signal_2511, signal_1053}), .clk ( clk ), .r ( Fresh[222] ), .c ({signal_2835, signal_1377}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1365 ( .a ({signal_2489, signal_1031}), .b ({signal_2502, signal_1044}), .clk ( clk ), .r ( Fresh[223] ), .c ({signal_2838, signal_1380}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1366 ( .a ({signal_2490, signal_1032}), .b ({signal_2510, signal_1052}), .clk ( clk ), .r ( Fresh[224] ), .c ({signal_2839, signal_1381}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1367 ( .a ({signal_2500, signal_1042}), .b ({signal_2501, signal_1043}), .clk ( clk ), .r ( Fresh[225] ), .c ({signal_2840, signal_1382}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1368 ( .a ({signal_2495, signal_1037}), .b ({signal_2503, signal_1045}), .clk ( clk ), .r ( Fresh[226] ), .c ({signal_2841, signal_1383}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1369 ( .a ({signal_2432, signal_974}), .b ({signal_2511, signal_1053}), .clk ( clk ), .r ( Fresh[227] ), .c ({signal_2842, signal_1384}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1375 ( .a ({signal_2498, signal_1040}), .b ({signal_2514, signal_1056}), .clk ( clk ), .r ( Fresh[228] ), .c ({signal_2848, signal_1390}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1376 ( .a ({signal_2503, signal_1045}), .b ({signal_2508, signal_1050}), .clk ( clk ), .r ( Fresh[229] ), .c ({signal_2849, signal_1391}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1383 ( .a ({signal_2491, signal_1033}), .b ({signal_2493, signal_1035}), .clk ( clk ), .r ( Fresh[230] ), .c ({signal_2856, signal_1398}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1395 ( .a ({signal_2429, signal_971}), .b ({signal_2507, signal_1049}), .clk ( clk ), .r ( Fresh[231] ), .c ({signal_2868, signal_1410}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1396 ( .a ({signal_2490, signal_1032}), .b ({signal_2505, signal_1047}), .clk ( clk ), .r ( Fresh[232] ), .c ({signal_2869, signal_1411}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1401 ( .a ({signal_2425, signal_967}), .b ({signal_2501, signal_1043}), .clk ( clk ), .r ( Fresh[233] ), .c ({signal_2874, signal_1416}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1402 ( .a ({signal_2508, signal_1050}), .b ({signal_2433, signal_975}), .clk ( clk ), .r ( Fresh[234] ), .c ({signal_2875, signal_1417}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1403 ( .a ({signal_2430, signal_972}), .b ({signal_2503, signal_1045}), .clk ( clk ), .r ( Fresh[235] ), .c ({signal_2876, signal_1418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1407 ( .a ({signal_2496, signal_1038}), .b ({signal_2504, signal_1046}), .clk ( clk ), .r ( Fresh[236] ), .c ({signal_2880, signal_1422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1408 ( .a ({signal_2498, signal_1040}), .b ({signal_2433, signal_975}), .clk ( clk ), .r ( Fresh[237] ), .c ({signal_2881, signal_1423}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1492 ( .a ({signal_2826, signal_1368}), .b ({signal_2965, signal_1507}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1493 ( .a ({signal_2827, signal_1369}), .b ({signal_2966, signal_1508}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1494 ( .a ({signal_2828, signal_1370}), .b ({signal_2967, signal_1509}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1495 ( .a ({signal_2829, signal_1371}), .b ({signal_2968, signal_1510}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1496 ( .a ({signal_2830, signal_1372}), .b ({signal_2969, signal_1511}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1499 ( .a ({signal_2833, signal_1375}), .b ({signal_2972, signal_1514}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1500 ( .a ({signal_2834, signal_1376}), .b ({signal_2973, signal_1515}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1501 ( .a ({signal_2835, signal_1377}), .b ({signal_2974, signal_1516}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1504 ( .a ({signal_2838, signal_1380}), .b ({signal_2977, signal_1519}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1505 ( .a ({signal_2839, signal_1381}), .b ({signal_2978, signal_1520}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1506 ( .a ({signal_2840, signal_1382}), .b ({signal_2979, signal_1521}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1507 ( .a ({signal_2842, signal_1384}), .b ({signal_2980, signal_1522}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1513 ( .a ({signal_2849, signal_1391}), .b ({signal_2986, signal_1528}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1520 ( .a ({signal_2856, signal_1398}), .b ({signal_2993, signal_1535}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1532 ( .a ({signal_2868, signal_1410}), .b ({signal_3005, signal_1547}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1533 ( .a ({signal_2869, signal_1411}), .b ({signal_3006, signal_1548}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1538 ( .a ({signal_2874, signal_1416}), .b ({signal_3011, signal_1553}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1539 ( .a ({signal_2875, signal_1417}), .b ({signal_3012, signal_1554}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1543 ( .a ({signal_2880, signal_1422}), .b ({signal_3016, signal_1558}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1544 ( .a ({signal_2881, signal_1423}), .b ({signal_3017, signal_1559}) ) ;
    buf_clk cell_2440 ( .C ( clk ), .D ( signal_4799 ), .Q ( signal_4800 ) ) ;
    buf_clk cell_2444 ( .C ( clk ), .D ( signal_4803 ), .Q ( signal_4804 ) ) ;
    buf_clk cell_2446 ( .C ( clk ), .D ( signal_4805 ), .Q ( signal_4806 ) ) ;
    buf_clk cell_2448 ( .C ( clk ), .D ( signal_4807 ), .Q ( signal_4808 ) ) ;
    buf_clk cell_2450 ( .C ( clk ), .D ( signal_4809 ), .Q ( signal_4810 ) ) ;
    buf_clk cell_2452 ( .C ( clk ), .D ( signal_4811 ), .Q ( signal_4812 ) ) ;
    buf_clk cell_2454 ( .C ( clk ), .D ( signal_4813 ), .Q ( signal_4814 ) ) ;
    buf_clk cell_2456 ( .C ( clk ), .D ( signal_4815 ), .Q ( signal_4816 ) ) ;
    buf_clk cell_2458 ( .C ( clk ), .D ( signal_4817 ), .Q ( signal_4818 ) ) ;
    buf_clk cell_2460 ( .C ( clk ), .D ( signal_4819 ), .Q ( signal_4820 ) ) ;
    buf_clk cell_2462 ( .C ( clk ), .D ( signal_4821 ), .Q ( signal_4822 ) ) ;
    buf_clk cell_2464 ( .C ( clk ), .D ( signal_4823 ), .Q ( signal_4824 ) ) ;
    buf_clk cell_2466 ( .C ( clk ), .D ( signal_4825 ), .Q ( signal_4826 ) ) ;
    buf_clk cell_2468 ( .C ( clk ), .D ( signal_4827 ), .Q ( signal_4828 ) ) ;
    buf_clk cell_2470 ( .C ( clk ), .D ( signal_4829 ), .Q ( signal_4830 ) ) ;
    buf_clk cell_2472 ( .C ( clk ), .D ( signal_4831 ), .Q ( signal_4832 ) ) ;
    buf_clk cell_2474 ( .C ( clk ), .D ( signal_4833 ), .Q ( signal_4834 ) ) ;
    buf_clk cell_2476 ( .C ( clk ), .D ( signal_4835 ), .Q ( signal_4836 ) ) ;
    buf_clk cell_2478 ( .C ( clk ), .D ( signal_4837 ), .Q ( signal_4838 ) ) ;
    buf_clk cell_2480 ( .C ( clk ), .D ( signal_4839 ), .Q ( signal_4840 ) ) ;
    buf_clk cell_2482 ( .C ( clk ), .D ( signal_4841 ), .Q ( signal_4842 ) ) ;
    buf_clk cell_2484 ( .C ( clk ), .D ( signal_4843 ), .Q ( signal_4844 ) ) ;
    buf_clk cell_2486 ( .C ( clk ), .D ( signal_4845 ), .Q ( signal_4846 ) ) ;
    buf_clk cell_2488 ( .C ( clk ), .D ( signal_4847 ), .Q ( signal_4848 ) ) ;
    buf_clk cell_2490 ( .C ( clk ), .D ( signal_4849 ), .Q ( signal_4850 ) ) ;
    buf_clk cell_2492 ( .C ( clk ), .D ( signal_4851 ), .Q ( signal_4852 ) ) ;
    buf_clk cell_2494 ( .C ( clk ), .D ( signal_4853 ), .Q ( signal_4854 ) ) ;
    buf_clk cell_2496 ( .C ( clk ), .D ( signal_4855 ), .Q ( signal_4856 ) ) ;
    buf_clk cell_2498 ( .C ( clk ), .D ( signal_4857 ), .Q ( signal_4858 ) ) ;
    buf_clk cell_2500 ( .C ( clk ), .D ( signal_4859 ), .Q ( signal_4860 ) ) ;
    buf_clk cell_2502 ( .C ( clk ), .D ( signal_4861 ), .Q ( signal_4862 ) ) ;
    buf_clk cell_2504 ( .C ( clk ), .D ( signal_4863 ), .Q ( signal_4864 ) ) ;
    buf_clk cell_2506 ( .C ( clk ), .D ( signal_4865 ), .Q ( signal_4866 ) ) ;
    buf_clk cell_2508 ( .C ( clk ), .D ( signal_4867 ), .Q ( signal_4868 ) ) ;
    buf_clk cell_2510 ( .C ( clk ), .D ( signal_4869 ), .Q ( signal_4870 ) ) ;
    buf_clk cell_2512 ( .C ( clk ), .D ( signal_4871 ), .Q ( signal_4872 ) ) ;
    buf_clk cell_2514 ( .C ( clk ), .D ( signal_4873 ), .Q ( signal_4874 ) ) ;
    buf_clk cell_2516 ( .C ( clk ), .D ( signal_4875 ), .Q ( signal_4876 ) ) ;
    buf_clk cell_2518 ( .C ( clk ), .D ( signal_4877 ), .Q ( signal_4878 ) ) ;
    buf_clk cell_2520 ( .C ( clk ), .D ( signal_4879 ), .Q ( signal_4880 ) ) ;
    buf_clk cell_2522 ( .C ( clk ), .D ( signal_4881 ), .Q ( signal_4882 ) ) ;
    buf_clk cell_2524 ( .C ( clk ), .D ( signal_4883 ), .Q ( signal_4884 ) ) ;
    buf_clk cell_2526 ( .C ( clk ), .D ( signal_4885 ), .Q ( signal_4886 ) ) ;
    buf_clk cell_2528 ( .C ( clk ), .D ( signal_4887 ), .Q ( signal_4888 ) ) ;
    buf_clk cell_2530 ( .C ( clk ), .D ( signal_4889 ), .Q ( signal_4890 ) ) ;
    buf_clk cell_2532 ( .C ( clk ), .D ( signal_4891 ), .Q ( signal_4892 ) ) ;
    buf_clk cell_2534 ( .C ( clk ), .D ( signal_4893 ), .Q ( signal_4894 ) ) ;
    buf_clk cell_2536 ( .C ( clk ), .D ( signal_4895 ), .Q ( signal_4896 ) ) ;
    buf_clk cell_2538 ( .C ( clk ), .D ( signal_4897 ), .Q ( signal_4898 ) ) ;
    buf_clk cell_2540 ( .C ( clk ), .D ( signal_4899 ), .Q ( signal_4900 ) ) ;
    buf_clk cell_2542 ( .C ( clk ), .D ( signal_4901 ), .Q ( signal_4902 ) ) ;
    buf_clk cell_2544 ( .C ( clk ), .D ( signal_4903 ), .Q ( signal_4904 ) ) ;
    buf_clk cell_2546 ( .C ( clk ), .D ( signal_4905 ), .Q ( signal_4906 ) ) ;
    buf_clk cell_2548 ( .C ( clk ), .D ( signal_4907 ), .Q ( signal_4908 ) ) ;
    buf_clk cell_2550 ( .C ( clk ), .D ( signal_4909 ), .Q ( signal_4910 ) ) ;
    buf_clk cell_2552 ( .C ( clk ), .D ( signal_4911 ), .Q ( signal_4912 ) ) ;
    buf_clk cell_2554 ( .C ( clk ), .D ( signal_4913 ), .Q ( signal_4914 ) ) ;
    buf_clk cell_2556 ( .C ( clk ), .D ( signal_4915 ), .Q ( signal_4916 ) ) ;
    buf_clk cell_2558 ( .C ( clk ), .D ( signal_4917 ), .Q ( signal_4918 ) ) ;
    buf_clk cell_2560 ( .C ( clk ), .D ( signal_4919 ), .Q ( signal_4920 ) ) ;
    buf_clk cell_2562 ( .C ( clk ), .D ( signal_4921 ), .Q ( signal_4922 ) ) ;
    buf_clk cell_2564 ( .C ( clk ), .D ( signal_4923 ), .Q ( signal_4924 ) ) ;
    buf_clk cell_2566 ( .C ( clk ), .D ( signal_4925 ), .Q ( signal_4926 ) ) ;
    buf_clk cell_2568 ( .C ( clk ), .D ( signal_4927 ), .Q ( signal_4928 ) ) ;
    buf_clk cell_2570 ( .C ( clk ), .D ( signal_4929 ), .Q ( signal_4930 ) ) ;
    buf_clk cell_2572 ( .C ( clk ), .D ( signal_4931 ), .Q ( signal_4932 ) ) ;
    buf_clk cell_2574 ( .C ( clk ), .D ( signal_4933 ), .Q ( signal_4934 ) ) ;
    buf_clk cell_2576 ( .C ( clk ), .D ( signal_4935 ), .Q ( signal_4936 ) ) ;
    buf_clk cell_2578 ( .C ( clk ), .D ( signal_4937 ), .Q ( signal_4938 ) ) ;
    buf_clk cell_2580 ( .C ( clk ), .D ( signal_4939 ), .Q ( signal_4940 ) ) ;
    buf_clk cell_2584 ( .C ( clk ), .D ( signal_4943 ), .Q ( signal_4944 ) ) ;
    buf_clk cell_2588 ( .C ( clk ), .D ( signal_4947 ), .Q ( signal_4948 ) ) ;
    buf_clk cell_2590 ( .C ( clk ), .D ( signal_4949 ), .Q ( signal_4950 ) ) ;
    buf_clk cell_2592 ( .C ( clk ), .D ( signal_4951 ), .Q ( signal_4952 ) ) ;
    buf_clk cell_2594 ( .C ( clk ), .D ( signal_4953 ), .Q ( signal_4954 ) ) ;
    buf_clk cell_2596 ( .C ( clk ), .D ( signal_4955 ), .Q ( signal_4956 ) ) ;
    buf_clk cell_2598 ( .C ( clk ), .D ( signal_4957 ), .Q ( signal_4958 ) ) ;
    buf_clk cell_2600 ( .C ( clk ), .D ( signal_4959 ), .Q ( signal_4960 ) ) ;
    buf_clk cell_2602 ( .C ( clk ), .D ( signal_4961 ), .Q ( signal_4962 ) ) ;
    buf_clk cell_2604 ( .C ( clk ), .D ( signal_4963 ), .Q ( signal_4964 ) ) ;
    buf_clk cell_2606 ( .C ( clk ), .D ( signal_4965 ), .Q ( signal_4966 ) ) ;
    buf_clk cell_2608 ( .C ( clk ), .D ( signal_4967 ), .Q ( signal_4968 ) ) ;
    buf_clk cell_2610 ( .C ( clk ), .D ( signal_4969 ), .Q ( signal_4970 ) ) ;
    buf_clk cell_2612 ( .C ( clk ), .D ( signal_4971 ), .Q ( signal_4972 ) ) ;
    buf_clk cell_2614 ( .C ( clk ), .D ( signal_4973 ), .Q ( signal_4974 ) ) ;
    buf_clk cell_2616 ( .C ( clk ), .D ( signal_4975 ), .Q ( signal_4976 ) ) ;
    buf_clk cell_2618 ( .C ( clk ), .D ( signal_4977 ), .Q ( signal_4978 ) ) ;
    buf_clk cell_2620 ( .C ( clk ), .D ( signal_4979 ), .Q ( signal_4980 ) ) ;
    buf_clk cell_2622 ( .C ( clk ), .D ( signal_4981 ), .Q ( signal_4982 ) ) ;
    buf_clk cell_2624 ( .C ( clk ), .D ( signal_4983 ), .Q ( signal_4984 ) ) ;
    buf_clk cell_2626 ( .C ( clk ), .D ( signal_4985 ), .Q ( signal_4986 ) ) ;
    buf_clk cell_2628 ( .C ( clk ), .D ( signal_4987 ), .Q ( signal_4988 ) ) ;
    buf_clk cell_2630 ( .C ( clk ), .D ( signal_4989 ), .Q ( signal_4990 ) ) ;
    buf_clk cell_2632 ( .C ( clk ), .D ( signal_4991 ), .Q ( signal_4992 ) ) ;
    buf_clk cell_2634 ( .C ( clk ), .D ( signal_4993 ), .Q ( signal_4994 ) ) ;
    buf_clk cell_2636 ( .C ( clk ), .D ( signal_4995 ), .Q ( signal_4996 ) ) ;
    buf_clk cell_2638 ( .C ( clk ), .D ( signal_4997 ), .Q ( signal_4998 ) ) ;
    buf_clk cell_2640 ( .C ( clk ), .D ( signal_4999 ), .Q ( signal_5000 ) ) ;
    buf_clk cell_2642 ( .C ( clk ), .D ( signal_5001 ), .Q ( signal_5002 ) ) ;
    buf_clk cell_2644 ( .C ( clk ), .D ( signal_5003 ), .Q ( signal_5004 ) ) ;
    buf_clk cell_2646 ( .C ( clk ), .D ( signal_5005 ), .Q ( signal_5006 ) ) ;
    buf_clk cell_2648 ( .C ( clk ), .D ( signal_5007 ), .Q ( signal_5008 ) ) ;
    buf_clk cell_2650 ( .C ( clk ), .D ( signal_5009 ), .Q ( signal_5010 ) ) ;
    buf_clk cell_2652 ( .C ( clk ), .D ( signal_5011 ), .Q ( signal_5012 ) ) ;
    buf_clk cell_2654 ( .C ( clk ), .D ( signal_5013 ), .Q ( signal_5014 ) ) ;
    buf_clk cell_2656 ( .C ( clk ), .D ( signal_5015 ), .Q ( signal_5016 ) ) ;
    buf_clk cell_2658 ( .C ( clk ), .D ( signal_5017 ), .Q ( signal_5018 ) ) ;
    buf_clk cell_2660 ( .C ( clk ), .D ( signal_5019 ), .Q ( signal_5020 ) ) ;
    buf_clk cell_2662 ( .C ( clk ), .D ( signal_5021 ), .Q ( signal_5022 ) ) ;
    buf_clk cell_2664 ( .C ( clk ), .D ( signal_5023 ), .Q ( signal_5024 ) ) ;
    buf_clk cell_2666 ( .C ( clk ), .D ( signal_5025 ), .Q ( signal_5026 ) ) ;
    buf_clk cell_2668 ( .C ( clk ), .D ( signal_5027 ), .Q ( signal_5028 ) ) ;
    buf_clk cell_2670 ( .C ( clk ), .D ( signal_5029 ), .Q ( signal_5030 ) ) ;
    buf_clk cell_2672 ( .C ( clk ), .D ( signal_5031 ), .Q ( signal_5032 ) ) ;
    buf_clk cell_2674 ( .C ( clk ), .D ( signal_5033 ), .Q ( signal_5034 ) ) ;
    buf_clk cell_2676 ( .C ( clk ), .D ( signal_5035 ), .Q ( signal_5036 ) ) ;
    buf_clk cell_2724 ( .C ( clk ), .D ( signal_5083 ), .Q ( signal_5084 ) ) ;
    buf_clk cell_2730 ( .C ( clk ), .D ( signal_5089 ), .Q ( signal_5090 ) ) ;
    buf_clk cell_2814 ( .C ( clk ), .D ( signal_5173 ), .Q ( signal_5174 ) ) ;
    buf_clk cell_2818 ( .C ( clk ), .D ( signal_5177 ), .Q ( signal_5178 ) ) ;
    buf_clk cell_2830 ( .C ( clk ), .D ( signal_5189 ), .Q ( signal_5190 ) ) ;
    buf_clk cell_2834 ( .C ( clk ), .D ( signal_5193 ), .Q ( signal_5194 ) ) ;
    buf_clk cell_2882 ( .C ( clk ), .D ( signal_5241 ), .Q ( signal_5242 ) ) ;
    buf_clk cell_2886 ( .C ( clk ), .D ( signal_5245 ), .Q ( signal_5246 ) ) ;
    buf_clk cell_2894 ( .C ( clk ), .D ( signal_5253 ), .Q ( signal_5254 ) ) ;
    buf_clk cell_2898 ( .C ( clk ), .D ( signal_5257 ), .Q ( signal_5258 ) ) ;
    buf_clk cell_2916 ( .C ( clk ), .D ( signal_5275 ), .Q ( signal_5276 ) ) ;
    buf_clk cell_2922 ( .C ( clk ), .D ( signal_5281 ), .Q ( signal_5282 ) ) ;
    buf_clk cell_2942 ( .C ( clk ), .D ( signal_5301 ), .Q ( signal_5302 ) ) ;
    buf_clk cell_2946 ( .C ( clk ), .D ( signal_5305 ), .Q ( signal_5306 ) ) ;
    buf_clk cell_2986 ( .C ( clk ), .D ( signal_5345 ), .Q ( signal_5346 ) ) ;
    buf_clk cell_2990 ( .C ( clk ), .D ( signal_5349 ), .Q ( signal_5350 ) ) ;
    buf_clk cell_3064 ( .C ( clk ), .D ( signal_5423 ), .Q ( signal_5424 ) ) ;
    buf_clk cell_3072 ( .C ( clk ), .D ( signal_5431 ), .Q ( signal_5432 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_2677 ( .C ( clk ), .D ( signal_1293 ), .Q ( signal_5037 ) ) ;
    buf_clk cell_2679 ( .C ( clk ), .D ( signal_2751 ), .Q ( signal_5039 ) ) ;
    buf_clk cell_2681 ( .C ( clk ), .D ( signal_4934 ), .Q ( signal_5041 ) ) ;
    buf_clk cell_2683 ( .C ( clk ), .D ( signal_4936 ), .Q ( signal_5043 ) ) ;
    buf_clk cell_2685 ( .C ( clk ), .D ( signal_1328 ), .Q ( signal_5045 ) ) ;
    buf_clk cell_2687 ( .C ( clk ), .D ( signal_2786 ), .Q ( signal_5047 ) ) ;
    buf_clk cell_2689 ( .C ( clk ), .D ( signal_1342 ), .Q ( signal_5049 ) ) ;
    buf_clk cell_2691 ( .C ( clk ), .D ( signal_2800 ), .Q ( signal_5051 ) ) ;
    buf_clk cell_2693 ( .C ( clk ), .D ( signal_1282 ), .Q ( signal_5053 ) ) ;
    buf_clk cell_2695 ( .C ( clk ), .D ( signal_2740 ), .Q ( signal_5055 ) ) ;
    buf_clk cell_2697 ( .C ( clk ), .D ( signal_1291 ), .Q ( signal_5057 ) ) ;
    buf_clk cell_2699 ( .C ( clk ), .D ( signal_2749 ), .Q ( signal_5059 ) ) ;
    buf_clk cell_2701 ( .C ( clk ), .D ( signal_4834 ), .Q ( signal_5061 ) ) ;
    buf_clk cell_2703 ( .C ( clk ), .D ( signal_4836 ), .Q ( signal_5063 ) ) ;
    buf_clk cell_2705 ( .C ( clk ), .D ( signal_4866 ), .Q ( signal_5065 ) ) ;
    buf_clk cell_2707 ( .C ( clk ), .D ( signal_4868 ), .Q ( signal_5067 ) ) ;
    buf_clk cell_2709 ( .C ( clk ), .D ( signal_4870 ), .Q ( signal_5069 ) ) ;
    buf_clk cell_2711 ( .C ( clk ), .D ( signal_4872 ), .Q ( signal_5071 ) ) ;
    buf_clk cell_2713 ( .C ( clk ), .D ( signal_4998 ), .Q ( signal_5073 ) ) ;
    buf_clk cell_2715 ( .C ( clk ), .D ( signal_5000 ), .Q ( signal_5075 ) ) ;
    buf_clk cell_2717 ( .C ( clk ), .D ( signal_4906 ), .Q ( signal_5077 ) ) ;
    buf_clk cell_2719 ( .C ( clk ), .D ( signal_4908 ), .Q ( signal_5079 ) ) ;
    buf_clk cell_2725 ( .C ( clk ), .D ( signal_5084 ), .Q ( signal_5085 ) ) ;
    buf_clk cell_2731 ( .C ( clk ), .D ( signal_5090 ), .Q ( signal_5091 ) ) ;
    buf_clk cell_2733 ( .C ( clk ), .D ( signal_4930 ), .Q ( signal_5093 ) ) ;
    buf_clk cell_2735 ( .C ( clk ), .D ( signal_4932 ), .Q ( signal_5095 ) ) ;
    buf_clk cell_2737 ( .C ( clk ), .D ( signal_5010 ), .Q ( signal_5097 ) ) ;
    buf_clk cell_2739 ( .C ( clk ), .D ( signal_5012 ), .Q ( signal_5099 ) ) ;
    buf_clk cell_2741 ( .C ( clk ), .D ( signal_4818 ), .Q ( signal_5101 ) ) ;
    buf_clk cell_2743 ( .C ( clk ), .D ( signal_4820 ), .Q ( signal_5103 ) ) ;
    buf_clk cell_2745 ( .C ( clk ), .D ( signal_4862 ), .Q ( signal_5105 ) ) ;
    buf_clk cell_2747 ( .C ( clk ), .D ( signal_4864 ), .Q ( signal_5107 ) ) ;
    buf_clk cell_2749 ( .C ( clk ), .D ( signal_1048 ), .Q ( signal_5109 ) ) ;
    buf_clk cell_2751 ( .C ( clk ), .D ( signal_2506 ), .Q ( signal_5111 ) ) ;
    buf_clk cell_2753 ( .C ( clk ), .D ( signal_4850 ), .Q ( signal_5113 ) ) ;
    buf_clk cell_2755 ( .C ( clk ), .D ( signal_4852 ), .Q ( signal_5115 ) ) ;
    buf_clk cell_2757 ( .C ( clk ), .D ( signal_1262 ), .Q ( signal_5117 ) ) ;
    buf_clk cell_2759 ( .C ( clk ), .D ( signal_2720 ), .Q ( signal_5119 ) ) ;
    buf_clk cell_2761 ( .C ( clk ), .D ( signal_1244 ), .Q ( signal_5121 ) ) ;
    buf_clk cell_2763 ( .C ( clk ), .D ( signal_2702 ), .Q ( signal_5123 ) ) ;
    buf_clk cell_2765 ( .C ( clk ), .D ( signal_1275 ), .Q ( signal_5125 ) ) ;
    buf_clk cell_2767 ( .C ( clk ), .D ( signal_2733 ), .Q ( signal_5127 ) ) ;
    buf_clk cell_2769 ( .C ( clk ), .D ( signal_1255 ), .Q ( signal_5129 ) ) ;
    buf_clk cell_2771 ( .C ( clk ), .D ( signal_2713 ), .Q ( signal_5131 ) ) ;
    buf_clk cell_2773 ( .C ( clk ), .D ( signal_1353 ), .Q ( signal_5133 ) ) ;
    buf_clk cell_2775 ( .C ( clk ), .D ( signal_2811 ), .Q ( signal_5135 ) ) ;
    buf_clk cell_2777 ( .C ( clk ), .D ( signal_1349 ), .Q ( signal_5137 ) ) ;
    buf_clk cell_2779 ( .C ( clk ), .D ( signal_2807 ), .Q ( signal_5139 ) ) ;
    buf_clk cell_2781 ( .C ( clk ), .D ( signal_1232 ), .Q ( signal_5141 ) ) ;
    buf_clk cell_2783 ( .C ( clk ), .D ( signal_2690 ), .Q ( signal_5143 ) ) ;
    buf_clk cell_2785 ( .C ( clk ), .D ( signal_1285 ), .Q ( signal_5145 ) ) ;
    buf_clk cell_2787 ( .C ( clk ), .D ( signal_2743 ), .Q ( signal_5147 ) ) ;
    buf_clk cell_2789 ( .C ( clk ), .D ( signal_1245 ), .Q ( signal_5149 ) ) ;
    buf_clk cell_2791 ( .C ( clk ), .D ( signal_2703 ), .Q ( signal_5151 ) ) ;
    buf_clk cell_2793 ( .C ( clk ), .D ( signal_1246 ), .Q ( signal_5153 ) ) ;
    buf_clk cell_2795 ( .C ( clk ), .D ( signal_2704 ), .Q ( signal_5155 ) ) ;
    buf_clk cell_2797 ( .C ( clk ), .D ( signal_1063 ), .Q ( signal_5157 ) ) ;
    buf_clk cell_2799 ( .C ( clk ), .D ( signal_2521 ), .Q ( signal_5159 ) ) ;
    buf_clk cell_2801 ( .C ( clk ), .D ( signal_1301 ), .Q ( signal_5161 ) ) ;
    buf_clk cell_2803 ( .C ( clk ), .D ( signal_2759 ), .Q ( signal_5163 ) ) ;
    buf_clk cell_2805 ( .C ( clk ), .D ( signal_1249 ), .Q ( signal_5165 ) ) ;
    buf_clk cell_2807 ( .C ( clk ), .D ( signal_2707 ), .Q ( signal_5167 ) ) ;
    buf_clk cell_2809 ( .C ( clk ), .D ( signal_1303 ), .Q ( signal_5169 ) ) ;
    buf_clk cell_2811 ( .C ( clk ), .D ( signal_2761 ), .Q ( signal_5171 ) ) ;
    buf_clk cell_2815 ( .C ( clk ), .D ( signal_5174 ), .Q ( signal_5175 ) ) ;
    buf_clk cell_2819 ( .C ( clk ), .D ( signal_5178 ), .Q ( signal_5179 ) ) ;
    buf_clk cell_2821 ( .C ( clk ), .D ( signal_1253 ), .Q ( signal_5181 ) ) ;
    buf_clk cell_2823 ( .C ( clk ), .D ( signal_2711 ), .Q ( signal_5183 ) ) ;
    buf_clk cell_2825 ( .C ( clk ), .D ( signal_1259 ), .Q ( signal_5185 ) ) ;
    buf_clk cell_2827 ( .C ( clk ), .D ( signal_2717 ), .Q ( signal_5187 ) ) ;
    buf_clk cell_2831 ( .C ( clk ), .D ( signal_5190 ), .Q ( signal_5191 ) ) ;
    buf_clk cell_2835 ( .C ( clk ), .D ( signal_5194 ), .Q ( signal_5195 ) ) ;
    buf_clk cell_2837 ( .C ( clk ), .D ( signal_1339 ), .Q ( signal_5197 ) ) ;
    buf_clk cell_2839 ( .C ( clk ), .D ( signal_2797 ), .Q ( signal_5199 ) ) ;
    buf_clk cell_2841 ( .C ( clk ), .D ( signal_4882 ), .Q ( signal_5201 ) ) ;
    buf_clk cell_2843 ( .C ( clk ), .D ( signal_4884 ), .Q ( signal_5203 ) ) ;
    buf_clk cell_2845 ( .C ( clk ), .D ( signal_1272 ), .Q ( signal_5205 ) ) ;
    buf_clk cell_2847 ( .C ( clk ), .D ( signal_2730 ), .Q ( signal_5207 ) ) ;
    buf_clk cell_2849 ( .C ( clk ), .D ( signal_1062 ), .Q ( signal_5209 ) ) ;
    buf_clk cell_2851 ( .C ( clk ), .D ( signal_2520 ), .Q ( signal_5211 ) ) ;
    buf_clk cell_2853 ( .C ( clk ), .D ( signal_1345 ), .Q ( signal_5213 ) ) ;
    buf_clk cell_2855 ( .C ( clk ), .D ( signal_2803 ), .Q ( signal_5215 ) ) ;
    buf_clk cell_2857 ( .C ( clk ), .D ( signal_1278 ), .Q ( signal_5217 ) ) ;
    buf_clk cell_2859 ( .C ( clk ), .D ( signal_2736 ), .Q ( signal_5219 ) ) ;
    buf_clk cell_2861 ( .C ( clk ), .D ( signal_1238 ), .Q ( signal_5221 ) ) ;
    buf_clk cell_2863 ( .C ( clk ), .D ( signal_2696 ), .Q ( signal_5223 ) ) ;
    buf_clk cell_2865 ( .C ( clk ), .D ( signal_1279 ), .Q ( signal_5225 ) ) ;
    buf_clk cell_2867 ( .C ( clk ), .D ( signal_2737 ), .Q ( signal_5227 ) ) ;
    buf_clk cell_2869 ( .C ( clk ), .D ( signal_1233 ), .Q ( signal_5229 ) ) ;
    buf_clk cell_2871 ( .C ( clk ), .D ( signal_2691 ), .Q ( signal_5231 ) ) ;
    buf_clk cell_2873 ( .C ( clk ), .D ( signal_1286 ), .Q ( signal_5233 ) ) ;
    buf_clk cell_2875 ( .C ( clk ), .D ( signal_2744 ), .Q ( signal_5235 ) ) ;
    buf_clk cell_2877 ( .C ( clk ), .D ( signal_1265 ), .Q ( signal_5237 ) ) ;
    buf_clk cell_2879 ( .C ( clk ), .D ( signal_2723 ), .Q ( signal_5239 ) ) ;
    buf_clk cell_2883 ( .C ( clk ), .D ( signal_5242 ), .Q ( signal_5243 ) ) ;
    buf_clk cell_2887 ( .C ( clk ), .D ( signal_5246 ), .Q ( signal_5247 ) ) ;
    buf_clk cell_2889 ( .C ( clk ), .D ( signal_4926 ), .Q ( signal_5249 ) ) ;
    buf_clk cell_2891 ( .C ( clk ), .D ( signal_4928 ), .Q ( signal_5251 ) ) ;
    buf_clk cell_2895 ( .C ( clk ), .D ( signal_5254 ), .Q ( signal_5255 ) ) ;
    buf_clk cell_2899 ( .C ( clk ), .D ( signal_5258 ), .Q ( signal_5259 ) ) ;
    buf_clk cell_2901 ( .C ( clk ), .D ( signal_1333 ), .Q ( signal_5261 ) ) ;
    buf_clk cell_2903 ( .C ( clk ), .D ( signal_2791 ), .Q ( signal_5263 ) ) ;
    buf_clk cell_2905 ( .C ( clk ), .D ( signal_4958 ), .Q ( signal_5265 ) ) ;
    buf_clk cell_2907 ( .C ( clk ), .D ( signal_4960 ), .Q ( signal_5267 ) ) ;
    buf_clk cell_2909 ( .C ( clk ), .D ( signal_4944 ), .Q ( signal_5269 ) ) ;
    buf_clk cell_2911 ( .C ( clk ), .D ( signal_4948 ), .Q ( signal_5271 ) ) ;
    buf_clk cell_2917 ( .C ( clk ), .D ( signal_5276 ), .Q ( signal_5277 ) ) ;
    buf_clk cell_2923 ( .C ( clk ), .D ( signal_5282 ), .Q ( signal_5283 ) ) ;
    buf_clk cell_2925 ( .C ( clk ), .D ( signal_4910 ), .Q ( signal_5285 ) ) ;
    buf_clk cell_2927 ( .C ( clk ), .D ( signal_4912 ), .Q ( signal_5287 ) ) ;
    buf_clk cell_2929 ( .C ( clk ), .D ( signal_4826 ), .Q ( signal_5289 ) ) ;
    buf_clk cell_2931 ( .C ( clk ), .D ( signal_4828 ), .Q ( signal_5291 ) ) ;
    buf_clk cell_2933 ( .C ( clk ), .D ( signal_4962 ), .Q ( signal_5293 ) ) ;
    buf_clk cell_2935 ( .C ( clk ), .D ( signal_4964 ), .Q ( signal_5295 ) ) ;
    buf_clk cell_2937 ( .C ( clk ), .D ( signal_1145 ), .Q ( signal_5297 ) ) ;
    buf_clk cell_2939 ( .C ( clk ), .D ( signal_2603 ), .Q ( signal_5299 ) ) ;
    buf_clk cell_2943 ( .C ( clk ), .D ( signal_5302 ), .Q ( signal_5303 ) ) ;
    buf_clk cell_2947 ( .C ( clk ), .D ( signal_5306 ), .Q ( signal_5307 ) ) ;
    buf_clk cell_2949 ( .C ( clk ), .D ( signal_1095 ), .Q ( signal_5309 ) ) ;
    buf_clk cell_2951 ( .C ( clk ), .D ( signal_2553 ), .Q ( signal_5311 ) ) ;
    buf_clk cell_2953 ( .C ( clk ), .D ( signal_1078 ), .Q ( signal_5313 ) ) ;
    buf_clk cell_2955 ( .C ( clk ), .D ( signal_2536 ), .Q ( signal_5315 ) ) ;
    buf_clk cell_2957 ( .C ( clk ), .D ( signal_1073 ), .Q ( signal_5317 ) ) ;
    buf_clk cell_2959 ( .C ( clk ), .D ( signal_2531 ), .Q ( signal_5319 ) ) ;
    buf_clk cell_2961 ( .C ( clk ), .D ( signal_1158 ), .Q ( signal_5321 ) ) ;
    buf_clk cell_2963 ( .C ( clk ), .D ( signal_2616 ), .Q ( signal_5323 ) ) ;
    buf_clk cell_2965 ( .C ( clk ), .D ( signal_1020 ), .Q ( signal_5325 ) ) ;
    buf_clk cell_2967 ( .C ( clk ), .D ( signal_2478 ), .Q ( signal_5327 ) ) ;
    buf_clk cell_2969 ( .C ( clk ), .D ( signal_5014 ), .Q ( signal_5329 ) ) ;
    buf_clk cell_2971 ( .C ( clk ), .D ( signal_5016 ), .Q ( signal_5331 ) ) ;
    buf_clk cell_2973 ( .C ( clk ), .D ( signal_4938 ), .Q ( signal_5333 ) ) ;
    buf_clk cell_2975 ( .C ( clk ), .D ( signal_4940 ), .Q ( signal_5335 ) ) ;
    buf_clk cell_2977 ( .C ( clk ), .D ( signal_1162 ), .Q ( signal_5337 ) ) ;
    buf_clk cell_2979 ( .C ( clk ), .D ( signal_2620 ), .Q ( signal_5339 ) ) ;
    buf_clk cell_2981 ( .C ( clk ), .D ( signal_1071 ), .Q ( signal_5341 ) ) ;
    buf_clk cell_2983 ( .C ( clk ), .D ( signal_2529 ), .Q ( signal_5343 ) ) ;
    buf_clk cell_2987 ( .C ( clk ), .D ( signal_5346 ), .Q ( signal_5347 ) ) ;
    buf_clk cell_2991 ( .C ( clk ), .D ( signal_5350 ), .Q ( signal_5351 ) ) ;
    buf_clk cell_2993 ( .C ( clk ), .D ( signal_1081 ), .Q ( signal_5353 ) ) ;
    buf_clk cell_2995 ( .C ( clk ), .D ( signal_2539 ), .Q ( signal_5355 ) ) ;
    buf_clk cell_2997 ( .C ( clk ), .D ( signal_4986 ), .Q ( signal_5357 ) ) ;
    buf_clk cell_2999 ( .C ( clk ), .D ( signal_4988 ), .Q ( signal_5359 ) ) ;
    buf_clk cell_3001 ( .C ( clk ), .D ( signal_4966 ), .Q ( signal_5361 ) ) ;
    buf_clk cell_3003 ( .C ( clk ), .D ( signal_4968 ), .Q ( signal_5363 ) ) ;
    buf_clk cell_3005 ( .C ( clk ), .D ( signal_1304 ), .Q ( signal_5365 ) ) ;
    buf_clk cell_3007 ( .C ( clk ), .D ( signal_2762 ), .Q ( signal_5367 ) ) ;
    buf_clk cell_3009 ( .C ( clk ), .D ( signal_1250 ), .Q ( signal_5369 ) ) ;
    buf_clk cell_3011 ( .C ( clk ), .D ( signal_2708 ), .Q ( signal_5371 ) ) ;
    buf_clk cell_3013 ( .C ( clk ), .D ( signal_1327 ), .Q ( signal_5373 ) ) ;
    buf_clk cell_3015 ( .C ( clk ), .D ( signal_2785 ), .Q ( signal_5375 ) ) ;
    buf_clk cell_3025 ( .C ( clk ), .D ( signal_5030 ), .Q ( signal_5385 ) ) ;
    buf_clk cell_3029 ( .C ( clk ), .D ( signal_5032 ), .Q ( signal_5389 ) ) ;
    buf_clk cell_3037 ( .C ( clk ), .D ( signal_1290 ), .Q ( signal_5397 ) ) ;
    buf_clk cell_3041 ( .C ( clk ), .D ( signal_2748 ), .Q ( signal_5401 ) ) ;
    buf_clk cell_3045 ( .C ( clk ), .D ( signal_1354 ), .Q ( signal_5405 ) ) ;
    buf_clk cell_3049 ( .C ( clk ), .D ( signal_2812 ), .Q ( signal_5409 ) ) ;
    buf_clk cell_3053 ( .C ( clk ), .D ( signal_1234 ), .Q ( signal_5413 ) ) ;
    buf_clk cell_3057 ( .C ( clk ), .D ( signal_2692 ), .Q ( signal_5417 ) ) ;
    buf_clk cell_3065 ( .C ( clk ), .D ( signal_5424 ), .Q ( signal_5425 ) ) ;
    buf_clk cell_3073 ( .C ( clk ), .D ( signal_5432 ), .Q ( signal_5433 ) ) ;
    buf_clk cell_3085 ( .C ( clk ), .D ( signal_1313 ), .Q ( signal_5445 ) ) ;
    buf_clk cell_3089 ( .C ( clk ), .D ( signal_2771 ), .Q ( signal_5449 ) ) ;
    buf_clk cell_3101 ( .C ( clk ), .D ( signal_1335 ), .Q ( signal_5461 ) ) ;
    buf_clk cell_3105 ( .C ( clk ), .D ( signal_2793 ), .Q ( signal_5465 ) ) ;
    buf_clk cell_3129 ( .C ( clk ), .D ( signal_1061 ), .Q ( signal_5489 ) ) ;
    buf_clk cell_3133 ( .C ( clk ), .D ( signal_2519 ), .Q ( signal_5493 ) ) ;
    buf_clk cell_3153 ( .C ( clk ), .D ( signal_1361 ), .Q ( signal_5513 ) ) ;
    buf_clk cell_3157 ( .C ( clk ), .D ( signal_2819 ), .Q ( signal_5517 ) ) ;
    buf_clk cell_3169 ( .C ( clk ), .D ( signal_4858 ), .Q ( signal_5529 ) ) ;
    buf_clk cell_3173 ( .C ( clk ), .D ( signal_4860 ), .Q ( signal_5533 ) ) ;
    buf_clk cell_3177 ( .C ( clk ), .D ( signal_4878 ), .Q ( signal_5537 ) ) ;
    buf_clk cell_3181 ( .C ( clk ), .D ( signal_4880 ), .Q ( signal_5541 ) ) ;
    buf_clk cell_3185 ( .C ( clk ), .D ( signal_4950 ), .Q ( signal_5545 ) ) ;
    buf_clk cell_3189 ( .C ( clk ), .D ( signal_4952 ), .Q ( signal_5549 ) ) ;
    buf_clk cell_3193 ( .C ( clk ), .D ( signal_4830 ), .Q ( signal_5553 ) ) ;
    buf_clk cell_3197 ( .C ( clk ), .D ( signal_4832 ), .Q ( signal_5557 ) ) ;
    buf_clk cell_3221 ( .C ( clk ), .D ( signal_4842 ), .Q ( signal_5581 ) ) ;
    buf_clk cell_3225 ( .C ( clk ), .D ( signal_4844 ), .Q ( signal_5585 ) ) ;
    buf_clk cell_3229 ( .C ( clk ), .D ( signal_4838 ), .Q ( signal_5589 ) ) ;
    buf_clk cell_3233 ( .C ( clk ), .D ( signal_4840 ), .Q ( signal_5593 ) ) ;
    buf_clk cell_3237 ( .C ( clk ), .D ( signal_4914 ), .Q ( signal_5597 ) ) ;
    buf_clk cell_3241 ( .C ( clk ), .D ( signal_4916 ), .Q ( signal_5601 ) ) ;
    buf_clk cell_3249 ( .C ( clk ), .D ( signal_4874 ), .Q ( signal_5609 ) ) ;
    buf_clk cell_3253 ( .C ( clk ), .D ( signal_4876 ), .Q ( signal_5613 ) ) ;
    buf_clk cell_3277 ( .C ( clk ), .D ( signal_1080 ), .Q ( signal_5637 ) ) ;
    buf_clk cell_3281 ( .C ( clk ), .D ( signal_2538 ), .Q ( signal_5641 ) ) ;
    buf_clk cell_3285 ( .C ( clk ), .D ( signal_1365 ), .Q ( signal_5645 ) ) ;
    buf_clk cell_3289 ( .C ( clk ), .D ( signal_2823 ), .Q ( signal_5649 ) ) ;
    buf_clk cell_3297 ( .C ( clk ), .D ( signal_1242 ), .Q ( signal_5657 ) ) ;
    buf_clk cell_3301 ( .C ( clk ), .D ( signal_2700 ), .Q ( signal_5661 ) ) ;
    buf_clk cell_3313 ( .C ( clk ), .D ( signal_1296 ), .Q ( signal_5673 ) ) ;
    buf_clk cell_3317 ( .C ( clk ), .D ( signal_2754 ), .Q ( signal_5677 ) ) ;
    buf_clk cell_3321 ( .C ( clk ), .D ( signal_1308 ), .Q ( signal_5681 ) ) ;
    buf_clk cell_3325 ( .C ( clk ), .D ( signal_2766 ), .Q ( signal_5685 ) ) ;
    buf_clk cell_3329 ( .C ( clk ), .D ( signal_1251 ), .Q ( signal_5689 ) ) ;
    buf_clk cell_3333 ( .C ( clk ), .D ( signal_2709 ), .Q ( signal_5693 ) ) ;
    buf_clk cell_3341 ( .C ( clk ), .D ( signal_1326 ), .Q ( signal_5701 ) ) ;
    buf_clk cell_3345 ( .C ( clk ), .D ( signal_2784 ), .Q ( signal_5705 ) ) ;
    buf_clk cell_3349 ( .C ( clk ), .D ( signal_1261 ), .Q ( signal_5709 ) ) ;
    buf_clk cell_3353 ( .C ( clk ), .D ( signal_2719 ), .Q ( signal_5713 ) ) ;
    buf_clk cell_3361 ( .C ( clk ), .D ( signal_1271 ), .Q ( signal_5721 ) ) ;
    buf_clk cell_3365 ( .C ( clk ), .D ( signal_2729 ), .Q ( signal_5725 ) ) ;
    buf_clk cell_3381 ( .C ( clk ), .D ( signal_4822 ), .Q ( signal_5741 ) ) ;
    buf_clk cell_3385 ( .C ( clk ), .D ( signal_4824 ), .Q ( signal_5745 ) ) ;
    buf_clk cell_3393 ( .C ( clk ), .D ( signal_5034 ), .Q ( signal_5753 ) ) ;
    buf_clk cell_3399 ( .C ( clk ), .D ( signal_5036 ), .Q ( signal_5759 ) ) ;
    buf_clk cell_3405 ( .C ( clk ), .D ( signal_1248 ), .Q ( signal_5765 ) ) ;
    buf_clk cell_3411 ( .C ( clk ), .D ( signal_2706 ), .Q ( signal_5771 ) ) ;
    buf_clk cell_3417 ( .C ( clk ), .D ( signal_1314 ), .Q ( signal_5777 ) ) ;
    buf_clk cell_3423 ( .C ( clk ), .D ( signal_2772 ), .Q ( signal_5783 ) ) ;
    buf_clk cell_3437 ( .C ( clk ), .D ( signal_1336 ), .Q ( signal_5797 ) ) ;
    buf_clk cell_3443 ( .C ( clk ), .D ( signal_2794 ), .Q ( signal_5803 ) ) ;
    buf_clk cell_3489 ( .C ( clk ), .D ( signal_4918 ), .Q ( signal_5849 ) ) ;
    buf_clk cell_3495 ( .C ( clk ), .D ( signal_4920 ), .Q ( signal_5855 ) ) ;
    buf_clk cell_3549 ( .C ( clk ), .D ( signal_4810 ), .Q ( signal_5909 ) ) ;
    buf_clk cell_3555 ( .C ( clk ), .D ( signal_4812 ), .Q ( signal_5915 ) ) ;
    buf_clk cell_3581 ( .C ( clk ), .D ( signal_1298 ), .Q ( signal_5941 ) ) ;
    buf_clk cell_3587 ( .C ( clk ), .D ( signal_2756 ), .Q ( signal_5947 ) ) ;
    buf_clk cell_3637 ( .C ( clk ), .D ( signal_1064 ), .Q ( signal_5997 ) ) ;
    buf_clk cell_3643 ( .C ( clk ), .D ( signal_2522 ), .Q ( signal_6003 ) ) ;
    buf_clk cell_3657 ( .C ( clk ), .D ( signal_1316 ), .Q ( signal_6017 ) ) ;
    buf_clk cell_3663 ( .C ( clk ), .D ( signal_2774 ), .Q ( signal_6023 ) ) ;
    buf_clk cell_3713 ( .C ( clk ), .D ( signal_1289 ), .Q ( signal_6073 ) ) ;
    buf_clk cell_3719 ( .C ( clk ), .D ( signal_2747 ), .Q ( signal_6079 ) ) ;
    buf_clk cell_3741 ( .C ( clk ), .D ( signal_1359 ), .Q ( signal_6101 ) ) ;
    buf_clk cell_3747 ( .C ( clk ), .D ( signal_2817 ), .Q ( signal_6107 ) ) ;
    buf_clk cell_3753 ( .C ( clk ), .D ( signal_1307 ), .Q ( signal_6113 ) ) ;
    buf_clk cell_3759 ( .C ( clk ), .D ( signal_2765 ), .Q ( signal_6119 ) ) ;
    buf_clk cell_3765 ( .C ( clk ), .D ( signal_4954 ), .Q ( signal_6125 ) ) ;
    buf_clk cell_3771 ( .C ( clk ), .D ( signal_4956 ), .Q ( signal_6131 ) ) ;
    buf_clk cell_3793 ( .C ( clk ), .D ( signal_1315 ), .Q ( signal_6153 ) ) ;
    buf_clk cell_3801 ( .C ( clk ), .D ( signal_2773 ), .Q ( signal_6161 ) ) ;
    buf_clk cell_3965 ( .C ( clk ), .D ( signal_1239 ), .Q ( signal_6325 ) ) ;
    buf_clk cell_3973 ( .C ( clk ), .D ( signal_2697 ), .Q ( signal_6333 ) ) ;
    buf_clk cell_4029 ( .C ( clk ), .D ( signal_1060 ), .Q ( signal_6389 ) ) ;
    buf_clk cell_4037 ( .C ( clk ), .D ( signal_2518 ), .Q ( signal_6397 ) ) ;
    buf_clk cell_4129 ( .C ( clk ), .D ( signal_1254 ), .Q ( signal_6489 ) ) ;
    buf_clk cell_4139 ( .C ( clk ), .D ( signal_2712 ), .Q ( signal_6499 ) ) ;
    buf_clk cell_4225 ( .C ( clk ), .D ( signal_1247 ), .Q ( signal_6585 ) ) ;
    buf_clk cell_4235 ( .C ( clk ), .D ( signal_2705 ), .Q ( signal_6595 ) ) ;
    buf_clk cell_4337 ( .C ( clk ), .D ( signal_1066 ), .Q ( signal_6697 ) ) ;
    buf_clk cell_4347 ( .C ( clk ), .D ( signal_2524 ), .Q ( signal_6707 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1085 ( .a ({signal_4804, signal_4800}), .b ({signal_2472, signal_1014}), .clk ( clk ), .r ( Fresh[238] ), .c ({signal_2558, signal_1100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1124 ( .a ({signal_4808, signal_4806}), .b ({signal_2477, signal_1019}), .clk ( clk ), .r ( Fresh[239] ), .c ({signal_2597, signal_1139}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1132 ( .a ({signal_4812, signal_4810}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[240] ), .c ({signal_2605, signal_1147}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1140 ( .a ({signal_4816, signal_4814}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[241] ), .c ({signal_2613, signal_1155}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1155 ( .a ({signal_4820, signal_4818}), .b ({signal_2478, signal_1020}), .clk ( clk ), .r ( Fresh[242] ), .c ({signal_2628, signal_1170}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1173 ( .a ({signal_4824, signal_4822}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[243] ), .c ({signal_2646, signal_1188}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1184 ( .a ({signal_4828, signal_4826}), .b ({signal_2482, signal_1024}), .clk ( clk ), .r ( Fresh[244] ), .c ({signal_2657, signal_1199}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1189 ( .a ({signal_4832, signal_4830}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[245] ), .c ({signal_2662, signal_1204}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1190 ( .a ({signal_4836, signal_4834}), .b ({signal_2482, signal_1024}), .clk ( clk ), .r ( Fresh[246] ), .c ({signal_2663, signal_1205}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1198 ( .a ({signal_4840, signal_4838}), .b ({signal_2482, signal_1024}), .clk ( clk ), .r ( Fresh[247] ), .c ({signal_2671, signal_1213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1207 ( .a ({signal_4844, signal_4842}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[248] ), .c ({signal_2680, signal_1222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1209 ( .a ({signal_4848, signal_4846}), .b ({signal_2484, signal_1026}), .clk ( clk ), .r ( Fresh[249] ), .c ({signal_2682, signal_1224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1211 ( .a ({signal_4852, signal_4850}), .b ({signal_2478, signal_1020}), .clk ( clk ), .r ( Fresh[250] ), .c ({signal_2684, signal_1226}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1212 ( .a ({signal_4856, signal_4854}), .b ({signal_2478, signal_1020}), .clk ( clk ), .r ( Fresh[251] ), .c ({signal_2685, signal_1227}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1243 ( .a ({signal_2558, signal_1100}), .b ({signal_2716, signal_1258}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1272 ( .a ({signal_2597, signal_1139}), .b ({signal_2745, signal_1287}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1277 ( .a ({signal_2605, signal_1147}), .b ({signal_2750, signal_1292}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1284 ( .a ({signal_2613, signal_1155}), .b ({signal_2757, signal_1299}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1297 ( .a ({signal_2628, signal_1170}), .b ({signal_2770, signal_1312}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1314 ( .a ({signal_2646, signal_1188}), .b ({signal_2787, signal_1329}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1323 ( .a ({signal_2657, signal_1199}), .b ({signal_2796, signal_1338}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1328 ( .a ({signal_2662, signal_1204}), .b ({signal_2801, signal_1343}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1329 ( .a ({signal_2663, signal_1205}), .b ({signal_2802, signal_1344}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1335 ( .a ({signal_2671, signal_1213}), .b ({signal_2808, signal_1350}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1343 ( .a ({signal_2680, signal_1222}), .b ({signal_2816, signal_1358}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1345 ( .a ({signal_2682, signal_1224}), .b ({signal_2818, signal_1360}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1347 ( .a ({signal_2684, signal_1226}), .b ({signal_2820, signal_1362}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1348 ( .a ({signal_2685, signal_1227}), .b ({signal_2821, signal_1363}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1351 ( .a ({signal_4860, signal_4858}), .b ({signal_2525, signal_1067}), .clk ( clk ), .r ( Fresh[252] ), .c ({signal_2824, signal_1366}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1352 ( .a ({signal_4864, signal_4862}), .b ({signal_2526, signal_1068}), .clk ( clk ), .r ( Fresh[253] ), .c ({signal_2825, signal_1367}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1358 ( .a ({signal_4824, signal_4822}), .b ({signal_2538, signal_1080}), .clk ( clk ), .r ( Fresh[254] ), .c ({signal_2831, signal_1373}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1359 ( .a ({signal_4844, signal_4842}), .b ({signal_2543, signal_1085}), .clk ( clk ), .r ( Fresh[255] ), .c ({signal_2832, signal_1374}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1363 ( .a ({signal_4836, signal_4834}), .b ({signal_2547, signal_1089}), .clk ( clk ), .r ( Fresh[256] ), .c ({signal_2836, signal_1378}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1364 ( .a ({signal_4868, signal_4866}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[257] ), .c ({signal_2837, signal_1379}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1370 ( .a ({signal_4872, signal_4870}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[258] ), .c ({signal_2843, signal_1385}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1371 ( .a ({signal_4876, signal_4874}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[259] ), .c ({signal_2844, signal_1386}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1372 ( .a ({signal_4880, signal_4878}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[260] ), .c ({signal_2845, signal_1387}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1373 ( .a ({signal_2531, signal_1073}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[261] ), .c ({signal_2846, signal_1388}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1374 ( .a ({signal_4884, signal_4882}), .b ({signal_2555, signal_1097}), .clk ( clk ), .r ( Fresh[262] ), .c ({signal_2847, signal_1389}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1377 ( .a ({signal_4888, signal_4886}), .b ({signal_2562, signal_1104}), .clk ( clk ), .r ( Fresh[263] ), .c ({signal_2850, signal_1392}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1378 ( .a ({signal_4892, signal_4890}), .b ({signal_2536, signal_1078}), .clk ( clk ), .r ( Fresh[264] ), .c ({signal_2851, signal_1393}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1379 ( .a ({signal_4852, signal_4850}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[265] ), .c ({signal_2852, signal_1394}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1380 ( .a ({signal_4884, signal_4882}), .b ({signal_2547, signal_1089}), .clk ( clk ), .r ( Fresh[266] ), .c ({signal_2853, signal_1395}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1381 ( .a ({signal_4836, signal_4834}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[267] ), .c ({signal_2854, signal_1396}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1382 ( .a ({signal_4896, signal_4894}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[268] ), .c ({signal_2855, signal_1397}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1384 ( .a ({signal_4900, signal_4898}), .b ({signal_2565, signal_1107}), .clk ( clk ), .r ( Fresh[269] ), .c ({signal_2857, signal_1399}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1385 ( .a ({signal_4828, signal_4826}), .b ({signal_2550, signal_1092}), .clk ( clk ), .r ( Fresh[270] ), .c ({signal_2858, signal_1400}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1386 ( .a ({signal_4904, signal_4902}), .b ({signal_2538, signal_1080}), .clk ( clk ), .r ( Fresh[271] ), .c ({signal_2859, signal_1401}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1387 ( .a ({signal_4908, signal_4906}), .b ({signal_2544, signal_1086}), .clk ( clk ), .r ( Fresh[272] ), .c ({signal_2860, signal_1402}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1388 ( .a ({signal_4912, signal_4910}), .b ({signal_2572, signal_1114}), .clk ( clk ), .r ( Fresh[273] ), .c ({signal_2861, signal_1403}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1389 ( .a ({signal_4916, signal_4914}), .b ({signal_2566, signal_1108}), .clk ( clk ), .r ( Fresh[274] ), .c ({signal_2862, signal_1404}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1390 ( .a ({signal_4872, signal_4870}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[275] ), .c ({signal_2863, signal_1405}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1391 ( .a ({signal_4820, signal_4818}), .b ({signal_2555, signal_1097}), .clk ( clk ), .r ( Fresh[276] ), .c ({signal_2864, signal_1406}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1392 ( .a ({signal_4912, signal_4910}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[277] ), .c ({signal_2865, signal_1407}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1393 ( .a ({signal_4920, signal_4918}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[278] ), .c ({signal_2866, signal_1408}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1394 ( .a ({signal_4872, signal_4870}), .b ({signal_2572, signal_1114}), .clk ( clk ), .r ( Fresh[279] ), .c ({signal_2867, signal_1409}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1397 ( .a ({signal_4852, signal_4850}), .b ({signal_2560, signal_1102}), .clk ( clk ), .r ( Fresh[280] ), .c ({signal_2870, signal_1412}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1398 ( .a ({signal_4856, signal_4854}), .b ({signal_2581, signal_1123}), .clk ( clk ), .r ( Fresh[281] ), .c ({signal_2871, signal_1413}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1399 ( .a ({signal_4924, signal_4922}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[282] ), .c ({signal_2872, signal_1414}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1400 ( .a ({signal_4872, signal_4870}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[283] ), .c ({signal_2873, signal_1415}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1404 ( .a ({signal_4880, signal_4878}), .b ({signal_2536, signal_1078}), .clk ( clk ), .r ( Fresh[284] ), .c ({signal_2877, signal_1419}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1405 ( .a ({signal_4836, signal_4834}), .b ({signal_2560, signal_1102}), .clk ( clk ), .r ( Fresh[285] ), .c ({signal_2878, signal_1420}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1406 ( .a ({signal_4928, signal_4926}), .b ({signal_2573, signal_1115}), .clk ( clk ), .r ( Fresh[286] ), .c ({signal_2879, signal_1421}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1409 ( .a ({signal_4932, signal_4930}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[287] ), .c ({signal_2882, signal_1424}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1410 ( .a ({signal_4808, signal_4806}), .b ({signal_2565, signal_1107}), .clk ( clk ), .r ( Fresh[288] ), .c ({signal_2883, signal_1425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1411 ( .a ({signal_4880, signal_4878}), .b ({signal_2544, signal_1086}), .clk ( clk ), .r ( Fresh[289] ), .c ({signal_2884, signal_1426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1412 ( .a ({signal_4820, signal_4818}), .b ({signal_2586, signal_1128}), .clk ( clk ), .r ( Fresh[290] ), .c ({signal_2885, signal_1427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1413 ( .a ({signal_4936, signal_4934}), .b ({signal_2530, signal_1072}), .clk ( clk ), .r ( Fresh[291] ), .c ({signal_2886, signal_1428}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1414 ( .a ({signal_4940, signal_4938}), .b ({signal_2591, signal_1133}), .clk ( clk ), .r ( Fresh[292] ), .c ({signal_2887, signal_1429}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1415 ( .a ({signal_4876, signal_4874}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[293] ), .c ({signal_2888, signal_1430}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1416 ( .a ({signal_4948, signal_4944}), .b ({signal_2596, signal_1138}), .clk ( clk ), .r ( Fresh[294] ), .c ({signal_2889, signal_1431}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1417 ( .a ({signal_4856, signal_4854}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[295] ), .c ({signal_2890, signal_1432}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1418 ( .a ({signal_4952, signal_4950}), .b ({signal_2598, signal_1140}), .clk ( clk ), .r ( Fresh[296] ), .c ({signal_2891, signal_1433}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1419 ( .a ({signal_4956, signal_4954}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[297] ), .c ({signal_2892, signal_1434}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1420 ( .a ({signal_4864, signal_4862}), .b ({signal_2600, signal_1142}), .clk ( clk ), .r ( Fresh[298] ), .c ({signal_2893, signal_1435}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1421 ( .a ({signal_4924, signal_4922}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[299] ), .c ({signal_2894, signal_1436}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1422 ( .a ({signal_4864, signal_4862}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[300] ), .c ({signal_2895, signal_1437}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1423 ( .a ({signal_4884, signal_4882}), .b ({signal_2609, signal_1151}), .clk ( clk ), .r ( Fresh[301] ), .c ({signal_2896, signal_1438}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1424 ( .a ({signal_4960, signal_4958}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[302] ), .c ({signal_2897, signal_1439}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1425 ( .a ({signal_4872, signal_4870}), .b ({signal_2614, signal_1156}), .clk ( clk ), .r ( Fresh[303] ), .c ({signal_2898, signal_1440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1426 ( .a ({signal_4888, signal_4886}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[304] ), .c ({signal_2899, signal_1441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1427 ( .a ({signal_4864, signal_4862}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[305] ), .c ({signal_2900, signal_1442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1428 ( .a ({signal_4928, signal_4926}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[306] ), .c ({signal_2901, signal_1443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1429 ( .a ({signal_4860, signal_4858}), .b ({signal_2624, signal_1166}), .clk ( clk ), .r ( Fresh[307] ), .c ({signal_2902, signal_1444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1430 ( .a ({signal_2544, signal_1086}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[308] ), .c ({signal_2903, signal_1445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1431 ( .a ({signal_4964, signal_4962}), .b ({signal_2626, signal_1168}), .clk ( clk ), .r ( Fresh[309] ), .c ({signal_2904, signal_1446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1432 ( .a ({signal_2480, signal_1022}), .b ({signal_2600, signal_1142}), .clk ( clk ), .r ( Fresh[310] ), .c ({signal_2905, signal_1447}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1433 ( .a ({signal_4828, signal_4826}), .b ({signal_2594, signal_1136}), .clk ( clk ), .r ( Fresh[311] ), .c ({signal_2906, signal_1448}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1434 ( .a ({signal_2601, signal_1143}), .b ({signal_2603, signal_1145}), .clk ( clk ), .r ( Fresh[312] ), .c ({signal_2907, signal_1449}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1435 ( .a ({signal_4900, signal_4898}), .b ({signal_2624, signal_1166}), .clk ( clk ), .r ( Fresh[313] ), .c ({signal_2908, signal_1450}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1436 ( .a ({signal_4968, signal_4966}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[314] ), .c ({signal_2909, signal_1451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1437 ( .a ({signal_4912, signal_4910}), .b ({signal_2634, signal_1176}), .clk ( clk ), .r ( Fresh[315] ), .c ({signal_2910, signal_1452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1438 ( .a ({signal_2594, signal_1136}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[316] ), .c ({signal_2911, signal_1453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1439 ( .a ({signal_2549, signal_1091}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[317] ), .c ({signal_2912, signal_1454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1440 ( .a ({signal_4848, signal_4846}), .b ({signal_2615, signal_1157}), .clk ( clk ), .r ( Fresh[318] ), .c ({signal_2913, signal_1455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1441 ( .a ({signal_4820, signal_4818}), .b ({signal_2636, signal_1178}), .clk ( clk ), .r ( Fresh[319] ), .c ({signal_2914, signal_1456}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1442 ( .a ({signal_4932, signal_4930}), .b ({signal_2540, signal_1082}), .clk ( clk ), .r ( Fresh[320] ), .c ({signal_2915, signal_1457}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1443 ( .a ({signal_4940, signal_4938}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[321] ), .c ({signal_2916, signal_1458}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1444 ( .a ({signal_4884, signal_4882}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[322] ), .c ({signal_2917, signal_1459}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1445 ( .a ({signal_4876, signal_4874}), .b ({signal_2647, signal_1189}), .clk ( clk ), .r ( Fresh[323] ), .c ({signal_2918, signal_1460}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1446 ( .a ({signal_4972, signal_4970}), .b ({signal_2648, signal_1190}), .clk ( clk ), .r ( Fresh[324] ), .c ({signal_2919, signal_1461}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1447 ( .a ({signal_4876, signal_4874}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[325] ), .c ({signal_2920, signal_1462}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1448 ( .a ({signal_4976, signal_4974}), .b ({signal_2615, signal_1157}), .clk ( clk ), .r ( Fresh[326] ), .c ({signal_2921, signal_1463}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1449 ( .a ({signal_4912, signal_4910}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[327] ), .c ({signal_2922, signal_1464}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1450 ( .a ({signal_4960, signal_4958}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[328] ), .c ({signal_2923, signal_1465}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1451 ( .a ({signal_4980, signal_4978}), .b ({signal_2656, signal_1198}), .clk ( clk ), .r ( Fresh[329] ), .c ({signal_2924, signal_1466}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1452 ( .a ({signal_4984, signal_4982}), .b ({signal_2603, signal_1145}), .clk ( clk ), .r ( Fresh[330] ), .c ({signal_2925, signal_1467}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1453 ( .a ({signal_4988, signal_4986}), .b ({signal_2650, signal_1192}), .clk ( clk ), .r ( Fresh[331] ), .c ({signal_2926, signal_1468}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1454 ( .a ({signal_2560, signal_1102}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[332] ), .c ({signal_2927, signal_1469}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1455 ( .a ({signal_4820, signal_4818}), .b ({signal_2635, signal_1177}), .clk ( clk ), .r ( Fresh[333] ), .c ({signal_2928, signal_1470}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1456 ( .a ({signal_4872, signal_4870}), .b ({signal_2540, signal_1082}), .clk ( clk ), .r ( Fresh[334] ), .c ({signal_2929, signal_1471}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1457 ( .a ({signal_4928, signal_4926}), .b ({signal_2649, signal_1191}), .clk ( clk ), .r ( Fresh[335] ), .c ({signal_2930, signal_1472}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1458 ( .a ({signal_4896, signal_4894}), .b ({signal_2602, signal_1144}), .clk ( clk ), .r ( Fresh[336] ), .c ({signal_2931, signal_1473}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1459 ( .a ({signal_4876, signal_4874}), .b ({signal_2635, signal_1177}), .clk ( clk ), .r ( Fresh[337] ), .c ({signal_2932, signal_1474}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1460 ( .a ({signal_4916, signal_4914}), .b ({signal_2644, signal_1186}), .clk ( clk ), .r ( Fresh[338] ), .c ({signal_2933, signal_1475}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1461 ( .a ({signal_4880, signal_4878}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[339] ), .c ({signal_2934, signal_1476}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1462 ( .a ({signal_4852, signal_4850}), .b ({signal_2540, signal_1082}), .clk ( clk ), .r ( Fresh[340] ), .c ({signal_2935, signal_1477}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1463 ( .a ({signal_4884, signal_4882}), .b ({signal_2664, signal_1206}), .clk ( clk ), .r ( Fresh[341] ), .c ({signal_2936, signal_1478}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1464 ( .a ({signal_4940, signal_4938}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[342] ), .c ({signal_2937, signal_1479}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1465 ( .a ({signal_4824, signal_4822}), .b ({signal_2644, signal_1186}), .clk ( clk ), .r ( Fresh[343] ), .c ({signal_2938, signal_1480}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1466 ( .a ({signal_2533, signal_1075}), .b ({signal_2539, signal_1081}), .clk ( clk ), .r ( Fresh[344] ), .c ({signal_2939, signal_1481}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1467 ( .a ({signal_4840, signal_4838}), .b ({signal_2626, signal_1168}), .clk ( clk ), .r ( Fresh[345] ), .c ({signal_2940, signal_1482}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1468 ( .a ({signal_4928, signal_4926}), .b ({signal_2619, signal_1161}), .clk ( clk ), .r ( Fresh[346] ), .c ({signal_2941, signal_1483}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1469 ( .a ({signal_2479, signal_1021}), .b ({signal_2590, signal_1132}), .clk ( clk ), .r ( Fresh[347] ), .c ({signal_2942, signal_1484}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1470 ( .a ({signal_4908, signal_4906}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[348] ), .c ({signal_2943, signal_1485}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1471 ( .a ({signal_4992, signal_4990}), .b ({signal_2666, signal_1208}), .clk ( clk ), .r ( Fresh[349] ), .c ({signal_2944, signal_1486}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1472 ( .a ({signal_4852, signal_4850}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[350] ), .c ({signal_2945, signal_1487}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1473 ( .a ({signal_4896, signal_4894}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[351] ), .c ({signal_2946, signal_1488}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1474 ( .a ({signal_4996, signal_4994}), .b ({signal_2659, signal_1201}), .clk ( clk ), .r ( Fresh[352] ), .c ({signal_2947, signal_1489}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1475 ( .a ({signal_4836, signal_4834}), .b ({signal_2619, signal_1161}), .clk ( clk ), .r ( Fresh[353] ), .c ({signal_2948, signal_1490}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1476 ( .a ({signal_4804, signal_4800}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[354] ), .c ({signal_2949, signal_1491}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1477 ( .a ({signal_4940, signal_4938}), .b ({signal_2675, signal_1217}), .clk ( clk ), .r ( Fresh[355] ), .c ({signal_2950, signal_1492}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1478 ( .a ({signal_4936, signal_4934}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[356] ), .c ({signal_2951, signal_1493}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1479 ( .a ({signal_4804, signal_4800}), .b ({signal_2647, signal_1189}), .clk ( clk ), .r ( Fresh[357] ), .c ({signal_2952, signal_1494}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1480 ( .a ({signal_5000, signal_4998}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[358] ), .c ({signal_2953, signal_1495}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1481 ( .a ({signal_4852, signal_4850}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[359] ), .c ({signal_2954, signal_1496}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1482 ( .a ({signal_4884, signal_4882}), .b ({signal_2602, signal_1144}), .clk ( clk ), .r ( Fresh[360] ), .c ({signal_2955, signal_1497}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1483 ( .a ({signal_4880, signal_4878}), .b ({signal_2602, signal_1144}), .clk ( clk ), .r ( Fresh[361] ), .c ({signal_2956, signal_1498}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1484 ( .a ({signal_4856, signal_4854}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[362] ), .c ({signal_2957, signal_1499}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1485 ( .a ({signal_4804, signal_4800}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[363] ), .c ({signal_2958, signal_1500}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1486 ( .a ({signal_4932, signal_4930}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[364] ), .c ({signal_2959, signal_1501}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1487 ( .a ({signal_4872, signal_4870}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[365] ), .c ({signal_2960, signal_1502}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1488 ( .a ({signal_4884, signal_4882}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[366] ), .c ({signal_2961, signal_1503}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1489 ( .a ({signal_4860, signal_4858}), .b ({signal_2577, signal_1119}), .clk ( clk ), .r ( Fresh[367] ), .c ({signal_2962, signal_1504}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1490 ( .a ({signal_2824, signal_1366}), .b ({signal_2963, signal_1505}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1491 ( .a ({signal_2825, signal_1367}), .b ({signal_2964, signal_1506}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1497 ( .a ({signal_2831, signal_1373}), .b ({signal_2970, signal_1512}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1498 ( .a ({signal_2832, signal_1374}), .b ({signal_2971, signal_1513}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1502 ( .a ({signal_2836, signal_1378}), .b ({signal_2975, signal_1517}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1503 ( .a ({signal_2837, signal_1379}), .b ({signal_2976, signal_1518}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1508 ( .a ({signal_2843, signal_1385}), .b ({signal_2981, signal_1523}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1509 ( .a ({signal_2844, signal_1386}), .b ({signal_2982, signal_1524}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1510 ( .a ({signal_2845, signal_1387}), .b ({signal_2983, signal_1525}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1511 ( .a ({signal_2846, signal_1388}), .b ({signal_2984, signal_1526}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1512 ( .a ({signal_2847, signal_1389}), .b ({signal_2985, signal_1527}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1514 ( .a ({signal_2850, signal_1392}), .b ({signal_2987, signal_1529}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1515 ( .a ({signal_2851, signal_1393}), .b ({signal_2988, signal_1530}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1516 ( .a ({signal_2852, signal_1394}), .b ({signal_2989, signal_1531}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1517 ( .a ({signal_2853, signal_1395}), .b ({signal_2990, signal_1532}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1518 ( .a ({signal_2854, signal_1396}), .b ({signal_2991, signal_1533}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1519 ( .a ({signal_2855, signal_1397}), .b ({signal_2992, signal_1534}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1521 ( .a ({signal_2857, signal_1399}), .b ({signal_2994, signal_1536}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1522 ( .a ({signal_2858, signal_1400}), .b ({signal_2995, signal_1537}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1523 ( .a ({signal_2859, signal_1401}), .b ({signal_2996, signal_1538}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1524 ( .a ({signal_2860, signal_1402}), .b ({signal_2997, signal_1539}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1525 ( .a ({signal_2861, signal_1403}), .b ({signal_2998, signal_1540}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1526 ( .a ({signal_2862, signal_1404}), .b ({signal_2999, signal_1541}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1527 ( .a ({signal_2863, signal_1405}), .b ({signal_3000, signal_1542}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1528 ( .a ({signal_2864, signal_1406}), .b ({signal_3001, signal_1543}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1529 ( .a ({signal_2865, signal_1407}), .b ({signal_3002, signal_1544}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1530 ( .a ({signal_2866, signal_1408}), .b ({signal_3003, signal_1545}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1531 ( .a ({signal_2867, signal_1409}), .b ({signal_3004, signal_1546}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1534 ( .a ({signal_2870, signal_1412}), .b ({signal_3007, signal_1549}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1535 ( .a ({signal_2871, signal_1413}), .b ({signal_3008, signal_1550}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1536 ( .a ({signal_2872, signal_1414}), .b ({signal_3009, signal_1551}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1537 ( .a ({signal_2873, signal_1415}), .b ({signal_3010, signal_1552}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1540 ( .a ({signal_2877, signal_1419}), .b ({signal_3013, signal_1555}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1541 ( .a ({signal_2878, signal_1420}), .b ({signal_3014, signal_1556}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1542 ( .a ({signal_2879, signal_1421}), .b ({signal_3015, signal_1557}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1545 ( .a ({signal_2882, signal_1424}), .b ({signal_3018, signal_1560}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1546 ( .a ({signal_2883, signal_1425}), .b ({signal_3019, signal_1561}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1547 ( .a ({signal_2884, signal_1426}), .b ({signal_3020, signal_1562}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1548 ( .a ({signal_2885, signal_1427}), .b ({signal_3021, signal_1563}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1549 ( .a ({signal_2886, signal_1428}), .b ({signal_3022, signal_1564}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1550 ( .a ({signal_2887, signal_1429}), .b ({signal_3023, signal_1565}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1551 ( .a ({signal_2888, signal_1430}), .b ({signal_3024, signal_1566}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1552 ( .a ({signal_2889, signal_1431}), .b ({signal_3025, signal_1567}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1553 ( .a ({signal_2890, signal_1432}), .b ({signal_3026, signal_1568}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1554 ( .a ({signal_2891, signal_1433}), .b ({signal_3027, signal_1569}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1555 ( .a ({signal_2892, signal_1434}), .b ({signal_3028, signal_1570}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1556 ( .a ({signal_2893, signal_1435}), .b ({signal_3029, signal_1571}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1557 ( .a ({signal_2894, signal_1436}), .b ({signal_3030, signal_1572}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1558 ( .a ({signal_2895, signal_1437}), .b ({signal_3031, signal_1573}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1559 ( .a ({signal_2896, signal_1438}), .b ({signal_3032, signal_1574}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1560 ( .a ({signal_2897, signal_1439}), .b ({signal_3033, signal_1575}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1561 ( .a ({signal_2898, signal_1440}), .b ({signal_3034, signal_1576}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1562 ( .a ({signal_2899, signal_1441}), .b ({signal_3035, signal_1577}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1563 ( .a ({signal_2900, signal_1442}), .b ({signal_3036, signal_1578}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1564 ( .a ({signal_2901, signal_1443}), .b ({signal_3037, signal_1579}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1565 ( .a ({signal_2902, signal_1444}), .b ({signal_3038, signal_1580}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1566 ( .a ({signal_2903, signal_1445}), .b ({signal_3039, signal_1581}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1567 ( .a ({signal_2905, signal_1447}), .b ({signal_3040, signal_1582}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1568 ( .a ({signal_2906, signal_1448}), .b ({signal_3041, signal_1583}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1569 ( .a ({signal_2907, signal_1449}), .b ({signal_3042, signal_1584}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1570 ( .a ({signal_2908, signal_1450}), .b ({signal_3043, signal_1585}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1571 ( .a ({signal_2909, signal_1451}), .b ({signal_3044, signal_1586}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1572 ( .a ({signal_2910, signal_1452}), .b ({signal_3045, signal_1587}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1573 ( .a ({signal_2911, signal_1453}), .b ({signal_3046, signal_1588}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1574 ( .a ({signal_2912, signal_1454}), .b ({signal_3047, signal_1589}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1575 ( .a ({signal_2913, signal_1455}), .b ({signal_3048, signal_1590}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1576 ( .a ({signal_2914, signal_1456}), .b ({signal_3049, signal_1591}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1577 ( .a ({signal_2915, signal_1457}), .b ({signal_3050, signal_1592}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1578 ( .a ({signal_2916, signal_1458}), .b ({signal_3051, signal_1593}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1579 ( .a ({signal_2917, signal_1459}), .b ({signal_3052, signal_1594}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1580 ( .a ({signal_2918, signal_1460}), .b ({signal_3053, signal_1595}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1581 ( .a ({signal_2920, signal_1462}), .b ({signal_3054, signal_1596}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1582 ( .a ({signal_2921, signal_1463}), .b ({signal_3055, signal_1597}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1583 ( .a ({signal_2922, signal_1464}), .b ({signal_3056, signal_1598}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1584 ( .a ({signal_2923, signal_1465}), .b ({signal_3057, signal_1599}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1585 ( .a ({signal_2924, signal_1466}), .b ({signal_3058, signal_1600}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1586 ( .a ({signal_2925, signal_1467}), .b ({signal_3059, signal_1601}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1587 ( .a ({signal_2926, signal_1468}), .b ({signal_3060, signal_1602}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1588 ( .a ({signal_2927, signal_1469}), .b ({signal_3061, signal_1603}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1589 ( .a ({signal_2928, signal_1470}), .b ({signal_3062, signal_1604}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1590 ( .a ({signal_2929, signal_1471}), .b ({signal_3063, signal_1605}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1591 ( .a ({signal_2930, signal_1472}), .b ({signal_3064, signal_1606}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1592 ( .a ({signal_2931, signal_1473}), .b ({signal_3065, signal_1607}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1593 ( .a ({signal_2932, signal_1474}), .b ({signal_3066, signal_1608}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1594 ( .a ({signal_2933, signal_1475}), .b ({signal_3067, signal_1609}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1595 ( .a ({signal_2934, signal_1476}), .b ({signal_3068, signal_1610}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1596 ( .a ({signal_2935, signal_1477}), .b ({signal_3069, signal_1611}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1597 ( .a ({signal_2937, signal_1479}), .b ({signal_3070, signal_1612}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1598 ( .a ({signal_2938, signal_1480}), .b ({signal_3071, signal_1613}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1599 ( .a ({signal_2939, signal_1481}), .b ({signal_3072, signal_1614}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1600 ( .a ({signal_2940, signal_1482}), .b ({signal_3073, signal_1615}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1601 ( .a ({signal_2941, signal_1483}), .b ({signal_3074, signal_1616}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1602 ( .a ({signal_2942, signal_1484}), .b ({signal_3075, signal_1617}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1603 ( .a ({signal_2943, signal_1485}), .b ({signal_3076, signal_1618}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1604 ( .a ({signal_2944, signal_1486}), .b ({signal_3077, signal_1619}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1605 ( .a ({signal_2945, signal_1487}), .b ({signal_3078, signal_1620}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1606 ( .a ({signal_2946, signal_1488}), .b ({signal_3079, signal_1621}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1607 ( .a ({signal_2947, signal_1489}), .b ({signal_3080, signal_1622}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1608 ( .a ({signal_2948, signal_1490}), .b ({signal_3081, signal_1623}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1609 ( .a ({signal_2949, signal_1491}), .b ({signal_3082, signal_1624}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1610 ( .a ({signal_2950, signal_1492}), .b ({signal_3083, signal_1625}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1611 ( .a ({signal_2951, signal_1493}), .b ({signal_3084, signal_1626}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1612 ( .a ({signal_2952, signal_1494}), .b ({signal_3085, signal_1627}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1613 ( .a ({signal_2953, signal_1495}), .b ({signal_3086, signal_1628}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1614 ( .a ({signal_2954, signal_1496}), .b ({signal_3087, signal_1629}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1615 ( .a ({signal_2955, signal_1497}), .b ({signal_3088, signal_1630}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1616 ( .a ({signal_2956, signal_1498}), .b ({signal_3089, signal_1631}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1617 ( .a ({signal_2957, signal_1499}), .b ({signal_3090, signal_1632}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1618 ( .a ({signal_2958, signal_1500}), .b ({signal_3091, signal_1633}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1619 ( .a ({signal_2959, signal_1501}), .b ({signal_3092, signal_1634}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1620 ( .a ({signal_2960, signal_1502}), .b ({signal_3093, signal_1635}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1621 ( .a ({signal_2961, signal_1503}), .b ({signal_3094, signal_1636}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1622 ( .a ({signal_2962, signal_1504}), .b ({signal_3095, signal_1637}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1623 ( .a ({signal_4988, signal_4986}), .b ({signal_2688, signal_1230}), .clk ( clk ), .r ( Fresh[368] ), .c ({signal_3096, signal_1638}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1624 ( .a ({signal_5004, signal_5002}), .b ({signal_2689, signal_1231}), .clk ( clk ), .r ( Fresh[369] ), .c ({signal_3097, signal_1639}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1625 ( .a ({signal_4932, signal_4930}), .b ({signal_2694, signal_1236}), .clk ( clk ), .r ( Fresh[370] ), .c ({signal_3098, signal_1640}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1626 ( .a ({signal_2693, signal_1235}), .b ({signal_2714, signal_1256}), .clk ( clk ), .r ( Fresh[371] ), .c ({signal_3099, signal_1641}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1627 ( .a ({signal_5008, signal_5006}), .b ({signal_2715, signal_1257}), .clk ( clk ), .r ( Fresh[372] ), .c ({signal_3100, signal_1642}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1628 ( .a ({signal_4996, signal_4994}), .b ({signal_2721, signal_1263}), .clk ( clk ), .r ( Fresh[373] ), .c ({signal_3101, signal_1643}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1629 ( .a ({signal_2708, signal_1250}), .b ({signal_2711, signal_1253}), .clk ( clk ), .r ( Fresh[374] ), .c ({signal_3102, signal_1644}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1630 ( .a ({signal_2725, signal_1267}), .b ({signal_2726, signal_1268}), .clk ( clk ), .r ( Fresh[375] ), .c ({signal_3103, signal_1645}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1631 ( .a ({signal_5012, signal_5010}), .b ({signal_2698, signal_1240}), .clk ( clk ), .r ( Fresh[376] ), .c ({signal_3104, signal_1646}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1632 ( .a ({signal_2727, signal_1269}), .b ({signal_2728, signal_1270}), .clk ( clk ), .r ( Fresh[377] ), .c ({signal_3105, signal_1647}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1633 ( .a ({signal_2693, signal_1235}), .b ({signal_2713, signal_1255}), .clk ( clk ), .r ( Fresh[378] ), .c ({signal_3106, signal_1648}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1634 ( .a ({signal_2731, signal_1273}), .b ({signal_2732, signal_1274}), .clk ( clk ), .r ( Fresh[379] ), .c ({signal_3107, signal_1649}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1635 ( .a ({signal_2513, signal_1055}), .b ({signal_2712, signal_1254}), .clk ( clk ), .r ( Fresh[380] ), .c ({signal_3108, signal_1650}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1636 ( .a ({signal_5000, signal_4998}), .b ({signal_2699, signal_1241}), .clk ( clk ), .r ( Fresh[381] ), .c ({signal_3109, signal_1651}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1637 ( .a ({signal_2694, signal_1236}), .b ({signal_2517, signal_1059}), .clk ( clk ), .r ( Fresh[382] ), .c ({signal_3110, signal_1652}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1638 ( .a ({signal_2738, signal_1280}), .b ({signal_2739, signal_1281}), .clk ( clk ), .r ( Fresh[383] ), .c ({signal_3111, signal_1653}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1639 ( .a ({signal_2741, signal_1283}), .b ({signal_2742, signal_1284}), .clk ( clk ), .r ( Fresh[384] ), .c ({signal_3112, signal_1654}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1640 ( .a ({signal_2691, signal_1233}), .b ({signal_2744, signal_1286}), .clk ( clk ), .r ( Fresh[385] ), .c ({signal_3113, signal_1655}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1641 ( .a ({signal_2695, signal_1237}), .b ({signal_2746, signal_1288}), .clk ( clk ), .r ( Fresh[386] ), .c ({signal_3114, signal_1656}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1642 ( .a ({signal_2517, signal_1059}), .b ({signal_2696, signal_1238}), .clk ( clk ), .r ( Fresh[387] ), .c ({signal_3115, signal_1657}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1643 ( .a ({signal_2700, signal_1242}), .b ({signal_2701, signal_1243}), .clk ( clk ), .r ( Fresh[388] ), .c ({signal_3116, signal_1658}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1645 ( .a ({signal_2752, signal_1294}), .b ({signal_2753, signal_1295}), .clk ( clk ), .r ( Fresh[389] ), .c ({signal_3118, signal_1660}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1646 ( .a ({signal_2696, signal_1238}), .b ({signal_2760, signal_1302}), .clk ( clk ), .r ( Fresh[390] ), .c ({signal_3119, signal_1661}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1647 ( .a ({signal_5016, signal_5014}), .b ({signal_2764, signal_1306}), .clk ( clk ), .r ( Fresh[391] ), .c ({signal_3120, signal_1662}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1648 ( .a ({signal_2710, signal_1252}), .b ({signal_2768, signal_1310}), .clk ( clk ), .r ( Fresh[392] ), .c ({signal_3121, signal_1663}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1649 ( .a ({signal_5020, signal_5018}), .b ({signal_2841, signal_1383}), .clk ( clk ), .r ( Fresh[393] ), .c ({signal_3122, signal_1664}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1650 ( .a ({signal_4804, signal_4800}), .b ({signal_2755, signal_1297}), .clk ( clk ), .r ( Fresh[394] ), .c ({signal_3123, signal_1665}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1651 ( .a ({signal_2702, signal_1244}), .b ({signal_2769, signal_1311}), .clk ( clk ), .r ( Fresh[395] ), .c ({signal_3124, signal_1666}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1653 ( .a ({signal_2834, signal_1376}), .b ({signal_2775, signal_1317}), .clk ( clk ), .r ( Fresh[396] ), .c ({signal_3126, signal_1668}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1654 ( .a ({signal_2693, signal_1235}), .b ({signal_2777, signal_1319}), .clk ( clk ), .r ( Fresh[397] ), .c ({signal_3127, signal_1669}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1655 ( .a ({signal_2848, signal_1390}), .b ({signal_2523, signal_1065}), .clk ( clk ), .r ( Fresh[398] ), .c ({signal_3128, signal_1670}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1656 ( .a ({signal_4912, signal_4910}), .b ({signal_2778, signal_1320}), .clk ( clk ), .r ( Fresh[399] ), .c ({signal_3129, signal_1671}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1657 ( .a ({signal_2718, signal_1260}), .b ({signal_2758, signal_1300}), .clk ( clk ), .r ( Fresh[400] ), .c ({signal_3130, signal_1672}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1658 ( .a ({signal_4912, signal_4910}), .b ({signal_2779, signal_1321}), .clk ( clk ), .r ( Fresh[401] ), .c ({signal_3131, signal_1673}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1659 ( .a ({signal_2774, signal_1316}), .b ({signal_2780, signal_1322}), .clk ( clk ), .r ( Fresh[402] ), .c ({signal_3132, signal_1674}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1660 ( .a ({signal_2521, signal_1063}), .b ({signal_2781, signal_1323}), .clk ( clk ), .r ( Fresh[403] ), .c ({signal_3133, signal_1675}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1661 ( .a ({signal_2782, signal_1324}), .b ({signal_2783, signal_1325}), .clk ( clk ), .r ( Fresh[404] ), .c ({signal_3134, signal_1676}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1663 ( .a ({signal_2698, signal_1240}), .b ({signal_2755, signal_1297}), .clk ( clk ), .r ( Fresh[405] ), .c ({signal_3136, signal_1678}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1664 ( .a ({signal_2722, signal_1264}), .b ({signal_2789, signal_1331}), .clk ( clk ), .r ( Fresh[406] ), .c ({signal_3137, signal_1679}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1665 ( .a ({signal_2700, signal_1242}), .b ({signal_2790, signal_1332}), .clk ( clk ), .r ( Fresh[407] ), .c ({signal_3138, signal_1680}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1666 ( .a ({signal_2724, signal_1266}), .b ({signal_2792, signal_1334}), .clk ( clk ), .r ( Fresh[408] ), .c ({signal_3139, signal_1681}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1667 ( .a ({signal_2755, signal_1297}), .b ({signal_2795, signal_1337}), .clk ( clk ), .r ( Fresh[409] ), .c ({signal_3140, signal_1682}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1668 ( .a ({signal_2729, signal_1271}), .b ({signal_2789, signal_1331}), .clk ( clk ), .r ( Fresh[410] ), .c ({signal_3141, signal_1683}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1669 ( .a ({signal_4848, signal_4846}), .b ({signal_2778, signal_1320}), .clk ( clk ), .r ( Fresh[411] ), .c ({signal_3142, signal_1684}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1670 ( .a ({signal_2747, signal_1289}), .b ({signal_2798, signal_1340}), .clk ( clk ), .r ( Fresh[412] ), .c ({signal_3143, signal_1685}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1671 ( .a ({signal_5024, signal_5022}), .b ({signal_2799, signal_1341}), .clk ( clk ), .r ( Fresh[413] ), .c ({signal_3144, signal_1686}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1673 ( .a ({signal_2734, signal_1276}), .b ({signal_2788, signal_1330}), .clk ( clk ), .r ( Fresh[414] ), .c ({signal_3146, signal_1688}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1674 ( .a ({signal_2776, signal_1318}), .b ({signal_2876, signal_1418}), .clk ( clk ), .r ( Fresh[415] ), .c ({signal_3147, signal_1689}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1675 ( .a ({signal_2717, signal_1259}), .b ({signal_2782, signal_1324}), .clk ( clk ), .r ( Fresh[416] ), .c ({signal_3148, signal_1690}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1676 ( .a ({signal_2735, signal_1277}), .b ({signal_2804, signal_1346}), .clk ( clk ), .r ( Fresh[417] ), .c ({signal_3149, signal_1691}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1677 ( .a ({signal_2805, signal_1347}), .b ({signal_2806, signal_1348}), .clk ( clk ), .r ( Fresh[418] ), .c ({signal_3150, signal_1692}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1678 ( .a ({signal_2708, signal_1250}), .b ({signal_2807, signal_1349}), .clk ( clk ), .r ( Fresh[419] ), .c ({signal_3151, signal_1693}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1679 ( .a ({signal_2809, signal_1351}), .b ({signal_2810, signal_1352}), .clk ( clk ), .r ( Fresh[420] ), .c ({signal_3152, signal_1694}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1680 ( .a ({signal_2693, signal_1235}), .b ({signal_2767, signal_1309}), .clk ( clk ), .r ( Fresh[421] ), .c ({signal_3153, signal_1695}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1681 ( .a ({signal_2813, signal_1355}), .b ({signal_2814, signal_1356}), .clk ( clk ), .r ( Fresh[422] ), .c ({signal_3154, signal_1696}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1682 ( .a ({signal_2773, signal_1315}), .b ({signal_2815, signal_1357}), .clk ( clk ), .r ( Fresh[423] ), .c ({signal_3155, signal_1697}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1684 ( .a ({signal_2747, signal_1289}), .b ({signal_2748, signal_1290}), .clk ( clk ), .r ( Fresh[424] ), .c ({signal_3157, signal_1699}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1687 ( .a ({signal_2701, signal_1243}), .b ({signal_2748, signal_1290}), .clk ( clk ), .r ( Fresh[425] ), .c ({signal_3160, signal_1702}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1693 ( .a ({signal_2748, signal_1290}), .b ({signal_2763, signal_1305}), .clk ( clk ), .r ( Fresh[426] ), .c ({signal_3166, signal_1708}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1698 ( .a ({signal_2751, signal_1293}), .b ({signal_2822, signal_1364}), .clk ( clk ), .r ( Fresh[427] ), .c ({signal_3171, signal_1713}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1700 ( .a ({signal_3096, signal_1638}), .b ({signal_3173, signal_1715}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1701 ( .a ({signal_3097, signal_1639}), .b ({signal_3174, signal_1716}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1702 ( .a ({signal_3099, signal_1641}), .b ({signal_3175, signal_1717}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1703 ( .a ({signal_3100, signal_1642}), .b ({signal_3176, signal_1718}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1704 ( .a ({signal_3101, signal_1643}), .b ({signal_3177, signal_1719}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1705 ( .a ({signal_3102, signal_1644}), .b ({signal_3178, signal_1720}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1706 ( .a ({signal_3104, signal_1646}), .b ({signal_3179, signal_1721}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1707 ( .a ({signal_3105, signal_1647}), .b ({signal_3180, signal_1722}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1708 ( .a ({signal_3106, signal_1648}), .b ({signal_3181, signal_1723}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1709 ( .a ({signal_3108, signal_1650}), .b ({signal_3182, signal_1724}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1710 ( .a ({signal_3109, signal_1651}), .b ({signal_3183, signal_1725}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1711 ( .a ({signal_3110, signal_1652}), .b ({signal_3184, signal_1726}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1712 ( .a ({signal_3114, signal_1656}), .b ({signal_3185, signal_1727}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1713 ( .a ({signal_3115, signal_1657}), .b ({signal_3186, signal_1728}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1714 ( .a ({signal_3116, signal_1658}), .b ({signal_3187, signal_1729}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1716 ( .a ({signal_3120, signal_1662}), .b ({signal_3189, signal_1731}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1717 ( .a ({signal_3121, signal_1663}), .b ({signal_3190, signal_1732}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1718 ( .a ({signal_3122, signal_1664}), .b ({signal_3191, signal_1733}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1719 ( .a ({signal_3123, signal_1665}), .b ({signal_3192, signal_1734}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1720 ( .a ({signal_3124, signal_1666}), .b ({signal_3193, signal_1735}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1722 ( .a ({signal_3127, signal_1669}), .b ({signal_3195, signal_1737}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1723 ( .a ({signal_3131, signal_1673}), .b ({signal_3196, signal_1738}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1724 ( .a ({signal_3134, signal_1676}), .b ({signal_3197, signal_1739}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1726 ( .a ({signal_3136, signal_1678}), .b ({signal_3199, signal_1741}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1727 ( .a ({signal_3137, signal_1679}), .b ({signal_3200, signal_1742}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1728 ( .a ({signal_3138, signal_1680}), .b ({signal_3201, signal_1743}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1729 ( .a ({signal_3139, signal_1681}), .b ({signal_3202, signal_1744}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1730 ( .a ({signal_3140, signal_1682}), .b ({signal_3203, signal_1745}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1731 ( .a ({signal_3144, signal_1686}), .b ({signal_3204, signal_1746}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1732 ( .a ({signal_3147, signal_1689}), .b ({signal_3205, signal_1747}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1733 ( .a ({signal_3151, signal_1693}), .b ({signal_3206, signal_1748}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1734 ( .a ({signal_3154, signal_1696}), .b ({signal_3207, signal_1749}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1735 ( .a ({signal_3155, signal_1697}), .b ({signal_3208, signal_1750}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1736 ( .a ({signal_3157, signal_1699}), .b ({signal_3209, signal_1751}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1739 ( .a ({signal_3160, signal_1702}), .b ({signal_3212, signal_1754}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1745 ( .a ({signal_3166, signal_1708}), .b ({signal_3218, signal_1760}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1749 ( .a ({signal_3171, signal_1713}), .b ({signal_3222, signal_1764}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1751 ( .a ({signal_2560, signal_1102}), .b ({signal_2965, signal_1507}), .clk ( clk ), .r ( Fresh[428] ), .c ({signal_3224, signal_1766}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1753 ( .a ({signal_4948, signal_4944}), .b ({signal_2966, signal_1508}), .clk ( clk ), .r ( Fresh[429] ), .c ({signal_3226, signal_1768}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1754 ( .a ({signal_4900, signal_4898}), .b ({signal_2967, signal_1509}), .clk ( clk ), .r ( Fresh[430] ), .c ({signal_3227, signal_1769}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1755 ( .a ({signal_2541, signal_1083}), .b ({signal_2968, signal_1510}), .clk ( clk ), .r ( Fresh[431] ), .c ({signal_3228, signal_1770}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1756 ( .a ({signal_4940, signal_4938}), .b ({signal_2965, signal_1507}), .clk ( clk ), .r ( Fresh[432] ), .c ({signal_3229, signal_1771}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1757 ( .a ({signal_2590, signal_1132}), .b ({signal_2969, signal_1511}), .clk ( clk ), .r ( Fresh[433] ), .c ({signal_3230, signal_1772}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1758 ( .a ({signal_4992, signal_4990}), .b ({signal_2969, signal_1511}), .clk ( clk ), .r ( Fresh[434] ), .c ({signal_3231, signal_1773}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1760 ( .a ({signal_5028, signal_5026}), .b ({signal_2972, signal_1514}), .clk ( clk ), .r ( Fresh[435] ), .c ({signal_3233, signal_1775}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1761 ( .a ({signal_5032, signal_5030}), .b ({signal_2973, signal_1515}), .clk ( clk ), .r ( Fresh[436] ), .c ({signal_3234, signal_1776}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1762 ( .a ({signal_4820, signal_4818}), .b ({signal_2974, signal_1516}), .clk ( clk ), .r ( Fresh[437] ), .c ({signal_3235, signal_1777}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1764 ( .a ({signal_4920, signal_4918}), .b ({signal_2977, signal_1519}), .clk ( clk ), .r ( Fresh[438] ), .c ({signal_3237, signal_1779}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1765 ( .a ({signal_5016, signal_5014}), .b ({signal_2978, signal_1520}), .clk ( clk ), .r ( Fresh[439] ), .c ({signal_3238, signal_1780}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1766 ( .a ({signal_4832, signal_4830}), .b ({signal_2979, signal_1521}), .clk ( clk ), .r ( Fresh[440] ), .c ({signal_3239, signal_1781}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1767 ( .a ({signal_4872, signal_4870}), .b ({signal_2980, signal_1522}), .clk ( clk ), .r ( Fresh[441] ), .c ({signal_3240, signal_1782}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1769 ( .a ({signal_2536, signal_1078}), .b ({signal_2980, signal_1522}), .clk ( clk ), .r ( Fresh[442] ), .c ({signal_3242, signal_1784}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1770 ( .a ({signal_2543, signal_1085}), .b ({signal_2986, signal_1528}), .clk ( clk ), .r ( Fresh[443] ), .c ({signal_3243, signal_1785}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1772 ( .a ({signal_4852, signal_4850}), .b ({signal_2979, signal_1521}), .clk ( clk ), .r ( Fresh[444] ), .c ({signal_3245, signal_1787}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1773 ( .a ({signal_2611, signal_1153}), .b ({signal_2993, signal_1535}), .clk ( clk ), .r ( Fresh[445] ), .c ({signal_3246, signal_1788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1776 ( .a ({signal_4968, signal_4966}), .b ({signal_2978, signal_1520}), .clk ( clk ), .r ( Fresh[446] ), .c ({signal_3249, signal_1791}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1778 ( .a ({signal_5036, signal_5034}), .b ({signal_3005, signal_1547}), .clk ( clk ), .r ( Fresh[447] ), .c ({signal_3251, signal_1793}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1779 ( .a ({signal_2544, signal_1086}), .b ({signal_3006, signal_1548}), .clk ( clk ), .r ( Fresh[448] ), .c ({signal_3252, signal_1794}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1782 ( .a ({signal_4912, signal_4910}), .b ({signal_3011, signal_1553}), .clk ( clk ), .r ( Fresh[449] ), .c ({signal_3255, signal_1797}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1783 ( .a ({signal_4828, signal_4826}), .b ({signal_3012, signal_1554}), .clk ( clk ), .r ( Fresh[450] ), .c ({signal_3256, signal_1798}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1784 ( .a ({signal_2540, signal_1082}), .b ({signal_2973, signal_1515}), .clk ( clk ), .r ( Fresh[451] ), .c ({signal_3257, signal_1799}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1785 ( .a ({signal_4960, signal_4958}), .b ({signal_3016, signal_1558}), .clk ( clk ), .r ( Fresh[452] ), .c ({signal_3258, signal_1800}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1786 ( .a ({signal_4912, signal_4910}), .b ({signal_3017, signal_1559}), .clk ( clk ), .r ( Fresh[453] ), .c ({signal_3259, signal_1801}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1835 ( .a ({signal_3224, signal_1766}), .b ({signal_3308, signal_1850}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1836 ( .a ({signal_3228, signal_1770}), .b ({signal_3309, signal_1851}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1837 ( .a ({signal_3230, signal_1772}), .b ({signal_3310, signal_1852}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1838 ( .a ({signal_3231, signal_1773}), .b ({signal_3311, signal_1853}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1839 ( .a ({signal_3233, signal_1775}), .b ({signal_3312, signal_1854}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1840 ( .a ({signal_3234, signal_1776}), .b ({signal_3313, signal_1855}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1841 ( .a ({signal_3235, signal_1777}), .b ({signal_3314, signal_1856}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1843 ( .a ({signal_3237, signal_1779}), .b ({signal_3316, signal_1858}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1844 ( .a ({signal_3238, signal_1780}), .b ({signal_3317, signal_1859}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1845 ( .a ({signal_3239, signal_1781}), .b ({signal_3318, signal_1860}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1846 ( .a ({signal_3242, signal_1784}), .b ({signal_3319, signal_1861}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1847 ( .a ({signal_3243, signal_1785}), .b ({signal_3320, signal_1862}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1848 ( .a ({signal_3245, signal_1787}), .b ({signal_3321, signal_1863}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1849 ( .a ({signal_3246, signal_1788}), .b ({signal_3322, signal_1864}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1850 ( .a ({signal_3249, signal_1791}), .b ({signal_3323, signal_1865}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1851 ( .a ({signal_3251, signal_1793}), .b ({signal_3324, signal_1866}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1852 ( .a ({signal_3252, signal_1794}), .b ({signal_3325, signal_1867}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1854 ( .a ({signal_3255, signal_1797}), .b ({signal_3327, signal_1869}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1855 ( .a ({signal_3256, signal_1798}), .b ({signal_3328, signal_1870}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1856 ( .a ({signal_3257, signal_1799}), .b ({signal_3329, signal_1871}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1857 ( .a ({signal_3258, signal_1800}), .b ({signal_3330, signal_1872}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1858 ( .a ({signal_3259, signal_1801}), .b ({signal_3331, signal_1873}) ) ;
    buf_clk cell_2678 ( .C ( clk ), .D ( signal_5037 ), .Q ( signal_5038 ) ) ;
    buf_clk cell_2680 ( .C ( clk ), .D ( signal_5039 ), .Q ( signal_5040 ) ) ;
    buf_clk cell_2682 ( .C ( clk ), .D ( signal_5041 ), .Q ( signal_5042 ) ) ;
    buf_clk cell_2684 ( .C ( clk ), .D ( signal_5043 ), .Q ( signal_5044 ) ) ;
    buf_clk cell_2686 ( .C ( clk ), .D ( signal_5045 ), .Q ( signal_5046 ) ) ;
    buf_clk cell_2688 ( .C ( clk ), .D ( signal_5047 ), .Q ( signal_5048 ) ) ;
    buf_clk cell_2690 ( .C ( clk ), .D ( signal_5049 ), .Q ( signal_5050 ) ) ;
    buf_clk cell_2692 ( .C ( clk ), .D ( signal_5051 ), .Q ( signal_5052 ) ) ;
    buf_clk cell_2694 ( .C ( clk ), .D ( signal_5053 ), .Q ( signal_5054 ) ) ;
    buf_clk cell_2696 ( .C ( clk ), .D ( signal_5055 ), .Q ( signal_5056 ) ) ;
    buf_clk cell_2698 ( .C ( clk ), .D ( signal_5057 ), .Q ( signal_5058 ) ) ;
    buf_clk cell_2700 ( .C ( clk ), .D ( signal_5059 ), .Q ( signal_5060 ) ) ;
    buf_clk cell_2702 ( .C ( clk ), .D ( signal_5061 ), .Q ( signal_5062 ) ) ;
    buf_clk cell_2704 ( .C ( clk ), .D ( signal_5063 ), .Q ( signal_5064 ) ) ;
    buf_clk cell_2706 ( .C ( clk ), .D ( signal_5065 ), .Q ( signal_5066 ) ) ;
    buf_clk cell_2708 ( .C ( clk ), .D ( signal_5067 ), .Q ( signal_5068 ) ) ;
    buf_clk cell_2710 ( .C ( clk ), .D ( signal_5069 ), .Q ( signal_5070 ) ) ;
    buf_clk cell_2712 ( .C ( clk ), .D ( signal_5071 ), .Q ( signal_5072 ) ) ;
    buf_clk cell_2714 ( .C ( clk ), .D ( signal_5073 ), .Q ( signal_5074 ) ) ;
    buf_clk cell_2716 ( .C ( clk ), .D ( signal_5075 ), .Q ( signal_5076 ) ) ;
    buf_clk cell_2718 ( .C ( clk ), .D ( signal_5077 ), .Q ( signal_5078 ) ) ;
    buf_clk cell_2720 ( .C ( clk ), .D ( signal_5079 ), .Q ( signal_5080 ) ) ;
    buf_clk cell_2726 ( .C ( clk ), .D ( signal_5085 ), .Q ( signal_5086 ) ) ;
    buf_clk cell_2732 ( .C ( clk ), .D ( signal_5091 ), .Q ( signal_5092 ) ) ;
    buf_clk cell_2734 ( .C ( clk ), .D ( signal_5093 ), .Q ( signal_5094 ) ) ;
    buf_clk cell_2736 ( .C ( clk ), .D ( signal_5095 ), .Q ( signal_5096 ) ) ;
    buf_clk cell_2738 ( .C ( clk ), .D ( signal_5097 ), .Q ( signal_5098 ) ) ;
    buf_clk cell_2740 ( .C ( clk ), .D ( signal_5099 ), .Q ( signal_5100 ) ) ;
    buf_clk cell_2742 ( .C ( clk ), .D ( signal_5101 ), .Q ( signal_5102 ) ) ;
    buf_clk cell_2744 ( .C ( clk ), .D ( signal_5103 ), .Q ( signal_5104 ) ) ;
    buf_clk cell_2746 ( .C ( clk ), .D ( signal_5105 ), .Q ( signal_5106 ) ) ;
    buf_clk cell_2748 ( .C ( clk ), .D ( signal_5107 ), .Q ( signal_5108 ) ) ;
    buf_clk cell_2750 ( .C ( clk ), .D ( signal_5109 ), .Q ( signal_5110 ) ) ;
    buf_clk cell_2752 ( .C ( clk ), .D ( signal_5111 ), .Q ( signal_5112 ) ) ;
    buf_clk cell_2754 ( .C ( clk ), .D ( signal_5113 ), .Q ( signal_5114 ) ) ;
    buf_clk cell_2756 ( .C ( clk ), .D ( signal_5115 ), .Q ( signal_5116 ) ) ;
    buf_clk cell_2758 ( .C ( clk ), .D ( signal_5117 ), .Q ( signal_5118 ) ) ;
    buf_clk cell_2760 ( .C ( clk ), .D ( signal_5119 ), .Q ( signal_5120 ) ) ;
    buf_clk cell_2762 ( .C ( clk ), .D ( signal_5121 ), .Q ( signal_5122 ) ) ;
    buf_clk cell_2764 ( .C ( clk ), .D ( signal_5123 ), .Q ( signal_5124 ) ) ;
    buf_clk cell_2766 ( .C ( clk ), .D ( signal_5125 ), .Q ( signal_5126 ) ) ;
    buf_clk cell_2768 ( .C ( clk ), .D ( signal_5127 ), .Q ( signal_5128 ) ) ;
    buf_clk cell_2770 ( .C ( clk ), .D ( signal_5129 ), .Q ( signal_5130 ) ) ;
    buf_clk cell_2772 ( .C ( clk ), .D ( signal_5131 ), .Q ( signal_5132 ) ) ;
    buf_clk cell_2774 ( .C ( clk ), .D ( signal_5133 ), .Q ( signal_5134 ) ) ;
    buf_clk cell_2776 ( .C ( clk ), .D ( signal_5135 ), .Q ( signal_5136 ) ) ;
    buf_clk cell_2778 ( .C ( clk ), .D ( signal_5137 ), .Q ( signal_5138 ) ) ;
    buf_clk cell_2780 ( .C ( clk ), .D ( signal_5139 ), .Q ( signal_5140 ) ) ;
    buf_clk cell_2782 ( .C ( clk ), .D ( signal_5141 ), .Q ( signal_5142 ) ) ;
    buf_clk cell_2784 ( .C ( clk ), .D ( signal_5143 ), .Q ( signal_5144 ) ) ;
    buf_clk cell_2786 ( .C ( clk ), .D ( signal_5145 ), .Q ( signal_5146 ) ) ;
    buf_clk cell_2788 ( .C ( clk ), .D ( signal_5147 ), .Q ( signal_5148 ) ) ;
    buf_clk cell_2790 ( .C ( clk ), .D ( signal_5149 ), .Q ( signal_5150 ) ) ;
    buf_clk cell_2792 ( .C ( clk ), .D ( signal_5151 ), .Q ( signal_5152 ) ) ;
    buf_clk cell_2794 ( .C ( clk ), .D ( signal_5153 ), .Q ( signal_5154 ) ) ;
    buf_clk cell_2796 ( .C ( clk ), .D ( signal_5155 ), .Q ( signal_5156 ) ) ;
    buf_clk cell_2798 ( .C ( clk ), .D ( signal_5157 ), .Q ( signal_5158 ) ) ;
    buf_clk cell_2800 ( .C ( clk ), .D ( signal_5159 ), .Q ( signal_5160 ) ) ;
    buf_clk cell_2802 ( .C ( clk ), .D ( signal_5161 ), .Q ( signal_5162 ) ) ;
    buf_clk cell_2804 ( .C ( clk ), .D ( signal_5163 ), .Q ( signal_5164 ) ) ;
    buf_clk cell_2806 ( .C ( clk ), .D ( signal_5165 ), .Q ( signal_5166 ) ) ;
    buf_clk cell_2808 ( .C ( clk ), .D ( signal_5167 ), .Q ( signal_5168 ) ) ;
    buf_clk cell_2810 ( .C ( clk ), .D ( signal_5169 ), .Q ( signal_5170 ) ) ;
    buf_clk cell_2812 ( .C ( clk ), .D ( signal_5171 ), .Q ( signal_5172 ) ) ;
    buf_clk cell_2816 ( .C ( clk ), .D ( signal_5175 ), .Q ( signal_5176 ) ) ;
    buf_clk cell_2820 ( .C ( clk ), .D ( signal_5179 ), .Q ( signal_5180 ) ) ;
    buf_clk cell_2822 ( .C ( clk ), .D ( signal_5181 ), .Q ( signal_5182 ) ) ;
    buf_clk cell_2824 ( .C ( clk ), .D ( signal_5183 ), .Q ( signal_5184 ) ) ;
    buf_clk cell_2826 ( .C ( clk ), .D ( signal_5185 ), .Q ( signal_5186 ) ) ;
    buf_clk cell_2828 ( .C ( clk ), .D ( signal_5187 ), .Q ( signal_5188 ) ) ;
    buf_clk cell_2832 ( .C ( clk ), .D ( signal_5191 ), .Q ( signal_5192 ) ) ;
    buf_clk cell_2836 ( .C ( clk ), .D ( signal_5195 ), .Q ( signal_5196 ) ) ;
    buf_clk cell_2838 ( .C ( clk ), .D ( signal_5197 ), .Q ( signal_5198 ) ) ;
    buf_clk cell_2840 ( .C ( clk ), .D ( signal_5199 ), .Q ( signal_5200 ) ) ;
    buf_clk cell_2842 ( .C ( clk ), .D ( signal_5201 ), .Q ( signal_5202 ) ) ;
    buf_clk cell_2844 ( .C ( clk ), .D ( signal_5203 ), .Q ( signal_5204 ) ) ;
    buf_clk cell_2846 ( .C ( clk ), .D ( signal_5205 ), .Q ( signal_5206 ) ) ;
    buf_clk cell_2848 ( .C ( clk ), .D ( signal_5207 ), .Q ( signal_5208 ) ) ;
    buf_clk cell_2850 ( .C ( clk ), .D ( signal_5209 ), .Q ( signal_5210 ) ) ;
    buf_clk cell_2852 ( .C ( clk ), .D ( signal_5211 ), .Q ( signal_5212 ) ) ;
    buf_clk cell_2854 ( .C ( clk ), .D ( signal_5213 ), .Q ( signal_5214 ) ) ;
    buf_clk cell_2856 ( .C ( clk ), .D ( signal_5215 ), .Q ( signal_5216 ) ) ;
    buf_clk cell_2858 ( .C ( clk ), .D ( signal_5217 ), .Q ( signal_5218 ) ) ;
    buf_clk cell_2860 ( .C ( clk ), .D ( signal_5219 ), .Q ( signal_5220 ) ) ;
    buf_clk cell_2862 ( .C ( clk ), .D ( signal_5221 ), .Q ( signal_5222 ) ) ;
    buf_clk cell_2864 ( .C ( clk ), .D ( signal_5223 ), .Q ( signal_5224 ) ) ;
    buf_clk cell_2866 ( .C ( clk ), .D ( signal_5225 ), .Q ( signal_5226 ) ) ;
    buf_clk cell_2868 ( .C ( clk ), .D ( signal_5227 ), .Q ( signal_5228 ) ) ;
    buf_clk cell_2870 ( .C ( clk ), .D ( signal_5229 ), .Q ( signal_5230 ) ) ;
    buf_clk cell_2872 ( .C ( clk ), .D ( signal_5231 ), .Q ( signal_5232 ) ) ;
    buf_clk cell_2874 ( .C ( clk ), .D ( signal_5233 ), .Q ( signal_5234 ) ) ;
    buf_clk cell_2876 ( .C ( clk ), .D ( signal_5235 ), .Q ( signal_5236 ) ) ;
    buf_clk cell_2878 ( .C ( clk ), .D ( signal_5237 ), .Q ( signal_5238 ) ) ;
    buf_clk cell_2880 ( .C ( clk ), .D ( signal_5239 ), .Q ( signal_5240 ) ) ;
    buf_clk cell_2884 ( .C ( clk ), .D ( signal_5243 ), .Q ( signal_5244 ) ) ;
    buf_clk cell_2888 ( .C ( clk ), .D ( signal_5247 ), .Q ( signal_5248 ) ) ;
    buf_clk cell_2890 ( .C ( clk ), .D ( signal_5249 ), .Q ( signal_5250 ) ) ;
    buf_clk cell_2892 ( .C ( clk ), .D ( signal_5251 ), .Q ( signal_5252 ) ) ;
    buf_clk cell_2896 ( .C ( clk ), .D ( signal_5255 ), .Q ( signal_5256 ) ) ;
    buf_clk cell_2900 ( .C ( clk ), .D ( signal_5259 ), .Q ( signal_5260 ) ) ;
    buf_clk cell_2902 ( .C ( clk ), .D ( signal_5261 ), .Q ( signal_5262 ) ) ;
    buf_clk cell_2904 ( .C ( clk ), .D ( signal_5263 ), .Q ( signal_5264 ) ) ;
    buf_clk cell_2906 ( .C ( clk ), .D ( signal_5265 ), .Q ( signal_5266 ) ) ;
    buf_clk cell_2908 ( .C ( clk ), .D ( signal_5267 ), .Q ( signal_5268 ) ) ;
    buf_clk cell_2910 ( .C ( clk ), .D ( signal_5269 ), .Q ( signal_5270 ) ) ;
    buf_clk cell_2912 ( .C ( clk ), .D ( signal_5271 ), .Q ( signal_5272 ) ) ;
    buf_clk cell_2918 ( .C ( clk ), .D ( signal_5277 ), .Q ( signal_5278 ) ) ;
    buf_clk cell_2924 ( .C ( clk ), .D ( signal_5283 ), .Q ( signal_5284 ) ) ;
    buf_clk cell_2926 ( .C ( clk ), .D ( signal_5285 ), .Q ( signal_5286 ) ) ;
    buf_clk cell_2928 ( .C ( clk ), .D ( signal_5287 ), .Q ( signal_5288 ) ) ;
    buf_clk cell_2930 ( .C ( clk ), .D ( signal_5289 ), .Q ( signal_5290 ) ) ;
    buf_clk cell_2932 ( .C ( clk ), .D ( signal_5291 ), .Q ( signal_5292 ) ) ;
    buf_clk cell_2934 ( .C ( clk ), .D ( signal_5293 ), .Q ( signal_5294 ) ) ;
    buf_clk cell_2936 ( .C ( clk ), .D ( signal_5295 ), .Q ( signal_5296 ) ) ;
    buf_clk cell_2938 ( .C ( clk ), .D ( signal_5297 ), .Q ( signal_5298 ) ) ;
    buf_clk cell_2940 ( .C ( clk ), .D ( signal_5299 ), .Q ( signal_5300 ) ) ;
    buf_clk cell_2944 ( .C ( clk ), .D ( signal_5303 ), .Q ( signal_5304 ) ) ;
    buf_clk cell_2948 ( .C ( clk ), .D ( signal_5307 ), .Q ( signal_5308 ) ) ;
    buf_clk cell_2950 ( .C ( clk ), .D ( signal_5309 ), .Q ( signal_5310 ) ) ;
    buf_clk cell_2952 ( .C ( clk ), .D ( signal_5311 ), .Q ( signal_5312 ) ) ;
    buf_clk cell_2954 ( .C ( clk ), .D ( signal_5313 ), .Q ( signal_5314 ) ) ;
    buf_clk cell_2956 ( .C ( clk ), .D ( signal_5315 ), .Q ( signal_5316 ) ) ;
    buf_clk cell_2958 ( .C ( clk ), .D ( signal_5317 ), .Q ( signal_5318 ) ) ;
    buf_clk cell_2960 ( .C ( clk ), .D ( signal_5319 ), .Q ( signal_5320 ) ) ;
    buf_clk cell_2962 ( .C ( clk ), .D ( signal_5321 ), .Q ( signal_5322 ) ) ;
    buf_clk cell_2964 ( .C ( clk ), .D ( signal_5323 ), .Q ( signal_5324 ) ) ;
    buf_clk cell_2966 ( .C ( clk ), .D ( signal_5325 ), .Q ( signal_5326 ) ) ;
    buf_clk cell_2968 ( .C ( clk ), .D ( signal_5327 ), .Q ( signal_5328 ) ) ;
    buf_clk cell_2970 ( .C ( clk ), .D ( signal_5329 ), .Q ( signal_5330 ) ) ;
    buf_clk cell_2972 ( .C ( clk ), .D ( signal_5331 ), .Q ( signal_5332 ) ) ;
    buf_clk cell_2974 ( .C ( clk ), .D ( signal_5333 ), .Q ( signal_5334 ) ) ;
    buf_clk cell_2976 ( .C ( clk ), .D ( signal_5335 ), .Q ( signal_5336 ) ) ;
    buf_clk cell_2978 ( .C ( clk ), .D ( signal_5337 ), .Q ( signal_5338 ) ) ;
    buf_clk cell_2980 ( .C ( clk ), .D ( signal_5339 ), .Q ( signal_5340 ) ) ;
    buf_clk cell_2982 ( .C ( clk ), .D ( signal_5341 ), .Q ( signal_5342 ) ) ;
    buf_clk cell_2984 ( .C ( clk ), .D ( signal_5343 ), .Q ( signal_5344 ) ) ;
    buf_clk cell_2988 ( .C ( clk ), .D ( signal_5347 ), .Q ( signal_5348 ) ) ;
    buf_clk cell_2992 ( .C ( clk ), .D ( signal_5351 ), .Q ( signal_5352 ) ) ;
    buf_clk cell_2994 ( .C ( clk ), .D ( signal_5353 ), .Q ( signal_5354 ) ) ;
    buf_clk cell_2996 ( .C ( clk ), .D ( signal_5355 ), .Q ( signal_5356 ) ) ;
    buf_clk cell_2998 ( .C ( clk ), .D ( signal_5357 ), .Q ( signal_5358 ) ) ;
    buf_clk cell_3000 ( .C ( clk ), .D ( signal_5359 ), .Q ( signal_5360 ) ) ;
    buf_clk cell_3002 ( .C ( clk ), .D ( signal_5361 ), .Q ( signal_5362 ) ) ;
    buf_clk cell_3004 ( .C ( clk ), .D ( signal_5363 ), .Q ( signal_5364 ) ) ;
    buf_clk cell_3006 ( .C ( clk ), .D ( signal_5365 ), .Q ( signal_5366 ) ) ;
    buf_clk cell_3008 ( .C ( clk ), .D ( signal_5367 ), .Q ( signal_5368 ) ) ;
    buf_clk cell_3010 ( .C ( clk ), .D ( signal_5369 ), .Q ( signal_5370 ) ) ;
    buf_clk cell_3012 ( .C ( clk ), .D ( signal_5371 ), .Q ( signal_5372 ) ) ;
    buf_clk cell_3014 ( .C ( clk ), .D ( signal_5373 ), .Q ( signal_5374 ) ) ;
    buf_clk cell_3016 ( .C ( clk ), .D ( signal_5375 ), .Q ( signal_5376 ) ) ;
    buf_clk cell_3026 ( .C ( clk ), .D ( signal_5385 ), .Q ( signal_5386 ) ) ;
    buf_clk cell_3030 ( .C ( clk ), .D ( signal_5389 ), .Q ( signal_5390 ) ) ;
    buf_clk cell_3038 ( .C ( clk ), .D ( signal_5397 ), .Q ( signal_5398 ) ) ;
    buf_clk cell_3042 ( .C ( clk ), .D ( signal_5401 ), .Q ( signal_5402 ) ) ;
    buf_clk cell_3046 ( .C ( clk ), .D ( signal_5405 ), .Q ( signal_5406 ) ) ;
    buf_clk cell_3050 ( .C ( clk ), .D ( signal_5409 ), .Q ( signal_5410 ) ) ;
    buf_clk cell_3054 ( .C ( clk ), .D ( signal_5413 ), .Q ( signal_5414 ) ) ;
    buf_clk cell_3058 ( .C ( clk ), .D ( signal_5417 ), .Q ( signal_5418 ) ) ;
    buf_clk cell_3066 ( .C ( clk ), .D ( signal_5425 ), .Q ( signal_5426 ) ) ;
    buf_clk cell_3074 ( .C ( clk ), .D ( signal_5433 ), .Q ( signal_5434 ) ) ;
    buf_clk cell_3086 ( .C ( clk ), .D ( signal_5445 ), .Q ( signal_5446 ) ) ;
    buf_clk cell_3090 ( .C ( clk ), .D ( signal_5449 ), .Q ( signal_5450 ) ) ;
    buf_clk cell_3102 ( .C ( clk ), .D ( signal_5461 ), .Q ( signal_5462 ) ) ;
    buf_clk cell_3106 ( .C ( clk ), .D ( signal_5465 ), .Q ( signal_5466 ) ) ;
    buf_clk cell_3130 ( .C ( clk ), .D ( signal_5489 ), .Q ( signal_5490 ) ) ;
    buf_clk cell_3134 ( .C ( clk ), .D ( signal_5493 ), .Q ( signal_5494 ) ) ;
    buf_clk cell_3154 ( .C ( clk ), .D ( signal_5513 ), .Q ( signal_5514 ) ) ;
    buf_clk cell_3158 ( .C ( clk ), .D ( signal_5517 ), .Q ( signal_5518 ) ) ;
    buf_clk cell_3170 ( .C ( clk ), .D ( signal_5529 ), .Q ( signal_5530 ) ) ;
    buf_clk cell_3174 ( .C ( clk ), .D ( signal_5533 ), .Q ( signal_5534 ) ) ;
    buf_clk cell_3178 ( .C ( clk ), .D ( signal_5537 ), .Q ( signal_5538 ) ) ;
    buf_clk cell_3182 ( .C ( clk ), .D ( signal_5541 ), .Q ( signal_5542 ) ) ;
    buf_clk cell_3186 ( .C ( clk ), .D ( signal_5545 ), .Q ( signal_5546 ) ) ;
    buf_clk cell_3190 ( .C ( clk ), .D ( signal_5549 ), .Q ( signal_5550 ) ) ;
    buf_clk cell_3194 ( .C ( clk ), .D ( signal_5553 ), .Q ( signal_5554 ) ) ;
    buf_clk cell_3198 ( .C ( clk ), .D ( signal_5557 ), .Q ( signal_5558 ) ) ;
    buf_clk cell_3222 ( .C ( clk ), .D ( signal_5581 ), .Q ( signal_5582 ) ) ;
    buf_clk cell_3226 ( .C ( clk ), .D ( signal_5585 ), .Q ( signal_5586 ) ) ;
    buf_clk cell_3230 ( .C ( clk ), .D ( signal_5589 ), .Q ( signal_5590 ) ) ;
    buf_clk cell_3234 ( .C ( clk ), .D ( signal_5593 ), .Q ( signal_5594 ) ) ;
    buf_clk cell_3238 ( .C ( clk ), .D ( signal_5597 ), .Q ( signal_5598 ) ) ;
    buf_clk cell_3242 ( .C ( clk ), .D ( signal_5601 ), .Q ( signal_5602 ) ) ;
    buf_clk cell_3250 ( .C ( clk ), .D ( signal_5609 ), .Q ( signal_5610 ) ) ;
    buf_clk cell_3254 ( .C ( clk ), .D ( signal_5613 ), .Q ( signal_5614 ) ) ;
    buf_clk cell_3278 ( .C ( clk ), .D ( signal_5637 ), .Q ( signal_5638 ) ) ;
    buf_clk cell_3282 ( .C ( clk ), .D ( signal_5641 ), .Q ( signal_5642 ) ) ;
    buf_clk cell_3286 ( .C ( clk ), .D ( signal_5645 ), .Q ( signal_5646 ) ) ;
    buf_clk cell_3290 ( .C ( clk ), .D ( signal_5649 ), .Q ( signal_5650 ) ) ;
    buf_clk cell_3298 ( .C ( clk ), .D ( signal_5657 ), .Q ( signal_5658 ) ) ;
    buf_clk cell_3302 ( .C ( clk ), .D ( signal_5661 ), .Q ( signal_5662 ) ) ;
    buf_clk cell_3314 ( .C ( clk ), .D ( signal_5673 ), .Q ( signal_5674 ) ) ;
    buf_clk cell_3318 ( .C ( clk ), .D ( signal_5677 ), .Q ( signal_5678 ) ) ;
    buf_clk cell_3322 ( .C ( clk ), .D ( signal_5681 ), .Q ( signal_5682 ) ) ;
    buf_clk cell_3326 ( .C ( clk ), .D ( signal_5685 ), .Q ( signal_5686 ) ) ;
    buf_clk cell_3330 ( .C ( clk ), .D ( signal_5689 ), .Q ( signal_5690 ) ) ;
    buf_clk cell_3334 ( .C ( clk ), .D ( signal_5693 ), .Q ( signal_5694 ) ) ;
    buf_clk cell_3342 ( .C ( clk ), .D ( signal_5701 ), .Q ( signal_5702 ) ) ;
    buf_clk cell_3346 ( .C ( clk ), .D ( signal_5705 ), .Q ( signal_5706 ) ) ;
    buf_clk cell_3350 ( .C ( clk ), .D ( signal_5709 ), .Q ( signal_5710 ) ) ;
    buf_clk cell_3354 ( .C ( clk ), .D ( signal_5713 ), .Q ( signal_5714 ) ) ;
    buf_clk cell_3362 ( .C ( clk ), .D ( signal_5721 ), .Q ( signal_5722 ) ) ;
    buf_clk cell_3366 ( .C ( clk ), .D ( signal_5725 ), .Q ( signal_5726 ) ) ;
    buf_clk cell_3382 ( .C ( clk ), .D ( signal_5741 ), .Q ( signal_5742 ) ) ;
    buf_clk cell_3386 ( .C ( clk ), .D ( signal_5745 ), .Q ( signal_5746 ) ) ;
    buf_clk cell_3394 ( .C ( clk ), .D ( signal_5753 ), .Q ( signal_5754 ) ) ;
    buf_clk cell_3400 ( .C ( clk ), .D ( signal_5759 ), .Q ( signal_5760 ) ) ;
    buf_clk cell_3406 ( .C ( clk ), .D ( signal_5765 ), .Q ( signal_5766 ) ) ;
    buf_clk cell_3412 ( .C ( clk ), .D ( signal_5771 ), .Q ( signal_5772 ) ) ;
    buf_clk cell_3418 ( .C ( clk ), .D ( signal_5777 ), .Q ( signal_5778 ) ) ;
    buf_clk cell_3424 ( .C ( clk ), .D ( signal_5783 ), .Q ( signal_5784 ) ) ;
    buf_clk cell_3438 ( .C ( clk ), .D ( signal_5797 ), .Q ( signal_5798 ) ) ;
    buf_clk cell_3444 ( .C ( clk ), .D ( signal_5803 ), .Q ( signal_5804 ) ) ;
    buf_clk cell_3490 ( .C ( clk ), .D ( signal_5849 ), .Q ( signal_5850 ) ) ;
    buf_clk cell_3496 ( .C ( clk ), .D ( signal_5855 ), .Q ( signal_5856 ) ) ;
    buf_clk cell_3550 ( .C ( clk ), .D ( signal_5909 ), .Q ( signal_5910 ) ) ;
    buf_clk cell_3556 ( .C ( clk ), .D ( signal_5915 ), .Q ( signal_5916 ) ) ;
    buf_clk cell_3582 ( .C ( clk ), .D ( signal_5941 ), .Q ( signal_5942 ) ) ;
    buf_clk cell_3588 ( .C ( clk ), .D ( signal_5947 ), .Q ( signal_5948 ) ) ;
    buf_clk cell_3638 ( .C ( clk ), .D ( signal_5997 ), .Q ( signal_5998 ) ) ;
    buf_clk cell_3644 ( .C ( clk ), .D ( signal_6003 ), .Q ( signal_6004 ) ) ;
    buf_clk cell_3658 ( .C ( clk ), .D ( signal_6017 ), .Q ( signal_6018 ) ) ;
    buf_clk cell_3664 ( .C ( clk ), .D ( signal_6023 ), .Q ( signal_6024 ) ) ;
    buf_clk cell_3714 ( .C ( clk ), .D ( signal_6073 ), .Q ( signal_6074 ) ) ;
    buf_clk cell_3720 ( .C ( clk ), .D ( signal_6079 ), .Q ( signal_6080 ) ) ;
    buf_clk cell_3742 ( .C ( clk ), .D ( signal_6101 ), .Q ( signal_6102 ) ) ;
    buf_clk cell_3748 ( .C ( clk ), .D ( signal_6107 ), .Q ( signal_6108 ) ) ;
    buf_clk cell_3754 ( .C ( clk ), .D ( signal_6113 ), .Q ( signal_6114 ) ) ;
    buf_clk cell_3760 ( .C ( clk ), .D ( signal_6119 ), .Q ( signal_6120 ) ) ;
    buf_clk cell_3766 ( .C ( clk ), .D ( signal_6125 ), .Q ( signal_6126 ) ) ;
    buf_clk cell_3772 ( .C ( clk ), .D ( signal_6131 ), .Q ( signal_6132 ) ) ;
    buf_clk cell_3794 ( .C ( clk ), .D ( signal_6153 ), .Q ( signal_6154 ) ) ;
    buf_clk cell_3802 ( .C ( clk ), .D ( signal_6161 ), .Q ( signal_6162 ) ) ;
    buf_clk cell_3966 ( .C ( clk ), .D ( signal_6325 ), .Q ( signal_6326 ) ) ;
    buf_clk cell_3974 ( .C ( clk ), .D ( signal_6333 ), .Q ( signal_6334 ) ) ;
    buf_clk cell_4030 ( .C ( clk ), .D ( signal_6389 ), .Q ( signal_6390 ) ) ;
    buf_clk cell_4038 ( .C ( clk ), .D ( signal_6397 ), .Q ( signal_6398 ) ) ;
    buf_clk cell_4130 ( .C ( clk ), .D ( signal_6489 ), .Q ( signal_6490 ) ) ;
    buf_clk cell_4140 ( .C ( clk ), .D ( signal_6499 ), .Q ( signal_6500 ) ) ;
    buf_clk cell_4226 ( .C ( clk ), .D ( signal_6585 ), .Q ( signal_6586 ) ) ;
    buf_clk cell_4236 ( .C ( clk ), .D ( signal_6595 ), .Q ( signal_6596 ) ) ;
    buf_clk cell_4338 ( .C ( clk ), .D ( signal_6697 ), .Q ( signal_6698 ) ) ;
    buf_clk cell_4348 ( .C ( clk ), .D ( signal_6707 ), .Q ( signal_6708 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_3017 ( .C ( clk ), .D ( signal_1550 ), .Q ( signal_5377 ) ) ;
    buf_clk cell_3019 ( .C ( clk ), .D ( signal_3008 ), .Q ( signal_5379 ) ) ;
    buf_clk cell_3021 ( .C ( clk ), .D ( signal_1566 ), .Q ( signal_5381 ) ) ;
    buf_clk cell_3023 ( .C ( clk ), .D ( signal_3024 ), .Q ( signal_5383 ) ) ;
    buf_clk cell_3027 ( .C ( clk ), .D ( signal_5386 ), .Q ( signal_5387 ) ) ;
    buf_clk cell_3031 ( .C ( clk ), .D ( signal_5390 ), .Q ( signal_5391 ) ) ;
    buf_clk cell_3033 ( .C ( clk ), .D ( signal_1604 ), .Q ( signal_5393 ) ) ;
    buf_clk cell_3035 ( .C ( clk ), .D ( signal_3062 ), .Q ( signal_5395 ) ) ;
    buf_clk cell_3039 ( .C ( clk ), .D ( signal_5398 ), .Q ( signal_5399 ) ) ;
    buf_clk cell_3043 ( .C ( clk ), .D ( signal_5402 ), .Q ( signal_5403 ) ) ;
    buf_clk cell_3047 ( .C ( clk ), .D ( signal_5406 ), .Q ( signal_5407 ) ) ;
    buf_clk cell_3051 ( .C ( clk ), .D ( signal_5410 ), .Q ( signal_5411 ) ) ;
    buf_clk cell_3055 ( .C ( clk ), .D ( signal_5414 ), .Q ( signal_5415 ) ) ;
    buf_clk cell_3059 ( .C ( clk ), .D ( signal_5418 ), .Q ( signal_5419 ) ) ;
    buf_clk cell_3067 ( .C ( clk ), .D ( signal_5426 ), .Q ( signal_5427 ) ) ;
    buf_clk cell_3075 ( .C ( clk ), .D ( signal_5434 ), .Q ( signal_5435 ) ) ;
    buf_clk cell_3077 ( .C ( clk ), .D ( signal_1576 ), .Q ( signal_5437 ) ) ;
    buf_clk cell_3079 ( .C ( clk ), .D ( signal_3034 ), .Q ( signal_5439 ) ) ;
    buf_clk cell_3081 ( .C ( clk ), .D ( signal_1582 ), .Q ( signal_5441 ) ) ;
    buf_clk cell_3083 ( .C ( clk ), .D ( signal_3040 ), .Q ( signal_5443 ) ) ;
    buf_clk cell_3087 ( .C ( clk ), .D ( signal_5446 ), .Q ( signal_5447 ) ) ;
    buf_clk cell_3091 ( .C ( clk ), .D ( signal_5450 ), .Q ( signal_5451 ) ) ;
    buf_clk cell_3093 ( .C ( clk ), .D ( signal_1632 ), .Q ( signal_5453 ) ) ;
    buf_clk cell_3095 ( .C ( clk ), .D ( signal_3090 ), .Q ( signal_5455 ) ) ;
    buf_clk cell_3097 ( .C ( clk ), .D ( signal_1597 ), .Q ( signal_5457 ) ) ;
    buf_clk cell_3099 ( .C ( clk ), .D ( signal_3055 ), .Q ( signal_5459 ) ) ;
    buf_clk cell_3103 ( .C ( clk ), .D ( signal_5462 ), .Q ( signal_5463 ) ) ;
    buf_clk cell_3107 ( .C ( clk ), .D ( signal_5466 ), .Q ( signal_5467 ) ) ;
    buf_clk cell_3109 ( .C ( clk ), .D ( signal_1595 ), .Q ( signal_5469 ) ) ;
    buf_clk cell_3111 ( .C ( clk ), .D ( signal_3053 ), .Q ( signal_5471 ) ) ;
    buf_clk cell_3113 ( .C ( clk ), .D ( signal_1551 ), .Q ( signal_5473 ) ) ;
    buf_clk cell_3115 ( .C ( clk ), .D ( signal_3009 ), .Q ( signal_5475 ) ) ;
    buf_clk cell_3117 ( .C ( clk ), .D ( signal_1613 ), .Q ( signal_5477 ) ) ;
    buf_clk cell_3119 ( .C ( clk ), .D ( signal_3071 ), .Q ( signal_5479 ) ) ;
    buf_clk cell_3121 ( .C ( clk ), .D ( signal_1690 ), .Q ( signal_5481 ) ) ;
    buf_clk cell_3123 ( .C ( clk ), .D ( signal_3148 ), .Q ( signal_5483 ) ) ;
    buf_clk cell_3125 ( .C ( clk ), .D ( signal_1555 ), .Q ( signal_5485 ) ) ;
    buf_clk cell_3127 ( .C ( clk ), .D ( signal_3013 ), .Q ( signal_5487 ) ) ;
    buf_clk cell_3131 ( .C ( clk ), .D ( signal_5490 ), .Q ( signal_5491 ) ) ;
    buf_clk cell_3135 ( .C ( clk ), .D ( signal_5494 ), .Q ( signal_5495 ) ) ;
    buf_clk cell_3137 ( .C ( clk ), .D ( signal_1562 ), .Q ( signal_5497 ) ) ;
    buf_clk cell_3139 ( .C ( clk ), .D ( signal_3020 ), .Q ( signal_5499 ) ) ;
    buf_clk cell_3141 ( .C ( clk ), .D ( signal_1694 ), .Q ( signal_5501 ) ) ;
    buf_clk cell_3143 ( .C ( clk ), .D ( signal_3152 ), .Q ( signal_5503 ) ) ;
    buf_clk cell_3145 ( .C ( clk ), .D ( signal_1636 ), .Q ( signal_5505 ) ) ;
    buf_clk cell_3147 ( .C ( clk ), .D ( signal_3094 ), .Q ( signal_5507 ) ) ;
    buf_clk cell_3149 ( .C ( clk ), .D ( signal_1568 ), .Q ( signal_5509 ) ) ;
    buf_clk cell_3151 ( .C ( clk ), .D ( signal_3026 ), .Q ( signal_5511 ) ) ;
    buf_clk cell_3155 ( .C ( clk ), .D ( signal_5514 ), .Q ( signal_5515 ) ) ;
    buf_clk cell_3159 ( .C ( clk ), .D ( signal_5518 ), .Q ( signal_5519 ) ) ;
    buf_clk cell_3161 ( .C ( clk ), .D ( signal_1853 ), .Q ( signal_5521 ) ) ;
    buf_clk cell_3163 ( .C ( clk ), .D ( signal_3311 ), .Q ( signal_5523 ) ) ;
    buf_clk cell_3165 ( .C ( clk ), .D ( signal_5334 ), .Q ( signal_5525 ) ) ;
    buf_clk cell_3167 ( .C ( clk ), .D ( signal_5336 ), .Q ( signal_5527 ) ) ;
    buf_clk cell_3171 ( .C ( clk ), .D ( signal_5530 ), .Q ( signal_5531 ) ) ;
    buf_clk cell_3175 ( .C ( clk ), .D ( signal_5534 ), .Q ( signal_5535 ) ) ;
    buf_clk cell_3179 ( .C ( clk ), .D ( signal_5538 ), .Q ( signal_5539 ) ) ;
    buf_clk cell_3183 ( .C ( clk ), .D ( signal_5542 ), .Q ( signal_5543 ) ) ;
    buf_clk cell_3187 ( .C ( clk ), .D ( signal_5546 ), .Q ( signal_5547 ) ) ;
    buf_clk cell_3191 ( .C ( clk ), .D ( signal_5550 ), .Q ( signal_5551 ) ) ;
    buf_clk cell_3195 ( .C ( clk ), .D ( signal_5554 ), .Q ( signal_5555 ) ) ;
    buf_clk cell_3199 ( .C ( clk ), .D ( signal_5558 ), .Q ( signal_5559 ) ) ;
    buf_clk cell_3201 ( .C ( clk ), .D ( signal_5286 ), .Q ( signal_5561 ) ) ;
    buf_clk cell_3203 ( .C ( clk ), .D ( signal_5288 ), .Q ( signal_5563 ) ) ;
    buf_clk cell_3205 ( .C ( clk ), .D ( signal_5202 ), .Q ( signal_5565 ) ) ;
    buf_clk cell_3207 ( .C ( clk ), .D ( signal_5204 ), .Q ( signal_5567 ) ) ;
    buf_clk cell_3209 ( .C ( clk ), .D ( signal_1854 ), .Q ( signal_5569 ) ) ;
    buf_clk cell_3211 ( .C ( clk ), .D ( signal_3312 ), .Q ( signal_5571 ) ) ;
    buf_clk cell_3213 ( .C ( clk ), .D ( signal_5062 ), .Q ( signal_5573 ) ) ;
    buf_clk cell_3215 ( .C ( clk ), .D ( signal_5064 ), .Q ( signal_5575 ) ) ;
    buf_clk cell_3217 ( .C ( clk ), .D ( signal_5358 ), .Q ( signal_5577 ) ) ;
    buf_clk cell_3219 ( .C ( clk ), .D ( signal_5360 ), .Q ( signal_5579 ) ) ;
    buf_clk cell_3223 ( .C ( clk ), .D ( signal_5582 ), .Q ( signal_5583 ) ) ;
    buf_clk cell_3227 ( .C ( clk ), .D ( signal_5586 ), .Q ( signal_5587 ) ) ;
    buf_clk cell_3231 ( .C ( clk ), .D ( signal_5590 ), .Q ( signal_5591 ) ) ;
    buf_clk cell_3235 ( .C ( clk ), .D ( signal_5594 ), .Q ( signal_5595 ) ) ;
    buf_clk cell_3239 ( .C ( clk ), .D ( signal_5598 ), .Q ( signal_5599 ) ) ;
    buf_clk cell_3243 ( .C ( clk ), .D ( signal_5602 ), .Q ( signal_5603 ) ) ;
    buf_clk cell_3245 ( .C ( clk ), .D ( signal_1862 ), .Q ( signal_5605 ) ) ;
    buf_clk cell_3247 ( .C ( clk ), .D ( signal_3320 ), .Q ( signal_5607 ) ) ;
    buf_clk cell_3251 ( .C ( clk ), .D ( signal_5610 ), .Q ( signal_5611 ) ) ;
    buf_clk cell_3255 ( .C ( clk ), .D ( signal_5614 ), .Q ( signal_5615 ) ) ;
    buf_clk cell_3257 ( .C ( clk ), .D ( signal_5094 ), .Q ( signal_5617 ) ) ;
    buf_clk cell_3259 ( .C ( clk ), .D ( signal_5096 ), .Q ( signal_5619 ) ) ;
    buf_clk cell_3261 ( .C ( clk ), .D ( signal_1866 ), .Q ( signal_5621 ) ) ;
    buf_clk cell_3263 ( .C ( clk ), .D ( signal_3324 ), .Q ( signal_5623 ) ) ;
    buf_clk cell_3265 ( .C ( clk ), .D ( signal_5042 ), .Q ( signal_5625 ) ) ;
    buf_clk cell_3267 ( .C ( clk ), .D ( signal_5044 ), .Q ( signal_5627 ) ) ;
    buf_clk cell_3269 ( .C ( clk ), .D ( signal_1873 ), .Q ( signal_5629 ) ) ;
    buf_clk cell_3271 ( .C ( clk ), .D ( signal_3331 ), .Q ( signal_5631 ) ) ;
    buf_clk cell_3273 ( .C ( clk ), .D ( signal_1851 ), .Q ( signal_5633 ) ) ;
    buf_clk cell_3275 ( .C ( clk ), .D ( signal_3309 ), .Q ( signal_5635 ) ) ;
    buf_clk cell_3279 ( .C ( clk ), .D ( signal_5638 ), .Q ( signal_5639 ) ) ;
    buf_clk cell_3283 ( .C ( clk ), .D ( signal_5642 ), .Q ( signal_5643 ) ) ;
    buf_clk cell_3287 ( .C ( clk ), .D ( signal_5646 ), .Q ( signal_5647 ) ) ;
    buf_clk cell_3291 ( .C ( clk ), .D ( signal_5650 ), .Q ( signal_5651 ) ) ;
    buf_clk cell_3293 ( .C ( clk ), .D ( signal_1571 ), .Q ( signal_5653 ) ) ;
    buf_clk cell_3295 ( .C ( clk ), .D ( signal_3029 ), .Q ( signal_5655 ) ) ;
    buf_clk cell_3299 ( .C ( clk ), .D ( signal_5658 ), .Q ( signal_5659 ) ) ;
    buf_clk cell_3303 ( .C ( clk ), .D ( signal_5662 ), .Q ( signal_5663 ) ) ;
    buf_clk cell_3305 ( .C ( clk ), .D ( signal_1540 ), .Q ( signal_5665 ) ) ;
    buf_clk cell_3307 ( .C ( clk ), .D ( signal_2998 ), .Q ( signal_5667 ) ) ;
    buf_clk cell_3309 ( .C ( clk ), .D ( signal_1872 ), .Q ( signal_5669 ) ) ;
    buf_clk cell_3311 ( .C ( clk ), .D ( signal_3330 ), .Q ( signal_5671 ) ) ;
    buf_clk cell_3315 ( .C ( clk ), .D ( signal_5674 ), .Q ( signal_5675 ) ) ;
    buf_clk cell_3319 ( .C ( clk ), .D ( signal_5678 ), .Q ( signal_5679 ) ) ;
    buf_clk cell_3323 ( .C ( clk ), .D ( signal_5682 ), .Q ( signal_5683 ) ) ;
    buf_clk cell_3327 ( .C ( clk ), .D ( signal_5686 ), .Q ( signal_5687 ) ) ;
    buf_clk cell_3331 ( .C ( clk ), .D ( signal_5690 ), .Q ( signal_5691 ) ) ;
    buf_clk cell_3335 ( .C ( clk ), .D ( signal_5694 ), .Q ( signal_5695 ) ) ;
    buf_clk cell_3337 ( .C ( clk ), .D ( signal_1583 ), .Q ( signal_5697 ) ) ;
    buf_clk cell_3339 ( .C ( clk ), .D ( signal_3041 ), .Q ( signal_5699 ) ) ;
    buf_clk cell_3343 ( .C ( clk ), .D ( signal_5702 ), .Q ( signal_5703 ) ) ;
    buf_clk cell_3347 ( .C ( clk ), .D ( signal_5706 ), .Q ( signal_5707 ) ) ;
    buf_clk cell_3351 ( .C ( clk ), .D ( signal_5710 ), .Q ( signal_5711 ) ) ;
    buf_clk cell_3355 ( .C ( clk ), .D ( signal_5714 ), .Q ( signal_5715 ) ) ;
    buf_clk cell_3357 ( .C ( clk ), .D ( signal_1600 ), .Q ( signal_5717 ) ) ;
    buf_clk cell_3359 ( .C ( clk ), .D ( signal_3058 ), .Q ( signal_5719 ) ) ;
    buf_clk cell_3363 ( .C ( clk ), .D ( signal_5722 ), .Q ( signal_5723 ) ) ;
    buf_clk cell_3367 ( .C ( clk ), .D ( signal_5726 ), .Q ( signal_5727 ) ) ;
    buf_clk cell_3369 ( .C ( clk ), .D ( signal_1870 ), .Q ( signal_5729 ) ) ;
    buf_clk cell_3371 ( .C ( clk ), .D ( signal_3328 ), .Q ( signal_5731 ) ) ;
    buf_clk cell_3373 ( .C ( clk ), .D ( signal_1312 ), .Q ( signal_5733 ) ) ;
    buf_clk cell_3375 ( .C ( clk ), .D ( signal_2770 ), .Q ( signal_5735 ) ) ;
    buf_clk cell_3377 ( .C ( clk ), .D ( signal_5078 ), .Q ( signal_5737 ) ) ;
    buf_clk cell_3379 ( .C ( clk ), .D ( signal_5080 ), .Q ( signal_5739 ) ) ;
    buf_clk cell_3383 ( .C ( clk ), .D ( signal_5742 ), .Q ( signal_5743 ) ) ;
    buf_clk cell_3387 ( .C ( clk ), .D ( signal_5746 ), .Q ( signal_5747 ) ) ;
    buf_clk cell_3395 ( .C ( clk ), .D ( signal_5754 ), .Q ( signal_5755 ) ) ;
    buf_clk cell_3401 ( .C ( clk ), .D ( signal_5760 ), .Q ( signal_5761 ) ) ;
    buf_clk cell_3407 ( .C ( clk ), .D ( signal_5766 ), .Q ( signal_5767 ) ) ;
    buf_clk cell_3413 ( .C ( clk ), .D ( signal_5772 ), .Q ( signal_5773 ) ) ;
    buf_clk cell_3419 ( .C ( clk ), .D ( signal_5778 ), .Q ( signal_5779 ) ) ;
    buf_clk cell_3425 ( .C ( clk ), .D ( signal_5784 ), .Q ( signal_5785 ) ) ;
    buf_clk cell_3429 ( .C ( clk ), .D ( signal_1537 ), .Q ( signal_5789 ) ) ;
    buf_clk cell_3433 ( .C ( clk ), .D ( signal_2995 ), .Q ( signal_5793 ) ) ;
    buf_clk cell_3439 ( .C ( clk ), .D ( signal_5798 ), .Q ( signal_5799 ) ) ;
    buf_clk cell_3445 ( .C ( clk ), .D ( signal_5804 ), .Q ( signal_5805 ) ) ;
    buf_clk cell_3449 ( .C ( clk ), .D ( signal_1552 ), .Q ( signal_5809 ) ) ;
    buf_clk cell_3453 ( .C ( clk ), .D ( signal_3010 ), .Q ( signal_5813 ) ) ;
    buf_clk cell_3457 ( .C ( clk ), .D ( signal_1618 ), .Q ( signal_5817 ) ) ;
    buf_clk cell_3461 ( .C ( clk ), .D ( signal_3076 ), .Q ( signal_5821 ) ) ;
    buf_clk cell_3465 ( .C ( clk ), .D ( signal_1560 ), .Q ( signal_5825 ) ) ;
    buf_clk cell_3469 ( .C ( clk ), .D ( signal_3018 ), .Q ( signal_5829 ) ) ;
    buf_clk cell_3473 ( .C ( clk ), .D ( signal_1622 ), .Q ( signal_5833 ) ) ;
    buf_clk cell_3477 ( .C ( clk ), .D ( signal_3080 ), .Q ( signal_5837 ) ) ;
    buf_clk cell_3481 ( .C ( clk ), .D ( signal_1533 ), .Q ( signal_5841 ) ) ;
    buf_clk cell_3485 ( .C ( clk ), .D ( signal_2991 ), .Q ( signal_5845 ) ) ;
    buf_clk cell_3491 ( .C ( clk ), .D ( signal_5850 ), .Q ( signal_5851 ) ) ;
    buf_clk cell_3497 ( .C ( clk ), .D ( signal_5856 ), .Q ( signal_5857 ) ) ;
    buf_clk cell_3501 ( .C ( clk ), .D ( signal_5106 ), .Q ( signal_5861 ) ) ;
    buf_clk cell_3505 ( .C ( clk ), .D ( signal_5108 ), .Q ( signal_5865 ) ) ;
    buf_clk cell_3529 ( .C ( clk ), .D ( signal_1591 ), .Q ( signal_5889 ) ) ;
    buf_clk cell_3533 ( .C ( clk ), .D ( signal_3049 ), .Q ( signal_5893 ) ) ;
    buf_clk cell_3551 ( .C ( clk ), .D ( signal_5910 ), .Q ( signal_5911 ) ) ;
    buf_clk cell_3557 ( .C ( clk ), .D ( signal_5916 ), .Q ( signal_5917 ) ) ;
    buf_clk cell_3565 ( .C ( clk ), .D ( signal_1621 ), .Q ( signal_5925 ) ) ;
    buf_clk cell_3569 ( .C ( clk ), .D ( signal_3079 ), .Q ( signal_5929 ) ) ;
    buf_clk cell_3583 ( .C ( clk ), .D ( signal_5942 ), .Q ( signal_5943 ) ) ;
    buf_clk cell_3589 ( .C ( clk ), .D ( signal_5948 ), .Q ( signal_5949 ) ) ;
    buf_clk cell_3593 ( .C ( clk ), .D ( signal_5362 ), .Q ( signal_5953 ) ) ;
    buf_clk cell_3597 ( .C ( clk ), .D ( signal_5364 ), .Q ( signal_5957 ) ) ;
    buf_clk cell_3609 ( .C ( clk ), .D ( signal_1606 ), .Q ( signal_5969 ) ) ;
    buf_clk cell_3613 ( .C ( clk ), .D ( signal_3064 ), .Q ( signal_5973 ) ) ;
    buf_clk cell_3617 ( .C ( clk ), .D ( signal_1691 ), .Q ( signal_5977 ) ) ;
    buf_clk cell_3621 ( .C ( clk ), .D ( signal_3149 ), .Q ( signal_5981 ) ) ;
    buf_clk cell_3625 ( .C ( clk ), .D ( signal_1570 ), .Q ( signal_5985 ) ) ;
    buf_clk cell_3629 ( .C ( clk ), .D ( signal_3028 ), .Q ( signal_5989 ) ) ;
    buf_clk cell_3639 ( .C ( clk ), .D ( signal_5998 ), .Q ( signal_5999 ) ) ;
    buf_clk cell_3645 ( .C ( clk ), .D ( signal_6004 ), .Q ( signal_6005 ) ) ;
    buf_clk cell_3649 ( .C ( clk ), .D ( signal_1584 ), .Q ( signal_6009 ) ) ;
    buf_clk cell_3653 ( .C ( clk ), .D ( signal_3042 ), .Q ( signal_6013 ) ) ;
    buf_clk cell_3659 ( .C ( clk ), .D ( signal_6018 ), .Q ( signal_6019 ) ) ;
    buf_clk cell_3665 ( .C ( clk ), .D ( signal_6024 ), .Q ( signal_6025 ) ) ;
    buf_clk cell_3669 ( .C ( clk ), .D ( signal_1590 ), .Q ( signal_6029 ) ) ;
    buf_clk cell_3673 ( .C ( clk ), .D ( signal_3048 ), .Q ( signal_6033 ) ) ;
    buf_clk cell_3677 ( .C ( clk ), .D ( signal_1675 ), .Q ( signal_6037 ) ) ;
    buf_clk cell_3681 ( .C ( clk ), .D ( signal_3133 ), .Q ( signal_6041 ) ) ;
    buf_clk cell_3685 ( .C ( clk ), .D ( signal_1598 ), .Q ( signal_6045 ) ) ;
    buf_clk cell_3689 ( .C ( clk ), .D ( signal_3056 ), .Q ( signal_6049 ) ) ;
    buf_clk cell_3697 ( .C ( clk ), .D ( signal_1601 ), .Q ( signal_6057 ) ) ;
    buf_clk cell_3701 ( .C ( clk ), .D ( signal_3059 ), .Q ( signal_6061 ) ) ;
    buf_clk cell_3705 ( .C ( clk ), .D ( signal_1543 ), .Q ( signal_6065 ) ) ;
    buf_clk cell_3709 ( .C ( clk ), .D ( signal_3001 ), .Q ( signal_6069 ) ) ;
    buf_clk cell_3715 ( .C ( clk ), .D ( signal_6074 ), .Q ( signal_6075 ) ) ;
    buf_clk cell_3721 ( .C ( clk ), .D ( signal_6080 ), .Q ( signal_6081 ) ) ;
    buf_clk cell_3733 ( .C ( clk ), .D ( signal_1625 ), .Q ( signal_6093 ) ) ;
    buf_clk cell_3737 ( .C ( clk ), .D ( signal_3083 ), .Q ( signal_6097 ) ) ;
    buf_clk cell_3743 ( .C ( clk ), .D ( signal_6102 ), .Q ( signal_6103 ) ) ;
    buf_clk cell_3749 ( .C ( clk ), .D ( signal_6108 ), .Q ( signal_6109 ) ) ;
    buf_clk cell_3755 ( .C ( clk ), .D ( signal_6114 ), .Q ( signal_6115 ) ) ;
    buf_clk cell_3761 ( .C ( clk ), .D ( signal_6120 ), .Q ( signal_6121 ) ) ;
    buf_clk cell_3767 ( .C ( clk ), .D ( signal_6126 ), .Q ( signal_6127 ) ) ;
    buf_clk cell_3773 ( .C ( clk ), .D ( signal_6132 ), .Q ( signal_6133 ) ) ;
    buf_clk cell_3777 ( .C ( clk ), .D ( signal_5278 ), .Q ( signal_6137 ) ) ;
    buf_clk cell_3781 ( .C ( clk ), .D ( signal_5284 ), .Q ( signal_6141 ) ) ;
    buf_clk cell_3795 ( .C ( clk ), .D ( signal_6154 ), .Q ( signal_6155 ) ) ;
    buf_clk cell_3803 ( .C ( clk ), .D ( signal_6162 ), .Q ( signal_6163 ) ) ;
    buf_clk cell_3817 ( .C ( clk ), .D ( signal_1645 ), .Q ( signal_6177 ) ) ;
    buf_clk cell_3823 ( .C ( clk ), .D ( signal_3103 ), .Q ( signal_6183 ) ) ;
    buf_clk cell_3829 ( .C ( clk ), .D ( signal_1616 ), .Q ( signal_6189 ) ) ;
    buf_clk cell_3835 ( .C ( clk ), .D ( signal_3074 ), .Q ( signal_6195 ) ) ;
    buf_clk cell_3849 ( .C ( clk ), .D ( signal_1534 ), .Q ( signal_6209 ) ) ;
    buf_clk cell_3855 ( .C ( clk ), .D ( signal_2992 ), .Q ( signal_6215 ) ) ;
    buf_clk cell_3885 ( .C ( clk ), .D ( signal_1850 ), .Q ( signal_6245 ) ) ;
    buf_clk cell_3891 ( .C ( clk ), .D ( signal_3308 ), .Q ( signal_6251 ) ) ;
    buf_clk cell_3897 ( .C ( clk ), .D ( signal_1631 ), .Q ( signal_6257 ) ) ;
    buf_clk cell_3903 ( .C ( clk ), .D ( signal_3089 ), .Q ( signal_6263 ) ) ;
    buf_clk cell_3909 ( .C ( clk ), .D ( signal_1683 ), .Q ( signal_6269 ) ) ;
    buf_clk cell_3915 ( .C ( clk ), .D ( signal_3141 ), .Q ( signal_6275 ) ) ;
    buf_clk cell_3933 ( .C ( clk ), .D ( signal_1299 ), .Q ( signal_6293 ) ) ;
    buf_clk cell_3939 ( .C ( clk ), .D ( signal_2757 ), .Q ( signal_6299 ) ) ;
    buf_clk cell_3949 ( .C ( clk ), .D ( signal_1557 ), .Q ( signal_6309 ) ) ;
    buf_clk cell_3955 ( .C ( clk ), .D ( signal_3015 ), .Q ( signal_6315 ) ) ;
    buf_clk cell_3967 ( .C ( clk ), .D ( signal_6326 ), .Q ( signal_6327 ) ) ;
    buf_clk cell_3975 ( .C ( clk ), .D ( signal_6334 ), .Q ( signal_6335 ) ) ;
    buf_clk cell_3997 ( .C ( clk ), .D ( signal_1506 ), .Q ( signal_6357 ) ) ;
    buf_clk cell_4003 ( .C ( clk ), .D ( signal_2964 ), .Q ( signal_6363 ) ) ;
    buf_clk cell_4009 ( .C ( clk ), .D ( signal_1593 ), .Q ( signal_6369 ) ) ;
    buf_clk cell_4015 ( .C ( clk ), .D ( signal_3051 ), .Q ( signal_6375 ) ) ;
    buf_clk cell_4031 ( .C ( clk ), .D ( signal_6390 ), .Q ( signal_6391 ) ) ;
    buf_clk cell_4039 ( .C ( clk ), .D ( signal_6398 ), .Q ( signal_6399 ) ) ;
    buf_clk cell_4045 ( .C ( clk ), .D ( signal_1338 ), .Q ( signal_6405 ) ) ;
    buf_clk cell_4051 ( .C ( clk ), .D ( signal_2796 ), .Q ( signal_6411 ) ) ;
    buf_clk cell_4057 ( .C ( clk ), .D ( signal_5070 ), .Q ( signal_6417 ) ) ;
    buf_clk cell_4063 ( .C ( clk ), .D ( signal_5072 ), .Q ( signal_6423 ) ) ;
    buf_clk cell_4077 ( .C ( clk ), .D ( signal_5250 ), .Q ( signal_6437 ) ) ;
    buf_clk cell_4083 ( .C ( clk ), .D ( signal_5252 ), .Q ( signal_6443 ) ) ;
    buf_clk cell_4097 ( .C ( clk ), .D ( signal_1637 ), .Q ( signal_6457 ) ) ;
    buf_clk cell_4103 ( .C ( clk ), .D ( signal_3095 ), .Q ( signal_6463 ) ) ;
    buf_clk cell_4109 ( .C ( clk ), .D ( signal_1518 ), .Q ( signal_6469 ) ) ;
    buf_clk cell_4115 ( .C ( clk ), .D ( signal_2976 ), .Q ( signal_6475 ) ) ;
    buf_clk cell_4131 ( .C ( clk ), .D ( signal_6490 ), .Q ( signal_6491 ) ) ;
    buf_clk cell_4141 ( .C ( clk ), .D ( signal_6500 ), .Q ( signal_6501 ) ) ;
    buf_clk cell_4161 ( .C ( clk ), .D ( signal_1619 ), .Q ( signal_6521 ) ) ;
    buf_clk cell_4169 ( .C ( clk ), .D ( signal_3077 ), .Q ( signal_6529 ) ) ;
    buf_clk cell_4177 ( .C ( clk ), .D ( signal_1350 ), .Q ( signal_6537 ) ) ;
    buf_clk cell_4185 ( .C ( clk ), .D ( signal_2808 ), .Q ( signal_6545 ) ) ;
    buf_clk cell_4227 ( .C ( clk ), .D ( signal_6586 ), .Q ( signal_6587 ) ) ;
    buf_clk cell_4237 ( .C ( clk ), .D ( signal_6596 ), .Q ( signal_6597 ) ) ;
    buf_clk cell_4261 ( .C ( clk ), .D ( signal_1575 ), .Q ( signal_6621 ) ) ;
    buf_clk cell_4269 ( .C ( clk ), .D ( signal_3033 ), .Q ( signal_6629 ) ) ;
    buf_clk cell_4289 ( .C ( clk ), .D ( signal_1587 ), .Q ( signal_6649 ) ) ;
    buf_clk cell_4297 ( .C ( clk ), .D ( signal_3045 ), .Q ( signal_6657 ) ) ;
    buf_clk cell_4305 ( .C ( clk ), .D ( signal_1861 ), .Q ( signal_6665 ) ) ;
    buf_clk cell_4313 ( .C ( clk ), .D ( signal_3319 ), .Q ( signal_6673 ) ) ;
    buf_clk cell_4321 ( .C ( clk ), .D ( signal_1258 ), .Q ( signal_6681 ) ) ;
    buf_clk cell_4329 ( .C ( clk ), .D ( signal_2716 ), .Q ( signal_6689 ) ) ;
    buf_clk cell_4339 ( .C ( clk ), .D ( signal_6698 ), .Q ( signal_6699 ) ) ;
    buf_clk cell_4349 ( .C ( clk ), .D ( signal_6708 ), .Q ( signal_6709 ) ) ;
    buf_clk cell_4357 ( .C ( clk ), .D ( signal_5102 ), .Q ( signal_6717 ) ) ;
    buf_clk cell_4365 ( .C ( clk ), .D ( signal_5104 ), .Q ( signal_6725 ) ) ;
    buf_clk cell_4373 ( .C ( clk ), .D ( signal_1614 ), .Q ( signal_6733 ) ) ;
    buf_clk cell_4381 ( .C ( clk ), .D ( signal_3072 ), .Q ( signal_6741 ) ) ;
    buf_clk cell_4393 ( .C ( clk ), .D ( signal_1549 ), .Q ( signal_6753 ) ) ;
    buf_clk cell_4401 ( .C ( clk ), .D ( signal_3007 ), .Q ( signal_6761 ) ) ;
    buf_clk cell_4409 ( .C ( clk ), .D ( signal_1578 ), .Q ( signal_6769 ) ) ;
    buf_clk cell_4417 ( .C ( clk ), .D ( signal_3036 ), .Q ( signal_6777 ) ) ;
    buf_clk cell_4425 ( .C ( clk ), .D ( signal_1581 ), .Q ( signal_6785 ) ) ;
    buf_clk cell_4433 ( .C ( clk ), .D ( signal_3039 ), .Q ( signal_6793 ) ) ;
    buf_clk cell_4509 ( .C ( clk ), .D ( signal_1505 ), .Q ( signal_6869 ) ) ;
    buf_clk cell_4519 ( .C ( clk ), .D ( signal_2963 ), .Q ( signal_6879 ) ) ;
    buf_clk cell_4561 ( .C ( clk ), .D ( signal_1589 ), .Q ( signal_6921 ) ) ;
    buf_clk cell_4571 ( .C ( clk ), .D ( signal_3047 ), .Q ( signal_6931 ) ) ;
    buf_clk cell_4965 ( .C ( clk ), .D ( signal_1527 ), .Q ( signal_7325 ) ) ;
    buf_clk cell_4979 ( .C ( clk ), .D ( signal_2985 ), .Q ( signal_7339 ) ) ;
    buf_clk cell_5009 ( .C ( clk ), .D ( signal_1633 ), .Q ( signal_7369 ) ) ;
    buf_clk cell_5023 ( .C ( clk ), .D ( signal_3091 ), .Q ( signal_7383 ) ) ;
    buf_clk cell_5089 ( .C ( clk ), .D ( signal_1588 ), .Q ( signal_7449 ) ) ;
    buf_clk cell_5105 ( .C ( clk ), .D ( signal_3046 ), .Q ( signal_7465 ) ) ;
    buf_clk cell_5129 ( .C ( clk ), .D ( signal_1602 ), .Q ( signal_7489 ) ) ;
    buf_clk cell_5145 ( .C ( clk ), .D ( signal_3060 ), .Q ( signal_7505 ) ) ;
    buf_clk cell_5285 ( .C ( clk ), .D ( signal_1539 ), .Q ( signal_7645 ) ) ;
    buf_clk cell_5303 ( .C ( clk ), .D ( signal_2997 ), .Q ( signal_7663 ) ) ;
    buf_clk cell_5385 ( .C ( clk ), .D ( signal_1603 ), .Q ( signal_7745 ) ) ;
    buf_clk cell_5405 ( .C ( clk ), .D ( signal_3061 ), .Q ( signal_7765 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1644 ( .a ({signal_2750, signal_1292}), .b ({signal_5040, signal_5038}), .clk ( clk ), .r ( Fresh[454] ), .c ({signal_3117, signal_1659}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1652 ( .a ({signal_5044, signal_5042}), .b ({signal_2843, signal_1385}), .clk ( clk ), .r ( Fresh[455] ), .c ({signal_3125, signal_1667}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1662 ( .a ({signal_5048, signal_5046}), .b ({signal_2787, signal_1329}), .clk ( clk ), .r ( Fresh[456] ), .c ({signal_3135, signal_1677}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1672 ( .a ({signal_5052, signal_5050}), .b ({signal_2801, signal_1343}), .clk ( clk ), .r ( Fresh[457] ), .c ({signal_3145, signal_1687}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1683 ( .a ({signal_5056, signal_5054}), .b ({signal_2816, signal_1358}), .clk ( clk ), .r ( Fresh[458] ), .c ({signal_3156, signal_1698}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1685 ( .a ({signal_5060, signal_5058}), .b ({signal_2818, signal_1360}), .clk ( clk ), .r ( Fresh[459] ), .c ({signal_3158, signal_1700}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1686 ( .a ({signal_5064, signal_5062}), .b ({signal_2904, signal_1446}), .clk ( clk ), .r ( Fresh[460] ), .c ({signal_3159, signal_1701}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1688 ( .a ({signal_5068, signal_5066}), .b ({signal_2904, signal_1446}), .clk ( clk ), .r ( Fresh[461] ), .c ({signal_3161, signal_1703}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1689 ( .a ({signal_5068, signal_5066}), .b ({signal_2918, signal_1460}), .clk ( clk ), .r ( Fresh[462] ), .c ({signal_3162, signal_1704}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1690 ( .a ({signal_5072, signal_5070}), .b ({signal_2919, signal_1461}), .clk ( clk ), .r ( Fresh[463] ), .c ({signal_3163, signal_1705}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1691 ( .a ({signal_5076, signal_5074}), .b ({signal_2920, signal_1462}), .clk ( clk ), .r ( Fresh[464] ), .c ({signal_3164, signal_1706}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1692 ( .a ({signal_5080, signal_5078}), .b ({signal_2908, signal_1450}), .clk ( clk ), .r ( Fresh[465] ), .c ({signal_3165, signal_1707}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1694 ( .a ({signal_5092, signal_5086}), .b ({signal_2936, signal_1478}), .clk ( clk ), .r ( Fresh[466] ), .c ({signal_3167, signal_1709}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1695 ( .a ({signal_5096, signal_5094}), .b ({signal_2821, signal_1363}), .clk ( clk ), .r ( Fresh[467] ), .c ({signal_3168, signal_1710}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1696 ( .a ({signal_5100, signal_5098}), .b ({signal_2893, signal_1435}), .clk ( clk ), .r ( Fresh[468] ), .c ({signal_3169, signal_1711}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1697 ( .a ({signal_5104, signal_5102}), .b ({signal_2932, signal_1474}), .clk ( clk ), .r ( Fresh[469] ), .c ({signal_3170, signal_1712}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1699 ( .a ({signal_5108, signal_5106}), .b ({signal_2955, signal_1497}), .clk ( clk ), .r ( Fresh[470] ), .c ({signal_3172, signal_1714}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1715 ( .a ({signal_3117, signal_1659}), .b ({signal_3188, signal_1730}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1721 ( .a ({signal_3125, signal_1667}), .b ({signal_3194, signal_1736}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1725 ( .a ({signal_3135, signal_1677}), .b ({signal_3198, signal_1740}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1737 ( .a ({signal_3158, signal_1700}), .b ({signal_3210, signal_1752}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1738 ( .a ({signal_3159, signal_1701}), .b ({signal_3211, signal_1753}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1740 ( .a ({signal_3161, signal_1703}), .b ({signal_3213, signal_1755}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1741 ( .a ({signal_3162, signal_1704}), .b ({signal_3214, signal_1756}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1742 ( .a ({signal_3163, signal_1705}), .b ({signal_3215, signal_1757}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1743 ( .a ({signal_3164, signal_1706}), .b ({signal_3216, signal_1758}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1744 ( .a ({signal_3165, signal_1707}), .b ({signal_3217, signal_1759}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1746 ( .a ({signal_3167, signal_1709}), .b ({signal_3219, signal_1761}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1747 ( .a ({signal_3169, signal_1711}), .b ({signal_3220, signal_1762}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1748 ( .a ({signal_3170, signal_1712}), .b ({signal_3221, signal_1763}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1750 ( .a ({signal_3172, signal_1714}), .b ({signal_3223, signal_1765}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1752 ( .a ({signal_2989, signal_1531}), .b ({signal_2990, signal_1532}), .clk ( clk ), .r ( Fresh[471] ), .c ({signal_3225, signal_1767}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1759 ( .a ({signal_5112, signal_5110}), .b ({signal_2970, signal_1512}), .clk ( clk ), .r ( Fresh[472] ), .c ({signal_3232, signal_1774}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1763 ( .a ({signal_5116, signal_5114}), .b ({signal_2975, signal_1517}), .clk ( clk ), .r ( Fresh[473] ), .c ({signal_3236, signal_1778}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1768 ( .a ({signal_2983, signal_1525}), .b ({signal_2984, signal_1526}), .clk ( clk ), .r ( Fresh[474] ), .c ({signal_3241, signal_1783}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1771 ( .a ({signal_2981, signal_1523}), .b ({signal_2988, signal_1530}), .clk ( clk ), .r ( Fresh[475] ), .c ({signal_3244, signal_1786}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1774 ( .a ({signal_5120, signal_5118}), .b ({signal_2994, signal_1536}), .clk ( clk ), .r ( Fresh[476] ), .c ({signal_3247, signal_1789}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1775 ( .a ({signal_2999, signal_1541}), .b ({signal_3000, signal_1542}), .clk ( clk ), .r ( Fresh[477] ), .c ({signal_3248, signal_1790}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1777 ( .a ({signal_5124, signal_5122}), .b ({signal_3004, signal_1546}), .clk ( clk ), .r ( Fresh[478] ), .c ({signal_3250, signal_1792}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1780 ( .a ({signal_5128, signal_5126}), .b ({signal_3107, signal_1649}), .clk ( clk ), .r ( Fresh[479] ), .c ({signal_3253, signal_1795}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1781 ( .a ({signal_3052, signal_1594}), .b ({signal_3069, signal_1611}), .clk ( clk ), .r ( Fresh[480] ), .c ({signal_3254, signal_1796}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1787 ( .a ({signal_5132, signal_5130}), .b ({signal_3019, signal_1561}), .clk ( clk ), .r ( Fresh[481] ), .c ({signal_3260, signal_1802}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1788 ( .a ({signal_3021, signal_1563}), .b ({signal_5136, signal_5134}), .clk ( clk ), .r ( Fresh[482] ), .c ({signal_3261, signal_1803}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1789 ( .a ({signal_5140, signal_5138}), .b ({signal_3111, signal_1653}), .clk ( clk ), .r ( Fresh[483] ), .c ({signal_3262, signal_1804}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1790 ( .a ({signal_5144, signal_5142}), .b ({signal_3112, signal_1654}), .clk ( clk ), .r ( Fresh[484] ), .c ({signal_3263, signal_1805}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1791 ( .a ({signal_5148, signal_5146}), .b ({signal_3113, signal_1655}), .clk ( clk ), .r ( Fresh[485] ), .c ({signal_3264, signal_1806}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1792 ( .a ({signal_3024, signal_1566}), .b ({signal_3025, signal_1567}), .clk ( clk ), .r ( Fresh[486] ), .c ({signal_3265, signal_1807}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1793 ( .a ({signal_2745, signal_1287}), .b ({signal_3026, signal_1568}), .clk ( clk ), .r ( Fresh[487] ), .c ({signal_3266, signal_1808}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1794 ( .a ({signal_3098, signal_1640}), .b ({signal_3027, signal_1569}), .clk ( clk ), .r ( Fresh[488] ), .c ({signal_3267, signal_1809}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1795 ( .a ({signal_5072, signal_5070}), .b ({signal_3029, signal_1571}), .clk ( clk ), .r ( Fresh[489] ), .c ({signal_3268, signal_1810}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1796 ( .a ({signal_2971, signal_1513}), .b ({signal_3030, signal_1572}), .clk ( clk ), .r ( Fresh[490] ), .c ({signal_3269, signal_1811}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1797 ( .a ({signal_5152, signal_5150}), .b ({signal_3031, signal_1573}), .clk ( clk ), .r ( Fresh[491] ), .c ({signal_3270, signal_1812}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1798 ( .a ({signal_5156, signal_5154}), .b ({signal_3118, signal_1660}), .clk ( clk ), .r ( Fresh[492] ), .c ({signal_3271, signal_1813}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1799 ( .a ({signal_5160, signal_5158}), .b ({signal_3032, signal_1574}), .clk ( clk ), .r ( Fresh[493] ), .c ({signal_3272, signal_1814}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1800 ( .a ({signal_5164, signal_5162}), .b ({signal_3035, signal_1577}), .clk ( clk ), .r ( Fresh[494] ), .c ({signal_3273, signal_1815}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1801 ( .a ({signal_5168, signal_5166}), .b ({signal_3119, signal_1661}), .clk ( clk ), .r ( Fresh[495] ), .c ({signal_3274, signal_1816}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1802 ( .a ({signal_5172, signal_5170}), .b ({signal_3024, signal_1566}), .clk ( clk ), .r ( Fresh[496] ), .c ({signal_3275, signal_1817}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1803 ( .a ({signal_3037, signal_1579}), .b ({signal_3038, signal_1580}), .clk ( clk ), .r ( Fresh[497] ), .c ({signal_3276, signal_1818}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1804 ( .a ({signal_2982, signal_1524}), .b ({signal_3043, signal_1585}), .clk ( clk ), .r ( Fresh[498] ), .c ({signal_3277, signal_1819}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1805 ( .a ({signal_3032, signal_1574}), .b ({signal_3044, signal_1586}), .clk ( clk ), .r ( Fresh[499] ), .c ({signal_3278, signal_1820}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1806 ( .a ({signal_5180, signal_5176}), .b ({signal_3126, signal_1668}), .clk ( clk ), .r ( Fresh[500] ), .c ({signal_3279, signal_1821}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1807 ( .a ({signal_5184, signal_5182}), .b ({signal_3124, signal_1666}), .clk ( clk ), .r ( Fresh[501] ), .c ({signal_3280, signal_1822}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1808 ( .a ({signal_5188, signal_5186}), .b ({signal_3128, signal_1670}), .clk ( clk ), .r ( Fresh[502] ), .c ({signal_3281, signal_1823}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1809 ( .a ({signal_5196, signal_5192}), .b ({signal_3129, signal_1671}), .clk ( clk ), .r ( Fresh[503] ), .c ({signal_3282, signal_1824}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1810 ( .a ({signal_3087, signal_1629}), .b ({signal_3088, signal_1630}), .clk ( clk ), .r ( Fresh[504] ), .c ({signal_3283, signal_1825}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1811 ( .a ({signal_2987, signal_1529}), .b ({signal_3130, signal_1672}), .clk ( clk ), .r ( Fresh[505] ), .c ({signal_3284, signal_1826}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1812 ( .a ({signal_2996, signal_1538}), .b ({signal_3057, signal_1599}), .clk ( clk ), .r ( Fresh[506] ), .c ({signal_3285, signal_1827}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1813 ( .a ({signal_3002, signal_1544}), .b ({signal_3063, signal_1605}), .clk ( clk ), .r ( Fresh[507] ), .c ({signal_3286, signal_1828}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1814 ( .a ({signal_3003, signal_1545}), .b ({signal_3065, signal_1607}), .clk ( clk ), .r ( Fresh[508] ), .c ({signal_3287, signal_1829}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1815 ( .a ({signal_5200, signal_5198}), .b ({signal_3066, signal_1608}), .clk ( clk ), .r ( Fresh[509] ), .c ({signal_3288, signal_1830}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1816 ( .a ({signal_5204, signal_5202}), .b ({signal_3142, signal_1684}), .clk ( clk ), .r ( Fresh[510] ), .c ({signal_3289, signal_1831}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1817 ( .a ({signal_5208, signal_5206}), .b ({signal_3143, signal_1685}), .clk ( clk ), .r ( Fresh[511] ), .c ({signal_3290, signal_1832}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1818 ( .a ({signal_3029, signal_1571}), .b ({signal_3054, signal_1596}), .clk ( clk ), .r ( Fresh[512] ), .c ({signal_3291, signal_1833}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1820 ( .a ({signal_2802, signal_1344}), .b ({signal_3068, signal_1610}), .clk ( clk ), .r ( Fresh[513] ), .c ({signal_3293, signal_1835}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1821 ( .a ({signal_5212, signal_5210}), .b ({signal_3070, signal_1612}), .clk ( clk ), .r ( Fresh[514] ), .c ({signal_3294, signal_1836}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1822 ( .a ({signal_5216, signal_5214}), .b ({signal_3073, signal_1615}), .clk ( clk ), .r ( Fresh[515] ), .c ({signal_3295, signal_1837}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1823 ( .a ({signal_3014, signal_1556}), .b ({signal_3075, signal_1617}), .clk ( clk ), .r ( Fresh[516] ), .c ({signal_3296, signal_1838}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1824 ( .a ({signal_5220, signal_5218}), .b ({signal_3150, signal_1692}), .clk ( clk ), .r ( Fresh[517] ), .c ({signal_3297, signal_1839}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1825 ( .a ({signal_5224, signal_5222}), .b ({signal_3078, signal_1620}), .clk ( clk ), .r ( Fresh[518] ), .c ({signal_3298, signal_1840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1826 ( .a ({signal_5228, signal_5226}), .b ({signal_3073, signal_1615}), .clk ( clk ), .r ( Fresh[519] ), .c ({signal_3299, signal_1841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1827 ( .a ({signal_5232, signal_5230}), .b ({signal_3153, signal_1695}), .clk ( clk ), .r ( Fresh[520] ), .c ({signal_3300, signal_1842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1828 ( .a ({signal_3022, signal_1564}), .b ({signal_3081, signal_1623}), .clk ( clk ), .r ( Fresh[521] ), .c ({signal_3301, signal_1843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1829 ( .a ({signal_5236, signal_5234}), .b ({signal_3082, signal_1624}), .clk ( clk ), .r ( Fresh[522] ), .c ({signal_3302, signal_1844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1830 ( .a ({signal_3084, signal_1626}), .b ({signal_3085, signal_1627}), .clk ( clk ), .r ( Fresh[523] ), .c ({signal_3303, signal_1845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1831 ( .a ({signal_3050, signal_1592}), .b ({signal_3086, signal_1628}), .clk ( clk ), .r ( Fresh[524] ), .c ({signal_3304, signal_1846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1832 ( .a ({signal_2981, signal_1523}), .b ({signal_3092, signal_1634}), .clk ( clk ), .r ( Fresh[525] ), .c ({signal_3305, signal_1847}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1833 ( .a ({signal_2820, signal_1362}), .b ({signal_3093, signal_1635}), .clk ( clk ), .r ( Fresh[526] ), .c ({signal_3306, signal_1848}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1842 ( .a ({signal_3236, signal_1778}), .b ({signal_3315, signal_1857}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1853 ( .a ({signal_3253, signal_1795}), .b ({signal_3326, signal_1868}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1859 ( .a ({signal_3263, signal_1805}), .b ({signal_3332, signal_1874}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1860 ( .a ({signal_3265, signal_1807}), .b ({signal_3333, signal_1875}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1861 ( .a ({signal_3270, signal_1812}), .b ({signal_3334, signal_1876}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1862 ( .a ({signal_3274, signal_1816}), .b ({signal_3335, signal_1877}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1863 ( .a ({signal_3275, signal_1817}), .b ({signal_3336, signal_1878}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1864 ( .a ({signal_3279, signal_1821}), .b ({signal_3337, signal_1879}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1865 ( .a ({signal_3280, signal_1822}), .b ({signal_3338, signal_1880}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1866 ( .a ({signal_3281, signal_1823}), .b ({signal_3339, signal_1881}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1867 ( .a ({signal_3282, signal_1824}), .b ({signal_3340, signal_1882}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1868 ( .a ({signal_3286, signal_1828}), .b ({signal_3341, signal_1883}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1869 ( .a ({signal_3287, signal_1829}), .b ({signal_3342, signal_1884}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1870 ( .a ({signal_3289, signal_1831}), .b ({signal_3343, signal_1885}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1871 ( .a ({signal_3290, signal_1832}), .b ({signal_3344, signal_1886}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1873 ( .a ({signal_3300, signal_1842}), .b ({signal_3346, signal_1888}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1874 ( .a ({signal_3302, signal_1844}), .b ({signal_3347, signal_1889}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1876 ( .a ({signal_3173, signal_1715}), .b ({signal_5240, signal_5238}), .clk ( clk ), .r ( Fresh[527] ), .c ({signal_3349, signal_1891}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1877 ( .a ({signal_5248, signal_5244}), .b ({signal_3174, signal_1716}), .clk ( clk ), .r ( Fresh[528] ), .c ({signal_3350, signal_1892}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1878 ( .a ({signal_5252, signal_5250}), .b ({signal_3175, signal_1717}), .clk ( clk ), .r ( Fresh[529] ), .c ({signal_3351, signal_1893}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1879 ( .a ({signal_5068, signal_5066}), .b ({signal_3176, signal_1718}), .clk ( clk ), .r ( Fresh[530] ), .c ({signal_3352, signal_1894}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1880 ( .a ({signal_5108, signal_5106}), .b ({signal_3226, signal_1768}), .clk ( clk ), .r ( Fresh[531] ), .c ({signal_3353, signal_1895}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1881 ( .a ({signal_5260, signal_5256}), .b ({signal_3177, signal_1719}), .clk ( clk ), .r ( Fresh[532] ), .c ({signal_3354, signal_1896}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1882 ( .a ({signal_3178, signal_1720}), .b ({signal_5264, signal_5262}), .clk ( clk ), .r ( Fresh[533] ), .c ({signal_3355, signal_1897}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1883 ( .a ({signal_5268, signal_5266}), .b ({signal_3179, signal_1721}), .clk ( clk ), .r ( Fresh[534] ), .c ({signal_3356, signal_1898}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1884 ( .a ({signal_5272, signal_5270}), .b ({signal_3180, signal_1722}), .clk ( clk ), .r ( Fresh[535] ), .c ({signal_3357, signal_1899}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1885 ( .a ({signal_5284, signal_5278}), .b ({signal_3181, signal_1723}), .clk ( clk ), .r ( Fresh[536] ), .c ({signal_3358, signal_1900}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1886 ( .a ({signal_5080, signal_5078}), .b ({signal_3227, signal_1769}), .clk ( clk ), .r ( Fresh[537] ), .c ({signal_3359, signal_1901}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1887 ( .a ({signal_5288, signal_5286}), .b ({signal_3182, signal_1724}), .clk ( clk ), .r ( Fresh[538] ), .c ({signal_3360, signal_1902}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1888 ( .a ({signal_5292, signal_5290}), .b ({signal_3184, signal_1726}), .clk ( clk ), .r ( Fresh[539] ), .c ({signal_3361, signal_1903}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1889 ( .a ({signal_5296, signal_5294}), .b ({signal_3229, signal_1771}), .clk ( clk ), .r ( Fresh[540] ), .c ({signal_3362, signal_1904}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1890 ( .a ({signal_5068, signal_5066}), .b ({signal_3185, signal_1727}), .clk ( clk ), .r ( Fresh[541] ), .c ({signal_3363, signal_1905}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1891 ( .a ({signal_5108, signal_5106}), .b ({signal_3186, signal_1728}), .clk ( clk ), .r ( Fresh[542] ), .c ({signal_3364, signal_1906}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1892 ( .a ({signal_5300, signal_5298}), .b ({signal_3187, signal_1729}), .clk ( clk ), .r ( Fresh[543] ), .c ({signal_3365, signal_1907}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1894 ( .a ({signal_5116, signal_5114}), .b ({signal_3189, signal_1731}), .clk ( clk ), .r ( Fresh[544] ), .c ({signal_3367, signal_1909}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1895 ( .a ({signal_5308, signal_5304}), .b ({signal_3190, signal_1732}), .clk ( clk ), .r ( Fresh[545] ), .c ({signal_3368, signal_1910}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1896 ( .a ({signal_5312, signal_5310}), .b ({signal_3191, signal_1733}), .clk ( clk ), .r ( Fresh[546] ), .c ({signal_3369, signal_1911}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1897 ( .a ({signal_5316, signal_5314}), .b ({signal_3192, signal_1734}), .clk ( clk ), .r ( Fresh[547] ), .c ({signal_3370, signal_1912}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1898 ( .a ({signal_5320, signal_5318}), .b ({signal_3240, signal_1782}), .clk ( clk ), .r ( Fresh[548] ), .c ({signal_3371, signal_1913}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1899 ( .a ({signal_5324, signal_5322}), .b ({signal_3193, signal_1735}), .clk ( clk ), .r ( Fresh[549] ), .c ({signal_3372, signal_1914}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1900 ( .a ({signal_5292, signal_5290}), .b ({signal_3195, signal_1737}), .clk ( clk ), .r ( Fresh[550] ), .c ({signal_3373, signal_1915}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1901 ( .a ({signal_3196, signal_1738}), .b ({signal_3132, signal_1674}), .clk ( clk ), .r ( Fresh[551] ), .c ({signal_3374, signal_1916}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1903 ( .a ({signal_5072, signal_5070}), .b ({signal_3197, signal_1739}), .clk ( clk ), .r ( Fresh[552] ), .c ({signal_3376, signal_1918}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1905 ( .a ({signal_5312, signal_5310}), .b ({signal_3199, signal_1741}), .clk ( clk ), .r ( Fresh[553] ), .c ({signal_3378, signal_1920}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1906 ( .a ({signal_5104, signal_5102}), .b ({signal_3200, signal_1742}), .clk ( clk ), .r ( Fresh[554] ), .c ({signal_3379, signal_1921}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1907 ( .a ({signal_5204, signal_5202}), .b ({signal_3201, signal_1743}), .clk ( clk ), .r ( Fresh[555] ), .c ({signal_3380, signal_1922}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1908 ( .a ({signal_5260, signal_5256}), .b ({signal_3202, signal_1744}), .clk ( clk ), .r ( Fresh[556] ), .c ({signal_3381, signal_1923}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1909 ( .a ({signal_5328, signal_5326}), .b ({signal_3240, signal_1782}), .clk ( clk ), .r ( Fresh[557] ), .c ({signal_3382, signal_1924}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1910 ( .a ({signal_5332, signal_5330}), .b ({signal_3203, signal_1745}), .clk ( clk ), .r ( Fresh[558] ), .c ({signal_3383, signal_1925}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1913 ( .a ({signal_5336, signal_5334}), .b ({signal_3204, signal_1746}), .clk ( clk ), .r ( Fresh[559] ), .c ({signal_3386, signal_1928}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1914 ( .a ({signal_5104, signal_5102}), .b ({signal_3205, signal_1747}), .clk ( clk ), .r ( Fresh[560] ), .c ({signal_3387, signal_1929}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1915 ( .a ({signal_5068, signal_5066}), .b ({signal_3206, signal_1748}), .clk ( clk ), .r ( Fresh[561] ), .c ({signal_3388, signal_1930}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1916 ( .a ({signal_5340, signal_5338}), .b ({signal_3183, signal_1725}), .clk ( clk ), .r ( Fresh[562] ), .c ({signal_3389, signal_1931}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1917 ( .a ({signal_5344, signal_5342}), .b ({signal_3187, signal_1729}), .clk ( clk ), .r ( Fresh[563] ), .c ({signal_3390, signal_1932}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1919 ( .a ({signal_5352, signal_5348}), .b ({signal_3207, signal_1749}), .clk ( clk ), .r ( Fresh[564] ), .c ({signal_3392, signal_1934}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1920 ( .a ({signal_5204, signal_5202}), .b ({signal_3208, signal_1750}), .clk ( clk ), .r ( Fresh[565] ), .c ({signal_3393, signal_1935}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1923 ( .a ({signal_5356, signal_5354}), .b ({signal_3209, signal_1751}), .clk ( clk ), .r ( Fresh[566] ), .c ({signal_3396, signal_1938}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1927 ( .a ({signal_5360, signal_5358}), .b ({signal_3212, signal_1754}), .clk ( clk ), .r ( Fresh[567] ), .c ({signal_3400, signal_1942}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1932 ( .a ({signal_5064, signal_5062}), .b ({signal_3218, signal_1760}), .clk ( clk ), .r ( Fresh[568] ), .c ({signal_3405, signal_1947}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1944 ( .a ({signal_5364, signal_5362}), .b ({signal_3222, signal_1764}), .clk ( clk ), .r ( Fresh[569] ), .c ({signal_3417, signal_1959}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1948 ( .a ({signal_3350, signal_1892}), .b ({signal_3421, signal_1963}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1949 ( .a ({signal_3351, signal_1893}), .b ({signal_3422, signal_1964}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1950 ( .a ({signal_3353, signal_1895}), .b ({signal_3423, signal_1965}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1951 ( .a ({signal_3355, signal_1897}), .b ({signal_3424, signal_1966}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1952 ( .a ({signal_3356, signal_1898}), .b ({signal_3425, signal_1967}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1953 ( .a ({signal_3358, signal_1900}), .b ({signal_3426, signal_1968}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1954 ( .a ({signal_3359, signal_1901}), .b ({signal_3427, signal_1969}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1955 ( .a ({signal_3360, signal_1902}), .b ({signal_3428, signal_1970}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1956 ( .a ({signal_3361, signal_1903}), .b ({signal_3429, signal_1971}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1957 ( .a ({signal_3362, signal_1904}), .b ({signal_3430, signal_1972}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1958 ( .a ({signal_3363, signal_1905}), .b ({signal_3431, signal_1973}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1959 ( .a ({signal_3364, signal_1906}), .b ({signal_3432, signal_1974}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1960 ( .a ({signal_3365, signal_1907}), .b ({signal_3433, signal_1975}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1962 ( .a ({signal_3367, signal_1909}), .b ({signal_3435, signal_1977}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1963 ( .a ({signal_3368, signal_1910}), .b ({signal_3436, signal_1978}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1964 ( .a ({signal_3369, signal_1911}), .b ({signal_3437, signal_1979}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1965 ( .a ({signal_3370, signal_1912}), .b ({signal_3438, signal_1980}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1966 ( .a ({signal_3371, signal_1913}), .b ({signal_3439, signal_1981}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1967 ( .a ({signal_3372, signal_1914}), .b ({signal_3440, signal_1982}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1968 ( .a ({signal_3373, signal_1915}), .b ({signal_3441, signal_1983}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1970 ( .a ({signal_3376, signal_1918}), .b ({signal_3443, signal_1985}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1972 ( .a ({signal_3378, signal_1920}), .b ({signal_3445, signal_1987}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1973 ( .a ({signal_3379, signal_1921}), .b ({signal_3446, signal_1988}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1974 ( .a ({signal_3380, signal_1922}), .b ({signal_3447, signal_1989}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1975 ( .a ({signal_3381, signal_1923}), .b ({signal_3448, signal_1990}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1976 ( .a ({signal_3382, signal_1924}), .b ({signal_3449, signal_1991}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1977 ( .a ({signal_3383, signal_1925}), .b ({signal_3450, signal_1992}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1979 ( .a ({signal_3386, signal_1928}), .b ({signal_3452, signal_1994}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1980 ( .a ({signal_3387, signal_1929}), .b ({signal_3453, signal_1995}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1981 ( .a ({signal_3388, signal_1930}), .b ({signal_3454, signal_1996}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1982 ( .a ({signal_3389, signal_1931}), .b ({signal_3455, signal_1997}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1983 ( .a ({signal_3390, signal_1932}), .b ({signal_3456, signal_1998}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1984 ( .a ({signal_3392, signal_1934}), .b ({signal_3457, signal_1999}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1985 ( .a ({signal_3393, signal_1935}), .b ({signal_3458, signal_2000}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1988 ( .a ({signal_3396, signal_1938}), .b ({signal_3461, signal_2003}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1990 ( .a ({signal_3400, signal_1942}), .b ({signal_3463, signal_2005}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1991 ( .a ({signal_3405, signal_1947}), .b ({signal_3464, signal_2006}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1996 ( .a ({signal_3417, signal_1959}), .b ({signal_3469, signal_2011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2000 ( .a ({signal_3321, signal_1863}), .b ({signal_3052, signal_1594}), .clk ( clk ), .r ( Fresh[570] ), .c ({signal_3473, signal_2015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2001 ( .a ({signal_3310, signal_1852}), .b ({signal_3023, signal_1565}), .clk ( clk ), .r ( Fresh[571] ), .c ({signal_3474, signal_2016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2003 ( .a ({signal_3313, signal_1855}), .b ({signal_3314, signal_1856}), .clk ( clk ), .r ( Fresh[572] ), .c ({signal_3476, signal_2018}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2004 ( .a ({signal_5368, signal_5366}), .b ({signal_3316, signal_1858}), .clk ( clk ), .r ( Fresh[573] ), .c ({signal_3477, signal_2019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2005 ( .a ({signal_5212, signal_5210}), .b ({signal_3317, signal_1859}), .clk ( clk ), .r ( Fresh[574] ), .c ({signal_3478, signal_2020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2006 ( .a ({signal_5372, signal_5370}), .b ({signal_3318, signal_1860}), .clk ( clk ), .r ( Fresh[575] ), .c ({signal_3479, signal_2021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2008 ( .a ({signal_5376, signal_5374}), .b ({signal_3322, signal_1864}), .clk ( clk ), .r ( Fresh[576] ), .c ({signal_3481, signal_2023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2011 ( .a ({signal_5212, signal_5210}), .b ({signal_3323, signal_1865}), .clk ( clk ), .r ( Fresh[577] ), .c ({signal_3484, signal_2026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2012 ( .a ({signal_3067, signal_1609}), .b ({signal_3325, signal_1867}), .clk ( clk ), .r ( Fresh[578] ), .c ({signal_3485, signal_2027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2014 ( .a ({signal_3327, signal_1869}), .b ({signal_3146, signal_1688}), .clk ( clk ), .r ( Fresh[579] ), .c ({signal_3487, signal_2029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2015 ( .a ({signal_3065, signal_1607}), .b ({signal_3329, signal_1871}), .clk ( clk ), .r ( Fresh[580] ), .c ({signal_3488, signal_2030}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2048 ( .a ({signal_3477, signal_2019}), .b ({signal_3521, signal_2063}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2052 ( .a ({signal_3484, signal_2026}), .b ({signal_3525, signal_2067}) ) ;
    buf_clk cell_3018 ( .C ( clk ), .D ( signal_5377 ), .Q ( signal_5378 ) ) ;
    buf_clk cell_3020 ( .C ( clk ), .D ( signal_5379 ), .Q ( signal_5380 ) ) ;
    buf_clk cell_3022 ( .C ( clk ), .D ( signal_5381 ), .Q ( signal_5382 ) ) ;
    buf_clk cell_3024 ( .C ( clk ), .D ( signal_5383 ), .Q ( signal_5384 ) ) ;
    buf_clk cell_3028 ( .C ( clk ), .D ( signal_5387 ), .Q ( signal_5388 ) ) ;
    buf_clk cell_3032 ( .C ( clk ), .D ( signal_5391 ), .Q ( signal_5392 ) ) ;
    buf_clk cell_3034 ( .C ( clk ), .D ( signal_5393 ), .Q ( signal_5394 ) ) ;
    buf_clk cell_3036 ( .C ( clk ), .D ( signal_5395 ), .Q ( signal_5396 ) ) ;
    buf_clk cell_3040 ( .C ( clk ), .D ( signal_5399 ), .Q ( signal_5400 ) ) ;
    buf_clk cell_3044 ( .C ( clk ), .D ( signal_5403 ), .Q ( signal_5404 ) ) ;
    buf_clk cell_3048 ( .C ( clk ), .D ( signal_5407 ), .Q ( signal_5408 ) ) ;
    buf_clk cell_3052 ( .C ( clk ), .D ( signal_5411 ), .Q ( signal_5412 ) ) ;
    buf_clk cell_3056 ( .C ( clk ), .D ( signal_5415 ), .Q ( signal_5416 ) ) ;
    buf_clk cell_3060 ( .C ( clk ), .D ( signal_5419 ), .Q ( signal_5420 ) ) ;
    buf_clk cell_3068 ( .C ( clk ), .D ( signal_5427 ), .Q ( signal_5428 ) ) ;
    buf_clk cell_3076 ( .C ( clk ), .D ( signal_5435 ), .Q ( signal_5436 ) ) ;
    buf_clk cell_3078 ( .C ( clk ), .D ( signal_5437 ), .Q ( signal_5438 ) ) ;
    buf_clk cell_3080 ( .C ( clk ), .D ( signal_5439 ), .Q ( signal_5440 ) ) ;
    buf_clk cell_3082 ( .C ( clk ), .D ( signal_5441 ), .Q ( signal_5442 ) ) ;
    buf_clk cell_3084 ( .C ( clk ), .D ( signal_5443 ), .Q ( signal_5444 ) ) ;
    buf_clk cell_3088 ( .C ( clk ), .D ( signal_5447 ), .Q ( signal_5448 ) ) ;
    buf_clk cell_3092 ( .C ( clk ), .D ( signal_5451 ), .Q ( signal_5452 ) ) ;
    buf_clk cell_3094 ( .C ( clk ), .D ( signal_5453 ), .Q ( signal_5454 ) ) ;
    buf_clk cell_3096 ( .C ( clk ), .D ( signal_5455 ), .Q ( signal_5456 ) ) ;
    buf_clk cell_3098 ( .C ( clk ), .D ( signal_5457 ), .Q ( signal_5458 ) ) ;
    buf_clk cell_3100 ( .C ( clk ), .D ( signal_5459 ), .Q ( signal_5460 ) ) ;
    buf_clk cell_3104 ( .C ( clk ), .D ( signal_5463 ), .Q ( signal_5464 ) ) ;
    buf_clk cell_3108 ( .C ( clk ), .D ( signal_5467 ), .Q ( signal_5468 ) ) ;
    buf_clk cell_3110 ( .C ( clk ), .D ( signal_5469 ), .Q ( signal_5470 ) ) ;
    buf_clk cell_3112 ( .C ( clk ), .D ( signal_5471 ), .Q ( signal_5472 ) ) ;
    buf_clk cell_3114 ( .C ( clk ), .D ( signal_5473 ), .Q ( signal_5474 ) ) ;
    buf_clk cell_3116 ( .C ( clk ), .D ( signal_5475 ), .Q ( signal_5476 ) ) ;
    buf_clk cell_3118 ( .C ( clk ), .D ( signal_5477 ), .Q ( signal_5478 ) ) ;
    buf_clk cell_3120 ( .C ( clk ), .D ( signal_5479 ), .Q ( signal_5480 ) ) ;
    buf_clk cell_3122 ( .C ( clk ), .D ( signal_5481 ), .Q ( signal_5482 ) ) ;
    buf_clk cell_3124 ( .C ( clk ), .D ( signal_5483 ), .Q ( signal_5484 ) ) ;
    buf_clk cell_3126 ( .C ( clk ), .D ( signal_5485 ), .Q ( signal_5486 ) ) ;
    buf_clk cell_3128 ( .C ( clk ), .D ( signal_5487 ), .Q ( signal_5488 ) ) ;
    buf_clk cell_3132 ( .C ( clk ), .D ( signal_5491 ), .Q ( signal_5492 ) ) ;
    buf_clk cell_3136 ( .C ( clk ), .D ( signal_5495 ), .Q ( signal_5496 ) ) ;
    buf_clk cell_3138 ( .C ( clk ), .D ( signal_5497 ), .Q ( signal_5498 ) ) ;
    buf_clk cell_3140 ( .C ( clk ), .D ( signal_5499 ), .Q ( signal_5500 ) ) ;
    buf_clk cell_3142 ( .C ( clk ), .D ( signal_5501 ), .Q ( signal_5502 ) ) ;
    buf_clk cell_3144 ( .C ( clk ), .D ( signal_5503 ), .Q ( signal_5504 ) ) ;
    buf_clk cell_3146 ( .C ( clk ), .D ( signal_5505 ), .Q ( signal_5506 ) ) ;
    buf_clk cell_3148 ( .C ( clk ), .D ( signal_5507 ), .Q ( signal_5508 ) ) ;
    buf_clk cell_3150 ( .C ( clk ), .D ( signal_5509 ), .Q ( signal_5510 ) ) ;
    buf_clk cell_3152 ( .C ( clk ), .D ( signal_5511 ), .Q ( signal_5512 ) ) ;
    buf_clk cell_3156 ( .C ( clk ), .D ( signal_5515 ), .Q ( signal_5516 ) ) ;
    buf_clk cell_3160 ( .C ( clk ), .D ( signal_5519 ), .Q ( signal_5520 ) ) ;
    buf_clk cell_3162 ( .C ( clk ), .D ( signal_5521 ), .Q ( signal_5522 ) ) ;
    buf_clk cell_3164 ( .C ( clk ), .D ( signal_5523 ), .Q ( signal_5524 ) ) ;
    buf_clk cell_3166 ( .C ( clk ), .D ( signal_5525 ), .Q ( signal_5526 ) ) ;
    buf_clk cell_3168 ( .C ( clk ), .D ( signal_5527 ), .Q ( signal_5528 ) ) ;
    buf_clk cell_3172 ( .C ( clk ), .D ( signal_5531 ), .Q ( signal_5532 ) ) ;
    buf_clk cell_3176 ( .C ( clk ), .D ( signal_5535 ), .Q ( signal_5536 ) ) ;
    buf_clk cell_3180 ( .C ( clk ), .D ( signal_5539 ), .Q ( signal_5540 ) ) ;
    buf_clk cell_3184 ( .C ( clk ), .D ( signal_5543 ), .Q ( signal_5544 ) ) ;
    buf_clk cell_3188 ( .C ( clk ), .D ( signal_5547 ), .Q ( signal_5548 ) ) ;
    buf_clk cell_3192 ( .C ( clk ), .D ( signal_5551 ), .Q ( signal_5552 ) ) ;
    buf_clk cell_3196 ( .C ( clk ), .D ( signal_5555 ), .Q ( signal_5556 ) ) ;
    buf_clk cell_3200 ( .C ( clk ), .D ( signal_5559 ), .Q ( signal_5560 ) ) ;
    buf_clk cell_3202 ( .C ( clk ), .D ( signal_5561 ), .Q ( signal_5562 ) ) ;
    buf_clk cell_3204 ( .C ( clk ), .D ( signal_5563 ), .Q ( signal_5564 ) ) ;
    buf_clk cell_3206 ( .C ( clk ), .D ( signal_5565 ), .Q ( signal_5566 ) ) ;
    buf_clk cell_3208 ( .C ( clk ), .D ( signal_5567 ), .Q ( signal_5568 ) ) ;
    buf_clk cell_3210 ( .C ( clk ), .D ( signal_5569 ), .Q ( signal_5570 ) ) ;
    buf_clk cell_3212 ( .C ( clk ), .D ( signal_5571 ), .Q ( signal_5572 ) ) ;
    buf_clk cell_3214 ( .C ( clk ), .D ( signal_5573 ), .Q ( signal_5574 ) ) ;
    buf_clk cell_3216 ( .C ( clk ), .D ( signal_5575 ), .Q ( signal_5576 ) ) ;
    buf_clk cell_3218 ( .C ( clk ), .D ( signal_5577 ), .Q ( signal_5578 ) ) ;
    buf_clk cell_3220 ( .C ( clk ), .D ( signal_5579 ), .Q ( signal_5580 ) ) ;
    buf_clk cell_3224 ( .C ( clk ), .D ( signal_5583 ), .Q ( signal_5584 ) ) ;
    buf_clk cell_3228 ( .C ( clk ), .D ( signal_5587 ), .Q ( signal_5588 ) ) ;
    buf_clk cell_3232 ( .C ( clk ), .D ( signal_5591 ), .Q ( signal_5592 ) ) ;
    buf_clk cell_3236 ( .C ( clk ), .D ( signal_5595 ), .Q ( signal_5596 ) ) ;
    buf_clk cell_3240 ( .C ( clk ), .D ( signal_5599 ), .Q ( signal_5600 ) ) ;
    buf_clk cell_3244 ( .C ( clk ), .D ( signal_5603 ), .Q ( signal_5604 ) ) ;
    buf_clk cell_3246 ( .C ( clk ), .D ( signal_5605 ), .Q ( signal_5606 ) ) ;
    buf_clk cell_3248 ( .C ( clk ), .D ( signal_5607 ), .Q ( signal_5608 ) ) ;
    buf_clk cell_3252 ( .C ( clk ), .D ( signal_5611 ), .Q ( signal_5612 ) ) ;
    buf_clk cell_3256 ( .C ( clk ), .D ( signal_5615 ), .Q ( signal_5616 ) ) ;
    buf_clk cell_3258 ( .C ( clk ), .D ( signal_5617 ), .Q ( signal_5618 ) ) ;
    buf_clk cell_3260 ( .C ( clk ), .D ( signal_5619 ), .Q ( signal_5620 ) ) ;
    buf_clk cell_3262 ( .C ( clk ), .D ( signal_5621 ), .Q ( signal_5622 ) ) ;
    buf_clk cell_3264 ( .C ( clk ), .D ( signal_5623 ), .Q ( signal_5624 ) ) ;
    buf_clk cell_3266 ( .C ( clk ), .D ( signal_5625 ), .Q ( signal_5626 ) ) ;
    buf_clk cell_3268 ( .C ( clk ), .D ( signal_5627 ), .Q ( signal_5628 ) ) ;
    buf_clk cell_3270 ( .C ( clk ), .D ( signal_5629 ), .Q ( signal_5630 ) ) ;
    buf_clk cell_3272 ( .C ( clk ), .D ( signal_5631 ), .Q ( signal_5632 ) ) ;
    buf_clk cell_3274 ( .C ( clk ), .D ( signal_5633 ), .Q ( signal_5634 ) ) ;
    buf_clk cell_3276 ( .C ( clk ), .D ( signal_5635 ), .Q ( signal_5636 ) ) ;
    buf_clk cell_3280 ( .C ( clk ), .D ( signal_5639 ), .Q ( signal_5640 ) ) ;
    buf_clk cell_3284 ( .C ( clk ), .D ( signal_5643 ), .Q ( signal_5644 ) ) ;
    buf_clk cell_3288 ( .C ( clk ), .D ( signal_5647 ), .Q ( signal_5648 ) ) ;
    buf_clk cell_3292 ( .C ( clk ), .D ( signal_5651 ), .Q ( signal_5652 ) ) ;
    buf_clk cell_3294 ( .C ( clk ), .D ( signal_5653 ), .Q ( signal_5654 ) ) ;
    buf_clk cell_3296 ( .C ( clk ), .D ( signal_5655 ), .Q ( signal_5656 ) ) ;
    buf_clk cell_3300 ( .C ( clk ), .D ( signal_5659 ), .Q ( signal_5660 ) ) ;
    buf_clk cell_3304 ( .C ( clk ), .D ( signal_5663 ), .Q ( signal_5664 ) ) ;
    buf_clk cell_3306 ( .C ( clk ), .D ( signal_5665 ), .Q ( signal_5666 ) ) ;
    buf_clk cell_3308 ( .C ( clk ), .D ( signal_5667 ), .Q ( signal_5668 ) ) ;
    buf_clk cell_3310 ( .C ( clk ), .D ( signal_5669 ), .Q ( signal_5670 ) ) ;
    buf_clk cell_3312 ( .C ( clk ), .D ( signal_5671 ), .Q ( signal_5672 ) ) ;
    buf_clk cell_3316 ( .C ( clk ), .D ( signal_5675 ), .Q ( signal_5676 ) ) ;
    buf_clk cell_3320 ( .C ( clk ), .D ( signal_5679 ), .Q ( signal_5680 ) ) ;
    buf_clk cell_3324 ( .C ( clk ), .D ( signal_5683 ), .Q ( signal_5684 ) ) ;
    buf_clk cell_3328 ( .C ( clk ), .D ( signal_5687 ), .Q ( signal_5688 ) ) ;
    buf_clk cell_3332 ( .C ( clk ), .D ( signal_5691 ), .Q ( signal_5692 ) ) ;
    buf_clk cell_3336 ( .C ( clk ), .D ( signal_5695 ), .Q ( signal_5696 ) ) ;
    buf_clk cell_3338 ( .C ( clk ), .D ( signal_5697 ), .Q ( signal_5698 ) ) ;
    buf_clk cell_3340 ( .C ( clk ), .D ( signal_5699 ), .Q ( signal_5700 ) ) ;
    buf_clk cell_3344 ( .C ( clk ), .D ( signal_5703 ), .Q ( signal_5704 ) ) ;
    buf_clk cell_3348 ( .C ( clk ), .D ( signal_5707 ), .Q ( signal_5708 ) ) ;
    buf_clk cell_3352 ( .C ( clk ), .D ( signal_5711 ), .Q ( signal_5712 ) ) ;
    buf_clk cell_3356 ( .C ( clk ), .D ( signal_5715 ), .Q ( signal_5716 ) ) ;
    buf_clk cell_3358 ( .C ( clk ), .D ( signal_5717 ), .Q ( signal_5718 ) ) ;
    buf_clk cell_3360 ( .C ( clk ), .D ( signal_5719 ), .Q ( signal_5720 ) ) ;
    buf_clk cell_3364 ( .C ( clk ), .D ( signal_5723 ), .Q ( signal_5724 ) ) ;
    buf_clk cell_3368 ( .C ( clk ), .D ( signal_5727 ), .Q ( signal_5728 ) ) ;
    buf_clk cell_3370 ( .C ( clk ), .D ( signal_5729 ), .Q ( signal_5730 ) ) ;
    buf_clk cell_3372 ( .C ( clk ), .D ( signal_5731 ), .Q ( signal_5732 ) ) ;
    buf_clk cell_3374 ( .C ( clk ), .D ( signal_5733 ), .Q ( signal_5734 ) ) ;
    buf_clk cell_3376 ( .C ( clk ), .D ( signal_5735 ), .Q ( signal_5736 ) ) ;
    buf_clk cell_3378 ( .C ( clk ), .D ( signal_5737 ), .Q ( signal_5738 ) ) ;
    buf_clk cell_3380 ( .C ( clk ), .D ( signal_5739 ), .Q ( signal_5740 ) ) ;
    buf_clk cell_3384 ( .C ( clk ), .D ( signal_5743 ), .Q ( signal_5744 ) ) ;
    buf_clk cell_3388 ( .C ( clk ), .D ( signal_5747 ), .Q ( signal_5748 ) ) ;
    buf_clk cell_3396 ( .C ( clk ), .D ( signal_5755 ), .Q ( signal_5756 ) ) ;
    buf_clk cell_3402 ( .C ( clk ), .D ( signal_5761 ), .Q ( signal_5762 ) ) ;
    buf_clk cell_3408 ( .C ( clk ), .D ( signal_5767 ), .Q ( signal_5768 ) ) ;
    buf_clk cell_3414 ( .C ( clk ), .D ( signal_5773 ), .Q ( signal_5774 ) ) ;
    buf_clk cell_3420 ( .C ( clk ), .D ( signal_5779 ), .Q ( signal_5780 ) ) ;
    buf_clk cell_3426 ( .C ( clk ), .D ( signal_5785 ), .Q ( signal_5786 ) ) ;
    buf_clk cell_3430 ( .C ( clk ), .D ( signal_5789 ), .Q ( signal_5790 ) ) ;
    buf_clk cell_3434 ( .C ( clk ), .D ( signal_5793 ), .Q ( signal_5794 ) ) ;
    buf_clk cell_3440 ( .C ( clk ), .D ( signal_5799 ), .Q ( signal_5800 ) ) ;
    buf_clk cell_3446 ( .C ( clk ), .D ( signal_5805 ), .Q ( signal_5806 ) ) ;
    buf_clk cell_3450 ( .C ( clk ), .D ( signal_5809 ), .Q ( signal_5810 ) ) ;
    buf_clk cell_3454 ( .C ( clk ), .D ( signal_5813 ), .Q ( signal_5814 ) ) ;
    buf_clk cell_3458 ( .C ( clk ), .D ( signal_5817 ), .Q ( signal_5818 ) ) ;
    buf_clk cell_3462 ( .C ( clk ), .D ( signal_5821 ), .Q ( signal_5822 ) ) ;
    buf_clk cell_3466 ( .C ( clk ), .D ( signal_5825 ), .Q ( signal_5826 ) ) ;
    buf_clk cell_3470 ( .C ( clk ), .D ( signal_5829 ), .Q ( signal_5830 ) ) ;
    buf_clk cell_3474 ( .C ( clk ), .D ( signal_5833 ), .Q ( signal_5834 ) ) ;
    buf_clk cell_3478 ( .C ( clk ), .D ( signal_5837 ), .Q ( signal_5838 ) ) ;
    buf_clk cell_3482 ( .C ( clk ), .D ( signal_5841 ), .Q ( signal_5842 ) ) ;
    buf_clk cell_3486 ( .C ( clk ), .D ( signal_5845 ), .Q ( signal_5846 ) ) ;
    buf_clk cell_3492 ( .C ( clk ), .D ( signal_5851 ), .Q ( signal_5852 ) ) ;
    buf_clk cell_3498 ( .C ( clk ), .D ( signal_5857 ), .Q ( signal_5858 ) ) ;
    buf_clk cell_3502 ( .C ( clk ), .D ( signal_5861 ), .Q ( signal_5862 ) ) ;
    buf_clk cell_3506 ( .C ( clk ), .D ( signal_5865 ), .Q ( signal_5866 ) ) ;
    buf_clk cell_3530 ( .C ( clk ), .D ( signal_5889 ), .Q ( signal_5890 ) ) ;
    buf_clk cell_3534 ( .C ( clk ), .D ( signal_5893 ), .Q ( signal_5894 ) ) ;
    buf_clk cell_3552 ( .C ( clk ), .D ( signal_5911 ), .Q ( signal_5912 ) ) ;
    buf_clk cell_3558 ( .C ( clk ), .D ( signal_5917 ), .Q ( signal_5918 ) ) ;
    buf_clk cell_3566 ( .C ( clk ), .D ( signal_5925 ), .Q ( signal_5926 ) ) ;
    buf_clk cell_3570 ( .C ( clk ), .D ( signal_5929 ), .Q ( signal_5930 ) ) ;
    buf_clk cell_3584 ( .C ( clk ), .D ( signal_5943 ), .Q ( signal_5944 ) ) ;
    buf_clk cell_3590 ( .C ( clk ), .D ( signal_5949 ), .Q ( signal_5950 ) ) ;
    buf_clk cell_3594 ( .C ( clk ), .D ( signal_5953 ), .Q ( signal_5954 ) ) ;
    buf_clk cell_3598 ( .C ( clk ), .D ( signal_5957 ), .Q ( signal_5958 ) ) ;
    buf_clk cell_3610 ( .C ( clk ), .D ( signal_5969 ), .Q ( signal_5970 ) ) ;
    buf_clk cell_3614 ( .C ( clk ), .D ( signal_5973 ), .Q ( signal_5974 ) ) ;
    buf_clk cell_3618 ( .C ( clk ), .D ( signal_5977 ), .Q ( signal_5978 ) ) ;
    buf_clk cell_3622 ( .C ( clk ), .D ( signal_5981 ), .Q ( signal_5982 ) ) ;
    buf_clk cell_3626 ( .C ( clk ), .D ( signal_5985 ), .Q ( signal_5986 ) ) ;
    buf_clk cell_3630 ( .C ( clk ), .D ( signal_5989 ), .Q ( signal_5990 ) ) ;
    buf_clk cell_3640 ( .C ( clk ), .D ( signal_5999 ), .Q ( signal_6000 ) ) ;
    buf_clk cell_3646 ( .C ( clk ), .D ( signal_6005 ), .Q ( signal_6006 ) ) ;
    buf_clk cell_3650 ( .C ( clk ), .D ( signal_6009 ), .Q ( signal_6010 ) ) ;
    buf_clk cell_3654 ( .C ( clk ), .D ( signal_6013 ), .Q ( signal_6014 ) ) ;
    buf_clk cell_3660 ( .C ( clk ), .D ( signal_6019 ), .Q ( signal_6020 ) ) ;
    buf_clk cell_3666 ( .C ( clk ), .D ( signal_6025 ), .Q ( signal_6026 ) ) ;
    buf_clk cell_3670 ( .C ( clk ), .D ( signal_6029 ), .Q ( signal_6030 ) ) ;
    buf_clk cell_3674 ( .C ( clk ), .D ( signal_6033 ), .Q ( signal_6034 ) ) ;
    buf_clk cell_3678 ( .C ( clk ), .D ( signal_6037 ), .Q ( signal_6038 ) ) ;
    buf_clk cell_3682 ( .C ( clk ), .D ( signal_6041 ), .Q ( signal_6042 ) ) ;
    buf_clk cell_3686 ( .C ( clk ), .D ( signal_6045 ), .Q ( signal_6046 ) ) ;
    buf_clk cell_3690 ( .C ( clk ), .D ( signal_6049 ), .Q ( signal_6050 ) ) ;
    buf_clk cell_3698 ( .C ( clk ), .D ( signal_6057 ), .Q ( signal_6058 ) ) ;
    buf_clk cell_3702 ( .C ( clk ), .D ( signal_6061 ), .Q ( signal_6062 ) ) ;
    buf_clk cell_3706 ( .C ( clk ), .D ( signal_6065 ), .Q ( signal_6066 ) ) ;
    buf_clk cell_3710 ( .C ( clk ), .D ( signal_6069 ), .Q ( signal_6070 ) ) ;
    buf_clk cell_3716 ( .C ( clk ), .D ( signal_6075 ), .Q ( signal_6076 ) ) ;
    buf_clk cell_3722 ( .C ( clk ), .D ( signal_6081 ), .Q ( signal_6082 ) ) ;
    buf_clk cell_3734 ( .C ( clk ), .D ( signal_6093 ), .Q ( signal_6094 ) ) ;
    buf_clk cell_3738 ( .C ( clk ), .D ( signal_6097 ), .Q ( signal_6098 ) ) ;
    buf_clk cell_3744 ( .C ( clk ), .D ( signal_6103 ), .Q ( signal_6104 ) ) ;
    buf_clk cell_3750 ( .C ( clk ), .D ( signal_6109 ), .Q ( signal_6110 ) ) ;
    buf_clk cell_3756 ( .C ( clk ), .D ( signal_6115 ), .Q ( signal_6116 ) ) ;
    buf_clk cell_3762 ( .C ( clk ), .D ( signal_6121 ), .Q ( signal_6122 ) ) ;
    buf_clk cell_3768 ( .C ( clk ), .D ( signal_6127 ), .Q ( signal_6128 ) ) ;
    buf_clk cell_3774 ( .C ( clk ), .D ( signal_6133 ), .Q ( signal_6134 ) ) ;
    buf_clk cell_3778 ( .C ( clk ), .D ( signal_6137 ), .Q ( signal_6138 ) ) ;
    buf_clk cell_3782 ( .C ( clk ), .D ( signal_6141 ), .Q ( signal_6142 ) ) ;
    buf_clk cell_3796 ( .C ( clk ), .D ( signal_6155 ), .Q ( signal_6156 ) ) ;
    buf_clk cell_3804 ( .C ( clk ), .D ( signal_6163 ), .Q ( signal_6164 ) ) ;
    buf_clk cell_3818 ( .C ( clk ), .D ( signal_6177 ), .Q ( signal_6178 ) ) ;
    buf_clk cell_3824 ( .C ( clk ), .D ( signal_6183 ), .Q ( signal_6184 ) ) ;
    buf_clk cell_3830 ( .C ( clk ), .D ( signal_6189 ), .Q ( signal_6190 ) ) ;
    buf_clk cell_3836 ( .C ( clk ), .D ( signal_6195 ), .Q ( signal_6196 ) ) ;
    buf_clk cell_3850 ( .C ( clk ), .D ( signal_6209 ), .Q ( signal_6210 ) ) ;
    buf_clk cell_3856 ( .C ( clk ), .D ( signal_6215 ), .Q ( signal_6216 ) ) ;
    buf_clk cell_3886 ( .C ( clk ), .D ( signal_6245 ), .Q ( signal_6246 ) ) ;
    buf_clk cell_3892 ( .C ( clk ), .D ( signal_6251 ), .Q ( signal_6252 ) ) ;
    buf_clk cell_3898 ( .C ( clk ), .D ( signal_6257 ), .Q ( signal_6258 ) ) ;
    buf_clk cell_3904 ( .C ( clk ), .D ( signal_6263 ), .Q ( signal_6264 ) ) ;
    buf_clk cell_3910 ( .C ( clk ), .D ( signal_6269 ), .Q ( signal_6270 ) ) ;
    buf_clk cell_3916 ( .C ( clk ), .D ( signal_6275 ), .Q ( signal_6276 ) ) ;
    buf_clk cell_3934 ( .C ( clk ), .D ( signal_6293 ), .Q ( signal_6294 ) ) ;
    buf_clk cell_3940 ( .C ( clk ), .D ( signal_6299 ), .Q ( signal_6300 ) ) ;
    buf_clk cell_3950 ( .C ( clk ), .D ( signal_6309 ), .Q ( signal_6310 ) ) ;
    buf_clk cell_3956 ( .C ( clk ), .D ( signal_6315 ), .Q ( signal_6316 ) ) ;
    buf_clk cell_3968 ( .C ( clk ), .D ( signal_6327 ), .Q ( signal_6328 ) ) ;
    buf_clk cell_3976 ( .C ( clk ), .D ( signal_6335 ), .Q ( signal_6336 ) ) ;
    buf_clk cell_3998 ( .C ( clk ), .D ( signal_6357 ), .Q ( signal_6358 ) ) ;
    buf_clk cell_4004 ( .C ( clk ), .D ( signal_6363 ), .Q ( signal_6364 ) ) ;
    buf_clk cell_4010 ( .C ( clk ), .D ( signal_6369 ), .Q ( signal_6370 ) ) ;
    buf_clk cell_4016 ( .C ( clk ), .D ( signal_6375 ), .Q ( signal_6376 ) ) ;
    buf_clk cell_4032 ( .C ( clk ), .D ( signal_6391 ), .Q ( signal_6392 ) ) ;
    buf_clk cell_4040 ( .C ( clk ), .D ( signal_6399 ), .Q ( signal_6400 ) ) ;
    buf_clk cell_4046 ( .C ( clk ), .D ( signal_6405 ), .Q ( signal_6406 ) ) ;
    buf_clk cell_4052 ( .C ( clk ), .D ( signal_6411 ), .Q ( signal_6412 ) ) ;
    buf_clk cell_4058 ( .C ( clk ), .D ( signal_6417 ), .Q ( signal_6418 ) ) ;
    buf_clk cell_4064 ( .C ( clk ), .D ( signal_6423 ), .Q ( signal_6424 ) ) ;
    buf_clk cell_4078 ( .C ( clk ), .D ( signal_6437 ), .Q ( signal_6438 ) ) ;
    buf_clk cell_4084 ( .C ( clk ), .D ( signal_6443 ), .Q ( signal_6444 ) ) ;
    buf_clk cell_4098 ( .C ( clk ), .D ( signal_6457 ), .Q ( signal_6458 ) ) ;
    buf_clk cell_4104 ( .C ( clk ), .D ( signal_6463 ), .Q ( signal_6464 ) ) ;
    buf_clk cell_4110 ( .C ( clk ), .D ( signal_6469 ), .Q ( signal_6470 ) ) ;
    buf_clk cell_4116 ( .C ( clk ), .D ( signal_6475 ), .Q ( signal_6476 ) ) ;
    buf_clk cell_4132 ( .C ( clk ), .D ( signal_6491 ), .Q ( signal_6492 ) ) ;
    buf_clk cell_4142 ( .C ( clk ), .D ( signal_6501 ), .Q ( signal_6502 ) ) ;
    buf_clk cell_4162 ( .C ( clk ), .D ( signal_6521 ), .Q ( signal_6522 ) ) ;
    buf_clk cell_4170 ( .C ( clk ), .D ( signal_6529 ), .Q ( signal_6530 ) ) ;
    buf_clk cell_4178 ( .C ( clk ), .D ( signal_6537 ), .Q ( signal_6538 ) ) ;
    buf_clk cell_4186 ( .C ( clk ), .D ( signal_6545 ), .Q ( signal_6546 ) ) ;
    buf_clk cell_4228 ( .C ( clk ), .D ( signal_6587 ), .Q ( signal_6588 ) ) ;
    buf_clk cell_4238 ( .C ( clk ), .D ( signal_6597 ), .Q ( signal_6598 ) ) ;
    buf_clk cell_4262 ( .C ( clk ), .D ( signal_6621 ), .Q ( signal_6622 ) ) ;
    buf_clk cell_4270 ( .C ( clk ), .D ( signal_6629 ), .Q ( signal_6630 ) ) ;
    buf_clk cell_4290 ( .C ( clk ), .D ( signal_6649 ), .Q ( signal_6650 ) ) ;
    buf_clk cell_4298 ( .C ( clk ), .D ( signal_6657 ), .Q ( signal_6658 ) ) ;
    buf_clk cell_4306 ( .C ( clk ), .D ( signal_6665 ), .Q ( signal_6666 ) ) ;
    buf_clk cell_4314 ( .C ( clk ), .D ( signal_6673 ), .Q ( signal_6674 ) ) ;
    buf_clk cell_4322 ( .C ( clk ), .D ( signal_6681 ), .Q ( signal_6682 ) ) ;
    buf_clk cell_4330 ( .C ( clk ), .D ( signal_6689 ), .Q ( signal_6690 ) ) ;
    buf_clk cell_4340 ( .C ( clk ), .D ( signal_6699 ), .Q ( signal_6700 ) ) ;
    buf_clk cell_4350 ( .C ( clk ), .D ( signal_6709 ), .Q ( signal_6710 ) ) ;
    buf_clk cell_4358 ( .C ( clk ), .D ( signal_6717 ), .Q ( signal_6718 ) ) ;
    buf_clk cell_4366 ( .C ( clk ), .D ( signal_6725 ), .Q ( signal_6726 ) ) ;
    buf_clk cell_4374 ( .C ( clk ), .D ( signal_6733 ), .Q ( signal_6734 ) ) ;
    buf_clk cell_4382 ( .C ( clk ), .D ( signal_6741 ), .Q ( signal_6742 ) ) ;
    buf_clk cell_4394 ( .C ( clk ), .D ( signal_6753 ), .Q ( signal_6754 ) ) ;
    buf_clk cell_4402 ( .C ( clk ), .D ( signal_6761 ), .Q ( signal_6762 ) ) ;
    buf_clk cell_4410 ( .C ( clk ), .D ( signal_6769 ), .Q ( signal_6770 ) ) ;
    buf_clk cell_4418 ( .C ( clk ), .D ( signal_6777 ), .Q ( signal_6778 ) ) ;
    buf_clk cell_4426 ( .C ( clk ), .D ( signal_6785 ), .Q ( signal_6786 ) ) ;
    buf_clk cell_4434 ( .C ( clk ), .D ( signal_6793 ), .Q ( signal_6794 ) ) ;
    buf_clk cell_4510 ( .C ( clk ), .D ( signal_6869 ), .Q ( signal_6870 ) ) ;
    buf_clk cell_4520 ( .C ( clk ), .D ( signal_6879 ), .Q ( signal_6880 ) ) ;
    buf_clk cell_4562 ( .C ( clk ), .D ( signal_6921 ), .Q ( signal_6922 ) ) ;
    buf_clk cell_4572 ( .C ( clk ), .D ( signal_6931 ), .Q ( signal_6932 ) ) ;
    buf_clk cell_4966 ( .C ( clk ), .D ( signal_7325 ), .Q ( signal_7326 ) ) ;
    buf_clk cell_4980 ( .C ( clk ), .D ( signal_7339 ), .Q ( signal_7340 ) ) ;
    buf_clk cell_5010 ( .C ( clk ), .D ( signal_7369 ), .Q ( signal_7370 ) ) ;
    buf_clk cell_5024 ( .C ( clk ), .D ( signal_7383 ), .Q ( signal_7384 ) ) ;
    buf_clk cell_5090 ( .C ( clk ), .D ( signal_7449 ), .Q ( signal_7450 ) ) ;
    buf_clk cell_5106 ( .C ( clk ), .D ( signal_7465 ), .Q ( signal_7466 ) ) ;
    buf_clk cell_5130 ( .C ( clk ), .D ( signal_7489 ), .Q ( signal_7490 ) ) ;
    buf_clk cell_5146 ( .C ( clk ), .D ( signal_7505 ), .Q ( signal_7506 ) ) ;
    buf_clk cell_5286 ( .C ( clk ), .D ( signal_7645 ), .Q ( signal_7646 ) ) ;
    buf_clk cell_5304 ( .C ( clk ), .D ( signal_7663 ), .Q ( signal_7664 ) ) ;
    buf_clk cell_5386 ( .C ( clk ), .D ( signal_7745 ), .Q ( signal_7746 ) ) ;
    buf_clk cell_5406 ( .C ( clk ), .D ( signal_7765 ), .Q ( signal_7766 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_3389 ( .C ( clk ), .D ( signal_5666 ), .Q ( signal_5749 ) ) ;
    buf_clk cell_3391 ( .C ( clk ), .D ( signal_5668 ), .Q ( signal_5751 ) ) ;
    buf_clk cell_3397 ( .C ( clk ), .D ( signal_5756 ), .Q ( signal_5757 ) ) ;
    buf_clk cell_3403 ( .C ( clk ), .D ( signal_5762 ), .Q ( signal_5763 ) ) ;
    buf_clk cell_3409 ( .C ( clk ), .D ( signal_5768 ), .Q ( signal_5769 ) ) ;
    buf_clk cell_3415 ( .C ( clk ), .D ( signal_5774 ), .Q ( signal_5775 ) ) ;
    buf_clk cell_3421 ( .C ( clk ), .D ( signal_5780 ), .Q ( signal_5781 ) ) ;
    buf_clk cell_3427 ( .C ( clk ), .D ( signal_5786 ), .Q ( signal_5787 ) ) ;
    buf_clk cell_3431 ( .C ( clk ), .D ( signal_5790 ), .Q ( signal_5791 ) ) ;
    buf_clk cell_3435 ( .C ( clk ), .D ( signal_5794 ), .Q ( signal_5795 ) ) ;
    buf_clk cell_3441 ( .C ( clk ), .D ( signal_5800 ), .Q ( signal_5801 ) ) ;
    buf_clk cell_3447 ( .C ( clk ), .D ( signal_5806 ), .Q ( signal_5807 ) ) ;
    buf_clk cell_3451 ( .C ( clk ), .D ( signal_5810 ), .Q ( signal_5811 ) ) ;
    buf_clk cell_3455 ( .C ( clk ), .D ( signal_5814 ), .Q ( signal_5815 ) ) ;
    buf_clk cell_3459 ( .C ( clk ), .D ( signal_5818 ), .Q ( signal_5819 ) ) ;
    buf_clk cell_3463 ( .C ( clk ), .D ( signal_5822 ), .Q ( signal_5823 ) ) ;
    buf_clk cell_3467 ( .C ( clk ), .D ( signal_5826 ), .Q ( signal_5827 ) ) ;
    buf_clk cell_3471 ( .C ( clk ), .D ( signal_5830 ), .Q ( signal_5831 ) ) ;
    buf_clk cell_3475 ( .C ( clk ), .D ( signal_5834 ), .Q ( signal_5835 ) ) ;
    buf_clk cell_3479 ( .C ( clk ), .D ( signal_5838 ), .Q ( signal_5839 ) ) ;
    buf_clk cell_3483 ( .C ( clk ), .D ( signal_5842 ), .Q ( signal_5843 ) ) ;
    buf_clk cell_3487 ( .C ( clk ), .D ( signal_5846 ), .Q ( signal_5847 ) ) ;
    buf_clk cell_3493 ( .C ( clk ), .D ( signal_5852 ), .Q ( signal_5853 ) ) ;
    buf_clk cell_3499 ( .C ( clk ), .D ( signal_5858 ), .Q ( signal_5859 ) ) ;
    buf_clk cell_3503 ( .C ( clk ), .D ( signal_5862 ), .Q ( signal_5863 ) ) ;
    buf_clk cell_3507 ( .C ( clk ), .D ( signal_5866 ), .Q ( signal_5867 ) ) ;
    buf_clk cell_3509 ( .C ( clk ), .D ( signal_1999 ), .Q ( signal_5869 ) ) ;
    buf_clk cell_3511 ( .C ( clk ), .D ( signal_3457 ), .Q ( signal_5871 ) ) ;
    buf_clk cell_3513 ( .C ( clk ), .D ( signal_5574 ), .Q ( signal_5873 ) ) ;
    buf_clk cell_3515 ( .C ( clk ), .D ( signal_5576 ), .Q ( signal_5875 ) ) ;
    buf_clk cell_3517 ( .C ( clk ), .D ( signal_1811 ), .Q ( signal_5877 ) ) ;
    buf_clk cell_3519 ( .C ( clk ), .D ( signal_3269 ), .Q ( signal_5879 ) ) ;
    buf_clk cell_3521 ( .C ( clk ), .D ( signal_1980 ), .Q ( signal_5881 ) ) ;
    buf_clk cell_3523 ( .C ( clk ), .D ( signal_3438 ), .Q ( signal_5883 ) ) ;
    buf_clk cell_3525 ( .C ( clk ), .D ( signal_1983 ), .Q ( signal_5885 ) ) ;
    buf_clk cell_3527 ( .C ( clk ), .D ( signal_3441 ), .Q ( signal_5887 ) ) ;
    buf_clk cell_3531 ( .C ( clk ), .D ( signal_5890 ), .Q ( signal_5891 ) ) ;
    buf_clk cell_3535 ( .C ( clk ), .D ( signal_5894 ), .Q ( signal_5895 ) ) ;
    buf_clk cell_3537 ( .C ( clk ), .D ( signal_1965 ), .Q ( signal_5897 ) ) ;
    buf_clk cell_3539 ( .C ( clk ), .D ( signal_3423 ), .Q ( signal_5899 ) ) ;
    buf_clk cell_3541 ( .C ( clk ), .D ( signal_1968 ), .Q ( signal_5901 ) ) ;
    buf_clk cell_3543 ( .C ( clk ), .D ( signal_3426 ), .Q ( signal_5903 ) ) ;
    buf_clk cell_3545 ( .C ( clk ), .D ( signal_5618 ), .Q ( signal_5905 ) ) ;
    buf_clk cell_3547 ( .C ( clk ), .D ( signal_5620 ), .Q ( signal_5907 ) ) ;
    buf_clk cell_3553 ( .C ( clk ), .D ( signal_5912 ), .Q ( signal_5913 ) ) ;
    buf_clk cell_3559 ( .C ( clk ), .D ( signal_5918 ), .Q ( signal_5919 ) ) ;
    buf_clk cell_3561 ( .C ( clk ), .D ( signal_1970 ), .Q ( signal_5921 ) ) ;
    buf_clk cell_3563 ( .C ( clk ), .D ( signal_3428 ), .Q ( signal_5923 ) ) ;
    buf_clk cell_3567 ( .C ( clk ), .D ( signal_5926 ), .Q ( signal_5927 ) ) ;
    buf_clk cell_3571 ( .C ( clk ), .D ( signal_5930 ), .Q ( signal_5931 ) ) ;
    buf_clk cell_3573 ( .C ( clk ), .D ( signal_5548 ), .Q ( signal_5933 ) ) ;
    buf_clk cell_3575 ( .C ( clk ), .D ( signal_5552 ), .Q ( signal_5935 ) ) ;
    buf_clk cell_3577 ( .C ( clk ), .D ( signal_5626 ), .Q ( signal_5937 ) ) ;
    buf_clk cell_3579 ( .C ( clk ), .D ( signal_5628 ), .Q ( signal_5939 ) ) ;
    buf_clk cell_3585 ( .C ( clk ), .D ( signal_5944 ), .Q ( signal_5945 ) ) ;
    buf_clk cell_3591 ( .C ( clk ), .D ( signal_5950 ), .Q ( signal_5951 ) ) ;
    buf_clk cell_3595 ( .C ( clk ), .D ( signal_5954 ), .Q ( signal_5955 ) ) ;
    buf_clk cell_3599 ( .C ( clk ), .D ( signal_5958 ), .Q ( signal_5959 ) ) ;
    buf_clk cell_3601 ( .C ( clk ), .D ( signal_1755 ), .Q ( signal_5961 ) ) ;
    buf_clk cell_3603 ( .C ( clk ), .D ( signal_3213 ), .Q ( signal_5963 ) ) ;
    buf_clk cell_3605 ( .C ( clk ), .D ( signal_1987 ), .Q ( signal_5965 ) ) ;
    buf_clk cell_3607 ( .C ( clk ), .D ( signal_3445 ), .Q ( signal_5967 ) ) ;
    buf_clk cell_3611 ( .C ( clk ), .D ( signal_5970 ), .Q ( signal_5971 ) ) ;
    buf_clk cell_3615 ( .C ( clk ), .D ( signal_5974 ), .Q ( signal_5975 ) ) ;
    buf_clk cell_3619 ( .C ( clk ), .D ( signal_5978 ), .Q ( signal_5979 ) ) ;
    buf_clk cell_3623 ( .C ( clk ), .D ( signal_5982 ), .Q ( signal_5983 ) ) ;
    buf_clk cell_3627 ( .C ( clk ), .D ( signal_5986 ), .Q ( signal_5987 ) ) ;
    buf_clk cell_3631 ( .C ( clk ), .D ( signal_5990 ), .Q ( signal_5991 ) ) ;
    buf_clk cell_3633 ( .C ( clk ), .D ( signal_5600 ), .Q ( signal_5993 ) ) ;
    buf_clk cell_3635 ( .C ( clk ), .D ( signal_5604 ), .Q ( signal_5995 ) ) ;
    buf_clk cell_3641 ( .C ( clk ), .D ( signal_6000 ), .Q ( signal_6001 ) ) ;
    buf_clk cell_3647 ( .C ( clk ), .D ( signal_6006 ), .Q ( signal_6007 ) ) ;
    buf_clk cell_3651 ( .C ( clk ), .D ( signal_6010 ), .Q ( signal_6011 ) ) ;
    buf_clk cell_3655 ( .C ( clk ), .D ( signal_6014 ), .Q ( signal_6015 ) ) ;
    buf_clk cell_3661 ( .C ( clk ), .D ( signal_6020 ), .Q ( signal_6021 ) ) ;
    buf_clk cell_3667 ( .C ( clk ), .D ( signal_6026 ), .Q ( signal_6027 ) ) ;
    buf_clk cell_3671 ( .C ( clk ), .D ( signal_6030 ), .Q ( signal_6031 ) ) ;
    buf_clk cell_3675 ( .C ( clk ), .D ( signal_6034 ), .Q ( signal_6035 ) ) ;
    buf_clk cell_3679 ( .C ( clk ), .D ( signal_6038 ), .Q ( signal_6039 ) ) ;
    buf_clk cell_3683 ( .C ( clk ), .D ( signal_6042 ), .Q ( signal_6043 ) ) ;
    buf_clk cell_3687 ( .C ( clk ), .D ( signal_6046 ), .Q ( signal_6047 ) ) ;
    buf_clk cell_3691 ( .C ( clk ), .D ( signal_6050 ), .Q ( signal_6051 ) ) ;
    buf_clk cell_3693 ( .C ( clk ), .D ( signal_1966 ), .Q ( signal_6053 ) ) ;
    buf_clk cell_3695 ( .C ( clk ), .D ( signal_3424 ), .Q ( signal_6055 ) ) ;
    buf_clk cell_3699 ( .C ( clk ), .D ( signal_6058 ), .Q ( signal_6059 ) ) ;
    buf_clk cell_3703 ( .C ( clk ), .D ( signal_6062 ), .Q ( signal_6063 ) ) ;
    buf_clk cell_3707 ( .C ( clk ), .D ( signal_6066 ), .Q ( signal_6067 ) ) ;
    buf_clk cell_3711 ( .C ( clk ), .D ( signal_6070 ), .Q ( signal_6071 ) ) ;
    buf_clk cell_3717 ( .C ( clk ), .D ( signal_6076 ), .Q ( signal_6077 ) ) ;
    buf_clk cell_3723 ( .C ( clk ), .D ( signal_6082 ), .Q ( signal_6083 ) ) ;
    buf_clk cell_3725 ( .C ( clk ), .D ( signal_2011 ), .Q ( signal_6085 ) ) ;
    buf_clk cell_3727 ( .C ( clk ), .D ( signal_3469 ), .Q ( signal_6087 ) ) ;
    buf_clk cell_3729 ( .C ( clk ), .D ( signal_1843 ), .Q ( signal_6089 ) ) ;
    buf_clk cell_3731 ( .C ( clk ), .D ( signal_3301 ), .Q ( signal_6091 ) ) ;
    buf_clk cell_3735 ( .C ( clk ), .D ( signal_6094 ), .Q ( signal_6095 ) ) ;
    buf_clk cell_3739 ( .C ( clk ), .D ( signal_6098 ), .Q ( signal_6099 ) ) ;
    buf_clk cell_3745 ( .C ( clk ), .D ( signal_6104 ), .Q ( signal_6105 ) ) ;
    buf_clk cell_3751 ( .C ( clk ), .D ( signal_6110 ), .Q ( signal_6111 ) ) ;
    buf_clk cell_3757 ( .C ( clk ), .D ( signal_6116 ), .Q ( signal_6117 ) ) ;
    buf_clk cell_3763 ( .C ( clk ), .D ( signal_6122 ), .Q ( signal_6123 ) ) ;
    buf_clk cell_3769 ( .C ( clk ), .D ( signal_6128 ), .Q ( signal_6129 ) ) ;
    buf_clk cell_3775 ( .C ( clk ), .D ( signal_6134 ), .Q ( signal_6135 ) ) ;
    buf_clk cell_3779 ( .C ( clk ), .D ( signal_6138 ), .Q ( signal_6139 ) ) ;
    buf_clk cell_3783 ( .C ( clk ), .D ( signal_6142 ), .Q ( signal_6143 ) ) ;
    buf_clk cell_3785 ( .C ( clk ), .D ( signal_5592 ), .Q ( signal_6145 ) ) ;
    buf_clk cell_3787 ( .C ( clk ), .D ( signal_5596 ), .Q ( signal_6147 ) ) ;
    buf_clk cell_3789 ( .C ( clk ), .D ( signal_5612 ), .Q ( signal_6149 ) ) ;
    buf_clk cell_3791 ( .C ( clk ), .D ( signal_5616 ), .Q ( signal_6151 ) ) ;
    buf_clk cell_3797 ( .C ( clk ), .D ( signal_6156 ), .Q ( signal_6157 ) ) ;
    buf_clk cell_3805 ( .C ( clk ), .D ( signal_6164 ), .Q ( signal_6165 ) ) ;
    buf_clk cell_3809 ( .C ( clk ), .D ( signal_1758 ), .Q ( signal_6169 ) ) ;
    buf_clk cell_3813 ( .C ( clk ), .D ( signal_3216 ), .Q ( signal_6173 ) ) ;
    buf_clk cell_3819 ( .C ( clk ), .D ( signal_6178 ), .Q ( signal_6179 ) ) ;
    buf_clk cell_3825 ( .C ( clk ), .D ( signal_6184 ), .Q ( signal_6185 ) ) ;
    buf_clk cell_3831 ( .C ( clk ), .D ( signal_6190 ), .Q ( signal_6191 ) ) ;
    buf_clk cell_3837 ( .C ( clk ), .D ( signal_6196 ), .Q ( signal_6197 ) ) ;
    buf_clk cell_3841 ( .C ( clk ), .D ( signal_1762 ), .Q ( signal_6201 ) ) ;
    buf_clk cell_3845 ( .C ( clk ), .D ( signal_3220 ), .Q ( signal_6205 ) ) ;
    buf_clk cell_3851 ( .C ( clk ), .D ( signal_6210 ), .Q ( signal_6211 ) ) ;
    buf_clk cell_3857 ( .C ( clk ), .D ( signal_6216 ), .Q ( signal_6217 ) ) ;
    buf_clk cell_3861 ( .C ( clk ), .D ( signal_5532 ), .Q ( signal_6221 ) ) ;
    buf_clk cell_3865 ( .C ( clk ), .D ( signal_5536 ), .Q ( signal_6225 ) ) ;
    buf_clk cell_3869 ( .C ( clk ), .D ( signal_1845 ), .Q ( signal_6229 ) ) ;
    buf_clk cell_3873 ( .C ( clk ), .D ( signal_3303 ), .Q ( signal_6233 ) ) ;
    buf_clk cell_3887 ( .C ( clk ), .D ( signal_6246 ), .Q ( signal_6247 ) ) ;
    buf_clk cell_3893 ( .C ( clk ), .D ( signal_6252 ), .Q ( signal_6253 ) ) ;
    buf_clk cell_3899 ( .C ( clk ), .D ( signal_6258 ), .Q ( signal_6259 ) ) ;
    buf_clk cell_3905 ( .C ( clk ), .D ( signal_6264 ), .Q ( signal_6265 ) ) ;
    buf_clk cell_3911 ( .C ( clk ), .D ( signal_6270 ), .Q ( signal_6271 ) ) ;
    buf_clk cell_3917 ( .C ( clk ), .D ( signal_6276 ), .Q ( signal_6277 ) ) ;
    buf_clk cell_3925 ( .C ( clk ), .D ( signal_1810 ), .Q ( signal_6285 ) ) ;
    buf_clk cell_3929 ( .C ( clk ), .D ( signal_3268 ), .Q ( signal_6289 ) ) ;
    buf_clk cell_3935 ( .C ( clk ), .D ( signal_6294 ), .Q ( signal_6295 ) ) ;
    buf_clk cell_3941 ( .C ( clk ), .D ( signal_6300 ), .Q ( signal_6301 ) ) ;
    buf_clk cell_3951 ( .C ( clk ), .D ( signal_6310 ), .Q ( signal_6311 ) ) ;
    buf_clk cell_3957 ( .C ( clk ), .D ( signal_6316 ), .Q ( signal_6317 ) ) ;
    buf_clk cell_3969 ( .C ( clk ), .D ( signal_6328 ), .Q ( signal_6329 ) ) ;
    buf_clk cell_3977 ( .C ( clk ), .D ( signal_6336 ), .Q ( signal_6337 ) ) ;
    buf_clk cell_3981 ( .C ( clk ), .D ( signal_1814 ), .Q ( signal_6341 ) ) ;
    buf_clk cell_3985 ( .C ( clk ), .D ( signal_3272 ), .Q ( signal_6345 ) ) ;
    buf_clk cell_3989 ( .C ( clk ), .D ( signal_1820 ), .Q ( signal_6349 ) ) ;
    buf_clk cell_3993 ( .C ( clk ), .D ( signal_3278 ), .Q ( signal_6353 ) ) ;
    buf_clk cell_3999 ( .C ( clk ), .D ( signal_6358 ), .Q ( signal_6359 ) ) ;
    buf_clk cell_4005 ( .C ( clk ), .D ( signal_6364 ), .Q ( signal_6365 ) ) ;
    buf_clk cell_4011 ( .C ( clk ), .D ( signal_6370 ), .Q ( signal_6371 ) ) ;
    buf_clk cell_4017 ( .C ( clk ), .D ( signal_6376 ), .Q ( signal_6377 ) ) ;
    buf_clk cell_4021 ( .C ( clk ), .D ( signal_2006 ), .Q ( signal_6381 ) ) ;
    buf_clk cell_4025 ( .C ( clk ), .D ( signal_3464 ), .Q ( signal_6385 ) ) ;
    buf_clk cell_4033 ( .C ( clk ), .D ( signal_6392 ), .Q ( signal_6393 ) ) ;
    buf_clk cell_4041 ( .C ( clk ), .D ( signal_6400 ), .Q ( signal_6401 ) ) ;
    buf_clk cell_4047 ( .C ( clk ), .D ( signal_6406 ), .Q ( signal_6407 ) ) ;
    buf_clk cell_4053 ( .C ( clk ), .D ( signal_6412 ), .Q ( signal_6413 ) ) ;
    buf_clk cell_4059 ( .C ( clk ), .D ( signal_6418 ), .Q ( signal_6419 ) ) ;
    buf_clk cell_4065 ( .C ( clk ), .D ( signal_6424 ), .Q ( signal_6425 ) ) ;
    buf_clk cell_4079 ( .C ( clk ), .D ( signal_6438 ), .Q ( signal_6439 ) ) ;
    buf_clk cell_4085 ( .C ( clk ), .D ( signal_6444 ), .Q ( signal_6445 ) ) ;
    buf_clk cell_4099 ( .C ( clk ), .D ( signal_6458 ), .Q ( signal_6459 ) ) ;
    buf_clk cell_4105 ( .C ( clk ), .D ( signal_6464 ), .Q ( signal_6465 ) ) ;
    buf_clk cell_4111 ( .C ( clk ), .D ( signal_6470 ), .Q ( signal_6471 ) ) ;
    buf_clk cell_4117 ( .C ( clk ), .D ( signal_6476 ), .Q ( signal_6477 ) ) ;
    buf_clk cell_4121 ( .C ( clk ), .D ( signal_1818 ), .Q ( signal_6481 ) ) ;
    buf_clk cell_4125 ( .C ( clk ), .D ( signal_3276 ), .Q ( signal_6485 ) ) ;
    buf_clk cell_4133 ( .C ( clk ), .D ( signal_6492 ), .Q ( signal_6493 ) ) ;
    buf_clk cell_4143 ( .C ( clk ), .D ( signal_6502 ), .Q ( signal_6503 ) ) ;
    buf_clk cell_4149 ( .C ( clk ), .D ( signal_1988 ), .Q ( signal_6509 ) ) ;
    buf_clk cell_4155 ( .C ( clk ), .D ( signal_3446 ), .Q ( signal_6515 ) ) ;
    buf_clk cell_4163 ( .C ( clk ), .D ( signal_6522 ), .Q ( signal_6523 ) ) ;
    buf_clk cell_4171 ( .C ( clk ), .D ( signal_6530 ), .Q ( signal_6531 ) ) ;
    buf_clk cell_4179 ( .C ( clk ), .D ( signal_6538 ), .Q ( signal_6539 ) ) ;
    buf_clk cell_4187 ( .C ( clk ), .D ( signal_6546 ), .Q ( signal_6547 ) ) ;
    buf_clk cell_4229 ( .C ( clk ), .D ( signal_6588 ), .Q ( signal_6589 ) ) ;
    buf_clk cell_4239 ( .C ( clk ), .D ( signal_6598 ), .Q ( signal_6599 ) ) ;
    buf_clk cell_4245 ( .C ( clk ), .D ( signal_2016 ), .Q ( signal_6605 ) ) ;
    buf_clk cell_4251 ( .C ( clk ), .D ( signal_3474 ), .Q ( signal_6611 ) ) ;
    buf_clk cell_4263 ( .C ( clk ), .D ( signal_6622 ), .Q ( signal_6623 ) ) ;
    buf_clk cell_4271 ( .C ( clk ), .D ( signal_6630 ), .Q ( signal_6631 ) ) ;
    buf_clk cell_4277 ( .C ( clk ), .D ( signal_1979 ), .Q ( signal_6637 ) ) ;
    buf_clk cell_4283 ( .C ( clk ), .D ( signal_3437 ), .Q ( signal_6643 ) ) ;
    buf_clk cell_4291 ( .C ( clk ), .D ( signal_6650 ), .Q ( signal_6651 ) ) ;
    buf_clk cell_4299 ( .C ( clk ), .D ( signal_6658 ), .Q ( signal_6659 ) ) ;
    buf_clk cell_4307 ( .C ( clk ), .D ( signal_6666 ), .Q ( signal_6667 ) ) ;
    buf_clk cell_4315 ( .C ( clk ), .D ( signal_6674 ), .Q ( signal_6675 ) ) ;
    buf_clk cell_4323 ( .C ( clk ), .D ( signal_6682 ), .Q ( signal_6683 ) ) ;
    buf_clk cell_4331 ( .C ( clk ), .D ( signal_6690 ), .Q ( signal_6691 ) ) ;
    buf_clk cell_4341 ( .C ( clk ), .D ( signal_6700 ), .Q ( signal_6701 ) ) ;
    buf_clk cell_4351 ( .C ( clk ), .D ( signal_6710 ), .Q ( signal_6711 ) ) ;
    buf_clk cell_4359 ( .C ( clk ), .D ( signal_6718 ), .Q ( signal_6719 ) ) ;
    buf_clk cell_4367 ( .C ( clk ), .D ( signal_6726 ), .Q ( signal_6727 ) ) ;
    buf_clk cell_4375 ( .C ( clk ), .D ( signal_6734 ), .Q ( signal_6735 ) ) ;
    buf_clk cell_4383 ( .C ( clk ), .D ( signal_6742 ), .Q ( signal_6743 ) ) ;
    buf_clk cell_4395 ( .C ( clk ), .D ( signal_6754 ), .Q ( signal_6755 ) ) ;
    buf_clk cell_4403 ( .C ( clk ), .D ( signal_6762 ), .Q ( signal_6763 ) ) ;
    buf_clk cell_4411 ( .C ( clk ), .D ( signal_6770 ), .Q ( signal_6771 ) ) ;
    buf_clk cell_4419 ( .C ( clk ), .D ( signal_6778 ), .Q ( signal_6779 ) ) ;
    buf_clk cell_4427 ( .C ( clk ), .D ( signal_6786 ), .Q ( signal_6787 ) ) ;
    buf_clk cell_4435 ( .C ( clk ), .D ( signal_6794 ), .Q ( signal_6795 ) ) ;
    buf_clk cell_4453 ( .C ( clk ), .D ( signal_2030 ), .Q ( signal_6813 ) ) ;
    buf_clk cell_4461 ( .C ( clk ), .D ( signal_3488 ), .Q ( signal_6821 ) ) ;
    buf_clk cell_4493 ( .C ( clk ), .D ( signal_5738 ), .Q ( signal_6853 ) ) ;
    buf_clk cell_4501 ( .C ( clk ), .D ( signal_5740 ), .Q ( signal_6861 ) ) ;
    buf_clk cell_4511 ( .C ( clk ), .D ( signal_6870 ), .Q ( signal_6871 ) ) ;
    buf_clk cell_4521 ( .C ( clk ), .D ( signal_6880 ), .Q ( signal_6881 ) ) ;
    buf_clk cell_4545 ( .C ( clk ), .D ( signal_1982 ), .Q ( signal_6905 ) ) ;
    buf_clk cell_4553 ( .C ( clk ), .D ( signal_3440 ), .Q ( signal_6913 ) ) ;
    buf_clk cell_4563 ( .C ( clk ), .D ( signal_6922 ), .Q ( signal_6923 ) ) ;
    buf_clk cell_4573 ( .C ( clk ), .D ( signal_6932 ), .Q ( signal_6933 ) ) ;
    buf_clk cell_4581 ( .C ( clk ), .D ( signal_1967 ), .Q ( signal_6941 ) ) ;
    buf_clk cell_4589 ( .C ( clk ), .D ( signal_3425 ), .Q ( signal_6949 ) ) ;
    buf_clk cell_4741 ( .C ( clk ), .D ( signal_1978 ), .Q ( signal_7101 ) ) ;
    buf_clk cell_4751 ( .C ( clk ), .D ( signal_3436 ), .Q ( signal_7111 ) ) ;
    buf_clk cell_4917 ( .C ( clk ), .D ( signal_1736 ), .Q ( signal_7277 ) ) ;
    buf_clk cell_4929 ( .C ( clk ), .D ( signal_3194 ), .Q ( signal_7289 ) ) ;
    buf_clk cell_4967 ( .C ( clk ), .D ( signal_7326 ), .Q ( signal_7327 ) ) ;
    buf_clk cell_4981 ( .C ( clk ), .D ( signal_7340 ), .Q ( signal_7341 ) ) ;
    buf_clk cell_5011 ( .C ( clk ), .D ( signal_7370 ), .Q ( signal_7371 ) ) ;
    buf_clk cell_5025 ( .C ( clk ), .D ( signal_7384 ), .Q ( signal_7385 ) ) ;
    buf_clk cell_5091 ( .C ( clk ), .D ( signal_7450 ), .Q ( signal_7451 ) ) ;
    buf_clk cell_5107 ( .C ( clk ), .D ( signal_7466 ), .Q ( signal_7467 ) ) ;
    buf_clk cell_5131 ( .C ( clk ), .D ( signal_7490 ), .Q ( signal_7491 ) ) ;
    buf_clk cell_5147 ( .C ( clk ), .D ( signal_7506 ), .Q ( signal_7507 ) ) ;
    buf_clk cell_5253 ( .C ( clk ), .D ( signal_1783 ), .Q ( signal_7613 ) ) ;
    buf_clk cell_5269 ( .C ( clk ), .D ( signal_3241 ), .Q ( signal_7629 ) ) ;
    buf_clk cell_5287 ( .C ( clk ), .D ( signal_7646 ), .Q ( signal_7647 ) ) ;
    buf_clk cell_5305 ( .C ( clk ), .D ( signal_7664 ), .Q ( signal_7665 ) ) ;
    buf_clk cell_5387 ( .C ( clk ), .D ( signal_7746 ), .Q ( signal_7747 ) ) ;
    buf_clk cell_5407 ( .C ( clk ), .D ( signal_7766 ), .Q ( signal_7767 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1819 ( .a ({signal_5380, signal_5378}), .b ({signal_3145, signal_1687}), .clk ( clk ), .r ( Fresh[581] ), .c ({signal_3292, signal_1834}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1834 ( .a ({signal_5384, signal_5382}), .b ({signal_3168, signal_1710}), .clk ( clk ), .r ( Fresh[582] ), .c ({signal_3307, signal_1849}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1872 ( .a ({signal_3292, signal_1834}), .b ({signal_3345, signal_1887}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1875 ( .a ({signal_3307, signal_1849}), .b ({signal_3348, signal_1890}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1893 ( .a ({signal_5392, signal_5388}), .b ({signal_3188, signal_1730}), .clk ( clk ), .r ( Fresh[583] ), .c ({signal_3366, signal_1908}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1902 ( .a ({signal_3225, signal_1767}), .b ({signal_3244, signal_1786}), .clk ( clk ), .r ( Fresh[584] ), .c ({signal_3375, signal_1917}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1904 ( .a ({signal_5392, signal_5388}), .b ({signal_3198, signal_1740}), .clk ( clk ), .r ( Fresh[585] ), .c ({signal_3377, signal_1919}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1911 ( .a ({signal_3248, signal_1790}), .b ({signal_5396, signal_5394}), .clk ( clk ), .r ( Fresh[586] ), .c ({signal_3384, signal_1926}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1912 ( .a ({signal_5404, signal_5400}), .b ({signal_3250, signal_1792}), .clk ( clk ), .r ( Fresh[587] ), .c ({signal_3385, signal_1927}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1918 ( .a ({signal_5412, signal_5408}), .b ({signal_3262, signal_1804}), .clk ( clk ), .r ( Fresh[588] ), .c ({signal_3391, signal_1933}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1921 ( .a ({signal_5420, signal_5416}), .b ({signal_3264, signal_1806}), .clk ( clk ), .r ( Fresh[589] ), .c ({signal_3394, signal_1936}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1922 ( .a ({signal_3266, signal_1808}), .b ({signal_3267, signal_1809}), .clk ( clk ), .r ( Fresh[590] ), .c ({signal_3395, signal_1937}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1924 ( .a ({signal_5436, signal_5428}), .b ({signal_3210, signal_1752}), .clk ( clk ), .r ( Fresh[591] ), .c ({signal_3397, signal_1939}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1925 ( .a ({signal_5440, signal_5438}), .b ({signal_3273, signal_1815}), .clk ( clk ), .r ( Fresh[592] ), .c ({signal_3398, signal_1940}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1926 ( .a ({signal_5444, signal_5442}), .b ({signal_3211, signal_1753}), .clk ( clk ), .r ( Fresh[593] ), .c ({signal_3399, signal_1941}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1928 ( .a ({signal_5452, signal_5448}), .b ({signal_3277, signal_1819}), .clk ( clk ), .r ( Fresh[594] ), .c ({signal_3401, signal_1943}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1929 ( .a ({signal_3247, signal_1789}), .b ({signal_5456, signal_5454}), .clk ( clk ), .r ( Fresh[595] ), .c ({signal_3402, signal_1944}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1930 ( .a ({signal_3214, signal_1756}), .b ({signal_3215, signal_1757}), .clk ( clk ), .r ( Fresh[596] ), .c ({signal_3403, signal_1945}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1931 ( .a ({signal_5460, signal_5458}), .b ({signal_3217, signal_1759}), .clk ( clk ), .r ( Fresh[597] ), .c ({signal_3404, signal_1946}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1933 ( .a ({signal_5468, signal_5464}), .b ({signal_3285, signal_1827}), .clk ( clk ), .r ( Fresh[598] ), .c ({signal_3406, signal_1948}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1934 ( .a ({signal_5472, signal_5470}), .b ({signal_3291, signal_1833}), .clk ( clk ), .r ( Fresh[599] ), .c ({signal_3407, signal_1949}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1935 ( .a ({signal_5476, signal_5474}), .b ({signal_3293, signal_1835}), .clk ( clk ), .r ( Fresh[600] ), .c ({signal_3408, signal_1950}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1936 ( .a ({signal_3219, signal_1761}), .b ({signal_3294, signal_1836}), .clk ( clk ), .r ( Fresh[601] ), .c ({signal_3409, signal_1951}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1937 ( .a ({signal_5480, signal_5478}), .b ({signal_3213, signal_1755}), .clk ( clk ), .r ( Fresh[602] ), .c ({signal_3410, signal_1952}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1938 ( .a ({signal_5484, signal_5482}), .b ({signal_3295, signal_1837}), .clk ( clk ), .r ( Fresh[603] ), .c ({signal_3411, signal_1953}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1939 ( .a ({signal_5488, signal_5486}), .b ({signal_3296, signal_1838}), .clk ( clk ), .r ( Fresh[604] ), .c ({signal_3412, signal_1954}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1940 ( .a ({signal_5496, signal_5492}), .b ({signal_3298, signal_1840}), .clk ( clk ), .r ( Fresh[605] ), .c ({signal_3413, signal_1955}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1941 ( .a ({signal_5500, signal_5498}), .b ({signal_3221, signal_1763}), .clk ( clk ), .r ( Fresh[606] ), .c ({signal_3414, signal_1956}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1942 ( .a ({signal_5504, signal_5502}), .b ({signal_3299, signal_1841}), .clk ( clk ), .r ( Fresh[607] ), .c ({signal_3415, signal_1957}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1943 ( .a ({signal_3261, signal_1803}), .b ({signal_5508, signal_5506}), .clk ( clk ), .r ( Fresh[608] ), .c ({signal_3416, signal_1958}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1945 ( .a ({signal_3283, signal_1825}), .b ({signal_3304, signal_1846}), .clk ( clk ), .r ( Fresh[609] ), .c ({signal_3418, signal_1960}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1946 ( .a ({signal_5512, signal_5510}), .b ({signal_3223, signal_1765}), .clk ( clk ), .r ( Fresh[610] ), .c ({signal_3419, signal_1961}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1947 ( .a ({signal_3254, signal_1796}), .b ({signal_3305, signal_1847}), .clk ( clk ), .r ( Fresh[611] ), .c ({signal_3420, signal_1962}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1961 ( .a ({signal_3366, signal_1908}), .b ({signal_3434, signal_1976}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1969 ( .a ({signal_3375, signal_1917}), .b ({signal_3442, signal_1984}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1971 ( .a ({signal_3377, signal_1919}), .b ({signal_3444, signal_1986}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1978 ( .a ({signal_3385, signal_1927}), .b ({signal_3451, signal_1993}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1986 ( .a ({signal_3394, signal_1936}), .b ({signal_3459, signal_2001}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1987 ( .a ({signal_3395, signal_1937}), .b ({signal_3460, signal_2002}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1989 ( .a ({signal_3397, signal_1939}), .b ({signal_3462, signal_2004}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1992 ( .a ({signal_3407, signal_1949}), .b ({signal_3465, signal_2007}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1993 ( .a ({signal_3409, signal_1951}), .b ({signal_3466, signal_2008}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1994 ( .a ({signal_3415, signal_1957}), .b ({signal_3467, signal_2009}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1995 ( .a ({signal_3416, signal_1958}), .b ({signal_3468, signal_2010}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1997 ( .a ({signal_3418, signal_1960}), .b ({signal_3470, signal_2012}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_1998 ( .a ({signal_3420, signal_1962}), .b ({signal_3471, signal_2013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_1999 ( .a ({signal_3315, signal_1857}), .b ({signal_5520, signal_5516}), .clk ( clk ), .r ( Fresh[612] ), .c ({signal_3472, signal_2014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2002 ( .a ({signal_5524, signal_5522}), .b ({signal_3232, signal_1774}), .clk ( clk ), .r ( Fresh[613] ), .c ({signal_3475, signal_2017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2007 ( .a ({signal_5528, signal_5526}), .b ({signal_3352, signal_1894}), .clk ( clk ), .r ( Fresh[614] ), .c ({signal_3480, signal_2022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2009 ( .a ({signal_5536, signal_5532}), .b ({signal_3354, signal_1896}), .clk ( clk ), .r ( Fresh[615] ), .c ({signal_3482, signal_2024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2010 ( .a ({signal_5544, signal_5540}), .b ({signal_3357, signal_1899}), .clk ( clk ), .r ( Fresh[616] ), .c ({signal_3483, signal_2025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2013 ( .a ({signal_5552, signal_5548}), .b ({signal_3326, signal_1868}), .clk ( clk ), .r ( Fresh[617] ), .c ({signal_3486, signal_2028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2016 ( .a ({signal_5560, signal_5556}), .b ({signal_3332, signal_1874}), .clk ( clk ), .r ( Fresh[618] ), .c ({signal_3489, signal_2031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2017 ( .a ({signal_5564, signal_5562}), .b ({signal_3333, signal_1875}), .clk ( clk ), .r ( Fresh[619] ), .c ({signal_3490, signal_2032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2018 ( .a ({signal_5568, signal_5566}), .b ({signal_3334, signal_1876}), .clk ( clk ), .r ( Fresh[620] ), .c ({signal_3491, signal_2033}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2019 ( .a ({signal_5572, signal_5570}), .b ({signal_3271, signal_1813}), .clk ( clk ), .r ( Fresh[621] ), .c ({signal_3492, signal_2034}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2020 ( .a ({signal_5576, signal_5574}), .b ({signal_3335, signal_1877}), .clk ( clk ), .r ( Fresh[622] ), .c ({signal_3493, signal_2035}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2021 ( .a ({signal_5580, signal_5578}), .b ({signal_3336, signal_1878}), .clk ( clk ), .r ( Fresh[623] ), .c ({signal_3494, signal_2036}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2022 ( .a ({signal_5588, signal_5584}), .b ({signal_3337, signal_1879}), .clk ( clk ), .r ( Fresh[624] ), .c ({signal_3495, signal_2037}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2023 ( .a ({signal_5596, signal_5592}), .b ({signal_3338, signal_1880}), .clk ( clk ), .r ( Fresh[625] ), .c ({signal_3496, signal_2038}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2024 ( .a ({signal_5604, signal_5600}), .b ({signal_3339, signal_1881}), .clk ( clk ), .r ( Fresh[626] ), .c ({signal_3497, signal_2039}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2025 ( .a ({signal_5608, signal_5606}), .b ({signal_3340, signal_1882}), .clk ( clk ), .r ( Fresh[627] ), .c ({signal_3498, signal_2040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2026 ( .a ({signal_3284, signal_1826}), .b ({signal_3374, signal_1916}), .clk ( clk ), .r ( Fresh[628] ), .c ({signal_3499, signal_2041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2028 ( .a ({signal_5616, signal_5612}), .b ({signal_3341, signal_1883}), .clk ( clk ), .r ( Fresh[629] ), .c ({signal_3501, signal_2043}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2029 ( .a ({signal_5620, signal_5618}), .b ({signal_3342, signal_1884}), .clk ( clk ), .r ( Fresh[630] ), .c ({signal_3502, signal_2044}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2030 ( .a ({signal_5624, signal_5622}), .b ({signal_3288, signal_1830}), .clk ( clk ), .r ( Fresh[631] ), .c ({signal_3503, signal_2045}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2031 ( .a ({signal_5628, signal_5626}), .b ({signal_3344, signal_1886}), .clk ( clk ), .r ( Fresh[632] ), .c ({signal_3504, signal_2046}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2033 ( .a ({signal_5632, signal_5630}), .b ({signal_3297, signal_1839}), .clk ( clk ), .r ( Fresh[633] ), .c ({signal_3506, signal_2048}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2034 ( .a ({signal_5636, signal_5634}), .b ({signal_3276, signal_1818}), .clk ( clk ), .r ( Fresh[634] ), .c ({signal_3507, signal_2049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2035 ( .a ({signal_5644, signal_5640}), .b ({signal_3346, signal_1888}), .clk ( clk ), .r ( Fresh[635] ), .c ({signal_3508, signal_2050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2036 ( .a ({signal_5536, signal_5532}), .b ({signal_3347, signal_1889}), .clk ( clk ), .r ( Fresh[636] ), .c ({signal_3509, signal_2051}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2046 ( .a ({signal_3472, signal_2014}), .b ({signal_3519, signal_2061}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2047 ( .a ({signal_3475, signal_2017}), .b ({signal_3520, signal_2062}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2049 ( .a ({signal_3480, signal_2022}), .b ({signal_3522, signal_2064}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2050 ( .a ({signal_3482, signal_2024}), .b ({signal_3523, signal_2065}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2051 ( .a ({signal_3483, signal_2025}), .b ({signal_3524, signal_2066}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2053 ( .a ({signal_3486, signal_2028}), .b ({signal_3526, signal_2068}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2054 ( .a ({signal_3489, signal_2031}), .b ({signal_3527, signal_2069}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2055 ( .a ({signal_3490, signal_2032}), .b ({signal_3528, signal_2070}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2056 ( .a ({signal_3491, signal_2033}), .b ({signal_3529, signal_2071}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2057 ( .a ({signal_3492, signal_2034}), .b ({signal_3530, signal_2072}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2058 ( .a ({signal_3493, signal_2035}), .b ({signal_3531, signal_2073}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2059 ( .a ({signal_3494, signal_2036}), .b ({signal_3532, signal_2074}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2060 ( .a ({signal_3495, signal_2037}), .b ({signal_3533, signal_2075}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2061 ( .a ({signal_3496, signal_2038}), .b ({signal_3534, signal_2076}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2062 ( .a ({signal_3497, signal_2039}), .b ({signal_3535, signal_2077}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2063 ( .a ({signal_3499, signal_2041}), .b ({signal_3536, signal_2078}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2065 ( .a ({signal_3501, signal_2043}), .b ({signal_3538, signal_2080}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2066 ( .a ({signal_3502, signal_2044}), .b ({signal_3539, signal_2081}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2067 ( .a ({signal_3504, signal_2046}), .b ({signal_3540, signal_2082}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2069 ( .a ({signal_3506, signal_2048}), .b ({signal_3542, signal_2084}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2070 ( .a ({signal_3508, signal_2050}), .b ({signal_3543, signal_2085}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2071 ( .a ({signal_3509, signal_2051}), .b ({signal_3544, signal_2086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2074 ( .a ({signal_3435, signal_1977}), .b ({signal_5652, signal_5648}), .clk ( clk ), .r ( Fresh[637] ), .c ({signal_3547, signal_2089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2075 ( .a ({signal_5656, signal_5654}), .b ({signal_3422, signal_1964}), .clk ( clk ), .r ( Fresh[638] ), .c ({signal_3548, signal_2090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2076 ( .a ({signal_5664, signal_5660}), .b ({signal_3473, signal_2015}), .clk ( clk ), .r ( Fresh[639] ), .c ({signal_3549, signal_2091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2077 ( .a ({signal_5668, signal_5666}), .b ({signal_3427, signal_1969}), .clk ( clk ), .r ( Fresh[640] ), .c ({signal_3550, signal_2092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2078 ( .a ({signal_3421, signal_1963}), .b ({signal_5672, signal_5670}), .clk ( clk ), .r ( Fresh[641] ), .c ({signal_3551, signal_2093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2079 ( .a ({signal_3431, signal_1973}), .b ({signal_3432, signal_1974}), .clk ( clk ), .r ( Fresh[642] ), .c ({signal_3552, signal_2094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2080 ( .a ({signal_5680, signal_5676}), .b ({signal_3476, signal_2018}), .clk ( clk ), .r ( Fresh[643] ), .c ({signal_3553, signal_2095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2081 ( .a ({signal_5688, signal_5684}), .b ({signal_3478, signal_2020}), .clk ( clk ), .r ( Fresh[644] ), .c ({signal_3554, signal_2096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2082 ( .a ({signal_5696, signal_5692}), .b ({signal_3479, signal_2021}), .clk ( clk ), .r ( Fresh[645] ), .c ({signal_3555, signal_2097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2083 ( .a ({signal_5700, signal_5698}), .b ({signal_3439, signal_1981}), .clk ( clk ), .r ( Fresh[646] ), .c ({signal_3556, signal_2098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2085 ( .a ({signal_5708, signal_5704}), .b ({signal_3443, signal_1985}), .clk ( clk ), .r ( Fresh[647] ), .c ({signal_3558, signal_2100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2086 ( .a ({signal_5716, signal_5712}), .b ({signal_3481, signal_2023}), .clk ( clk ), .r ( Fresh[648] ), .c ({signal_3559, signal_2101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2087 ( .a ({signal_3349, signal_1891}), .b ({signal_3447, signal_1989}), .clk ( clk ), .r ( Fresh[649] ), .c ({signal_3560, signal_2102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2088 ( .a ({signal_3448, signal_1990}), .b ({signal_3449, signal_1991}), .clk ( clk ), .r ( Fresh[650] ), .c ({signal_3561, signal_2103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2089 ( .a ({signal_5720, signal_5718}), .b ({signal_3450, signal_1992}), .clk ( clk ), .r ( Fresh[651] ), .c ({signal_3562, signal_2104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2091 ( .a ({signal_3485, signal_2027}), .b ({signal_3343, signal_1885}), .clk ( clk ), .r ( Fresh[652] ), .c ({signal_3564, signal_2106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2092 ( .a ({signal_5728, signal_5724}), .b ({signal_3452, signal_1994}), .clk ( clk ), .r ( Fresh[653] ), .c ({signal_3565, signal_2107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2093 ( .a ({signal_5732, signal_5730}), .b ({signal_3453, signal_1995}), .clk ( clk ), .r ( Fresh[654] ), .c ({signal_3566, signal_2108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2094 ( .a ({signal_3260, signal_1802}), .b ({signal_3454, signal_1996}), .clk ( clk ), .r ( Fresh[655] ), .c ({signal_3567, signal_2109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2095 ( .a ({signal_3429, signal_1971}), .b ({signal_3455, signal_1997}), .clk ( clk ), .r ( Fresh[656] ), .c ({signal_3568, signal_2110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2096 ( .a ({signal_3214, signal_1756}), .b ({signal_3456, signal_1998}), .clk ( clk ), .r ( Fresh[657] ), .c ({signal_3569, signal_2111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2097 ( .a ({signal_3430, signal_1972}), .b ({signal_5456, signal_5454}), .clk ( clk ), .r ( Fresh[658] ), .c ({signal_3570, signal_2112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2099 ( .a ({signal_3156, signal_1698}), .b ({signal_3458, signal_2000}), .clk ( clk ), .r ( Fresh[659] ), .c ({signal_3572, signal_2114}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2101 ( .a ({signal_3433, signal_1975}), .b ({signal_3461, signal_2003}), .clk ( clk ), .r ( Fresh[660] ), .c ({signal_3574, signal_2116}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2104 ( .a ({signal_5736, signal_5734}), .b ({signal_3463, signal_2005}), .clk ( clk ), .r ( Fresh[661] ), .c ({signal_3577, signal_2119}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2110 ( .a ({signal_3487, signal_2029}), .b ({signal_3306, signal_1848}), .clk ( clk ), .r ( Fresh[662] ), .c ({signal_3583, signal_2125}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2124 ( .a ({signal_3547, signal_2089}), .b ({signal_3597, signal_2139}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2125 ( .a ({signal_3549, signal_2091}), .b ({signal_3598, signal_2140}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2126 ( .a ({signal_3550, signal_2092}), .b ({signal_3599, signal_2141}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2127 ( .a ({signal_3554, signal_2096}), .b ({signal_3600, signal_2142}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2128 ( .a ({signal_3555, signal_2097}), .b ({signal_3601, signal_2143}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2130 ( .a ({signal_3559, signal_2101}), .b ({signal_3603, signal_2145}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2133 ( .a ({signal_3577, signal_2119}), .b ({signal_3606, signal_2148}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2135 ( .a ({signal_3583, signal_2125}), .b ({signal_3608, signal_2150}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2144 ( .a ({signal_5740, signal_5738}), .b ({signal_3521, signal_2063}), .clk ( clk ), .r ( Fresh[663] ), .c ({signal_3617, signal_2159}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2148 ( .a ({signal_5748, signal_5744}), .b ({signal_3525, signal_2067}), .clk ( clk ), .r ( Fresh[664] ), .c ({signal_3621, signal_2163}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2185 ( .a ({signal_3617, signal_2159}), .b ({signal_3658, signal_2200}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2186 ( .a ({signal_3621, signal_2163}), .b ({signal_3659, signal_2201}) ) ;
    buf_clk cell_3390 ( .C ( clk ), .D ( signal_5749 ), .Q ( signal_5750 ) ) ;
    buf_clk cell_3392 ( .C ( clk ), .D ( signal_5751 ), .Q ( signal_5752 ) ) ;
    buf_clk cell_3398 ( .C ( clk ), .D ( signal_5757 ), .Q ( signal_5758 ) ) ;
    buf_clk cell_3404 ( .C ( clk ), .D ( signal_5763 ), .Q ( signal_5764 ) ) ;
    buf_clk cell_3410 ( .C ( clk ), .D ( signal_5769 ), .Q ( signal_5770 ) ) ;
    buf_clk cell_3416 ( .C ( clk ), .D ( signal_5775 ), .Q ( signal_5776 ) ) ;
    buf_clk cell_3422 ( .C ( clk ), .D ( signal_5781 ), .Q ( signal_5782 ) ) ;
    buf_clk cell_3428 ( .C ( clk ), .D ( signal_5787 ), .Q ( signal_5788 ) ) ;
    buf_clk cell_3432 ( .C ( clk ), .D ( signal_5791 ), .Q ( signal_5792 ) ) ;
    buf_clk cell_3436 ( .C ( clk ), .D ( signal_5795 ), .Q ( signal_5796 ) ) ;
    buf_clk cell_3442 ( .C ( clk ), .D ( signal_5801 ), .Q ( signal_5802 ) ) ;
    buf_clk cell_3448 ( .C ( clk ), .D ( signal_5807 ), .Q ( signal_5808 ) ) ;
    buf_clk cell_3452 ( .C ( clk ), .D ( signal_5811 ), .Q ( signal_5812 ) ) ;
    buf_clk cell_3456 ( .C ( clk ), .D ( signal_5815 ), .Q ( signal_5816 ) ) ;
    buf_clk cell_3460 ( .C ( clk ), .D ( signal_5819 ), .Q ( signal_5820 ) ) ;
    buf_clk cell_3464 ( .C ( clk ), .D ( signal_5823 ), .Q ( signal_5824 ) ) ;
    buf_clk cell_3468 ( .C ( clk ), .D ( signal_5827 ), .Q ( signal_5828 ) ) ;
    buf_clk cell_3472 ( .C ( clk ), .D ( signal_5831 ), .Q ( signal_5832 ) ) ;
    buf_clk cell_3476 ( .C ( clk ), .D ( signal_5835 ), .Q ( signal_5836 ) ) ;
    buf_clk cell_3480 ( .C ( clk ), .D ( signal_5839 ), .Q ( signal_5840 ) ) ;
    buf_clk cell_3484 ( .C ( clk ), .D ( signal_5843 ), .Q ( signal_5844 ) ) ;
    buf_clk cell_3488 ( .C ( clk ), .D ( signal_5847 ), .Q ( signal_5848 ) ) ;
    buf_clk cell_3494 ( .C ( clk ), .D ( signal_5853 ), .Q ( signal_5854 ) ) ;
    buf_clk cell_3500 ( .C ( clk ), .D ( signal_5859 ), .Q ( signal_5860 ) ) ;
    buf_clk cell_3504 ( .C ( clk ), .D ( signal_5863 ), .Q ( signal_5864 ) ) ;
    buf_clk cell_3508 ( .C ( clk ), .D ( signal_5867 ), .Q ( signal_5868 ) ) ;
    buf_clk cell_3510 ( .C ( clk ), .D ( signal_5869 ), .Q ( signal_5870 ) ) ;
    buf_clk cell_3512 ( .C ( clk ), .D ( signal_5871 ), .Q ( signal_5872 ) ) ;
    buf_clk cell_3514 ( .C ( clk ), .D ( signal_5873 ), .Q ( signal_5874 ) ) ;
    buf_clk cell_3516 ( .C ( clk ), .D ( signal_5875 ), .Q ( signal_5876 ) ) ;
    buf_clk cell_3518 ( .C ( clk ), .D ( signal_5877 ), .Q ( signal_5878 ) ) ;
    buf_clk cell_3520 ( .C ( clk ), .D ( signal_5879 ), .Q ( signal_5880 ) ) ;
    buf_clk cell_3522 ( .C ( clk ), .D ( signal_5881 ), .Q ( signal_5882 ) ) ;
    buf_clk cell_3524 ( .C ( clk ), .D ( signal_5883 ), .Q ( signal_5884 ) ) ;
    buf_clk cell_3526 ( .C ( clk ), .D ( signal_5885 ), .Q ( signal_5886 ) ) ;
    buf_clk cell_3528 ( .C ( clk ), .D ( signal_5887 ), .Q ( signal_5888 ) ) ;
    buf_clk cell_3532 ( .C ( clk ), .D ( signal_5891 ), .Q ( signal_5892 ) ) ;
    buf_clk cell_3536 ( .C ( clk ), .D ( signal_5895 ), .Q ( signal_5896 ) ) ;
    buf_clk cell_3538 ( .C ( clk ), .D ( signal_5897 ), .Q ( signal_5898 ) ) ;
    buf_clk cell_3540 ( .C ( clk ), .D ( signal_5899 ), .Q ( signal_5900 ) ) ;
    buf_clk cell_3542 ( .C ( clk ), .D ( signal_5901 ), .Q ( signal_5902 ) ) ;
    buf_clk cell_3544 ( .C ( clk ), .D ( signal_5903 ), .Q ( signal_5904 ) ) ;
    buf_clk cell_3546 ( .C ( clk ), .D ( signal_5905 ), .Q ( signal_5906 ) ) ;
    buf_clk cell_3548 ( .C ( clk ), .D ( signal_5907 ), .Q ( signal_5908 ) ) ;
    buf_clk cell_3554 ( .C ( clk ), .D ( signal_5913 ), .Q ( signal_5914 ) ) ;
    buf_clk cell_3560 ( .C ( clk ), .D ( signal_5919 ), .Q ( signal_5920 ) ) ;
    buf_clk cell_3562 ( .C ( clk ), .D ( signal_5921 ), .Q ( signal_5922 ) ) ;
    buf_clk cell_3564 ( .C ( clk ), .D ( signal_5923 ), .Q ( signal_5924 ) ) ;
    buf_clk cell_3568 ( .C ( clk ), .D ( signal_5927 ), .Q ( signal_5928 ) ) ;
    buf_clk cell_3572 ( .C ( clk ), .D ( signal_5931 ), .Q ( signal_5932 ) ) ;
    buf_clk cell_3574 ( .C ( clk ), .D ( signal_5933 ), .Q ( signal_5934 ) ) ;
    buf_clk cell_3576 ( .C ( clk ), .D ( signal_5935 ), .Q ( signal_5936 ) ) ;
    buf_clk cell_3578 ( .C ( clk ), .D ( signal_5937 ), .Q ( signal_5938 ) ) ;
    buf_clk cell_3580 ( .C ( clk ), .D ( signal_5939 ), .Q ( signal_5940 ) ) ;
    buf_clk cell_3586 ( .C ( clk ), .D ( signal_5945 ), .Q ( signal_5946 ) ) ;
    buf_clk cell_3592 ( .C ( clk ), .D ( signal_5951 ), .Q ( signal_5952 ) ) ;
    buf_clk cell_3596 ( .C ( clk ), .D ( signal_5955 ), .Q ( signal_5956 ) ) ;
    buf_clk cell_3600 ( .C ( clk ), .D ( signal_5959 ), .Q ( signal_5960 ) ) ;
    buf_clk cell_3602 ( .C ( clk ), .D ( signal_5961 ), .Q ( signal_5962 ) ) ;
    buf_clk cell_3604 ( .C ( clk ), .D ( signal_5963 ), .Q ( signal_5964 ) ) ;
    buf_clk cell_3606 ( .C ( clk ), .D ( signal_5965 ), .Q ( signal_5966 ) ) ;
    buf_clk cell_3608 ( .C ( clk ), .D ( signal_5967 ), .Q ( signal_5968 ) ) ;
    buf_clk cell_3612 ( .C ( clk ), .D ( signal_5971 ), .Q ( signal_5972 ) ) ;
    buf_clk cell_3616 ( .C ( clk ), .D ( signal_5975 ), .Q ( signal_5976 ) ) ;
    buf_clk cell_3620 ( .C ( clk ), .D ( signal_5979 ), .Q ( signal_5980 ) ) ;
    buf_clk cell_3624 ( .C ( clk ), .D ( signal_5983 ), .Q ( signal_5984 ) ) ;
    buf_clk cell_3628 ( .C ( clk ), .D ( signal_5987 ), .Q ( signal_5988 ) ) ;
    buf_clk cell_3632 ( .C ( clk ), .D ( signal_5991 ), .Q ( signal_5992 ) ) ;
    buf_clk cell_3634 ( .C ( clk ), .D ( signal_5993 ), .Q ( signal_5994 ) ) ;
    buf_clk cell_3636 ( .C ( clk ), .D ( signal_5995 ), .Q ( signal_5996 ) ) ;
    buf_clk cell_3642 ( .C ( clk ), .D ( signal_6001 ), .Q ( signal_6002 ) ) ;
    buf_clk cell_3648 ( .C ( clk ), .D ( signal_6007 ), .Q ( signal_6008 ) ) ;
    buf_clk cell_3652 ( .C ( clk ), .D ( signal_6011 ), .Q ( signal_6012 ) ) ;
    buf_clk cell_3656 ( .C ( clk ), .D ( signal_6015 ), .Q ( signal_6016 ) ) ;
    buf_clk cell_3662 ( .C ( clk ), .D ( signal_6021 ), .Q ( signal_6022 ) ) ;
    buf_clk cell_3668 ( .C ( clk ), .D ( signal_6027 ), .Q ( signal_6028 ) ) ;
    buf_clk cell_3672 ( .C ( clk ), .D ( signal_6031 ), .Q ( signal_6032 ) ) ;
    buf_clk cell_3676 ( .C ( clk ), .D ( signal_6035 ), .Q ( signal_6036 ) ) ;
    buf_clk cell_3680 ( .C ( clk ), .D ( signal_6039 ), .Q ( signal_6040 ) ) ;
    buf_clk cell_3684 ( .C ( clk ), .D ( signal_6043 ), .Q ( signal_6044 ) ) ;
    buf_clk cell_3688 ( .C ( clk ), .D ( signal_6047 ), .Q ( signal_6048 ) ) ;
    buf_clk cell_3692 ( .C ( clk ), .D ( signal_6051 ), .Q ( signal_6052 ) ) ;
    buf_clk cell_3694 ( .C ( clk ), .D ( signal_6053 ), .Q ( signal_6054 ) ) ;
    buf_clk cell_3696 ( .C ( clk ), .D ( signal_6055 ), .Q ( signal_6056 ) ) ;
    buf_clk cell_3700 ( .C ( clk ), .D ( signal_6059 ), .Q ( signal_6060 ) ) ;
    buf_clk cell_3704 ( .C ( clk ), .D ( signal_6063 ), .Q ( signal_6064 ) ) ;
    buf_clk cell_3708 ( .C ( clk ), .D ( signal_6067 ), .Q ( signal_6068 ) ) ;
    buf_clk cell_3712 ( .C ( clk ), .D ( signal_6071 ), .Q ( signal_6072 ) ) ;
    buf_clk cell_3718 ( .C ( clk ), .D ( signal_6077 ), .Q ( signal_6078 ) ) ;
    buf_clk cell_3724 ( .C ( clk ), .D ( signal_6083 ), .Q ( signal_6084 ) ) ;
    buf_clk cell_3726 ( .C ( clk ), .D ( signal_6085 ), .Q ( signal_6086 ) ) ;
    buf_clk cell_3728 ( .C ( clk ), .D ( signal_6087 ), .Q ( signal_6088 ) ) ;
    buf_clk cell_3730 ( .C ( clk ), .D ( signal_6089 ), .Q ( signal_6090 ) ) ;
    buf_clk cell_3732 ( .C ( clk ), .D ( signal_6091 ), .Q ( signal_6092 ) ) ;
    buf_clk cell_3736 ( .C ( clk ), .D ( signal_6095 ), .Q ( signal_6096 ) ) ;
    buf_clk cell_3740 ( .C ( clk ), .D ( signal_6099 ), .Q ( signal_6100 ) ) ;
    buf_clk cell_3746 ( .C ( clk ), .D ( signal_6105 ), .Q ( signal_6106 ) ) ;
    buf_clk cell_3752 ( .C ( clk ), .D ( signal_6111 ), .Q ( signal_6112 ) ) ;
    buf_clk cell_3758 ( .C ( clk ), .D ( signal_6117 ), .Q ( signal_6118 ) ) ;
    buf_clk cell_3764 ( .C ( clk ), .D ( signal_6123 ), .Q ( signal_6124 ) ) ;
    buf_clk cell_3770 ( .C ( clk ), .D ( signal_6129 ), .Q ( signal_6130 ) ) ;
    buf_clk cell_3776 ( .C ( clk ), .D ( signal_6135 ), .Q ( signal_6136 ) ) ;
    buf_clk cell_3780 ( .C ( clk ), .D ( signal_6139 ), .Q ( signal_6140 ) ) ;
    buf_clk cell_3784 ( .C ( clk ), .D ( signal_6143 ), .Q ( signal_6144 ) ) ;
    buf_clk cell_3786 ( .C ( clk ), .D ( signal_6145 ), .Q ( signal_6146 ) ) ;
    buf_clk cell_3788 ( .C ( clk ), .D ( signal_6147 ), .Q ( signal_6148 ) ) ;
    buf_clk cell_3790 ( .C ( clk ), .D ( signal_6149 ), .Q ( signal_6150 ) ) ;
    buf_clk cell_3792 ( .C ( clk ), .D ( signal_6151 ), .Q ( signal_6152 ) ) ;
    buf_clk cell_3798 ( .C ( clk ), .D ( signal_6157 ), .Q ( signal_6158 ) ) ;
    buf_clk cell_3806 ( .C ( clk ), .D ( signal_6165 ), .Q ( signal_6166 ) ) ;
    buf_clk cell_3810 ( .C ( clk ), .D ( signal_6169 ), .Q ( signal_6170 ) ) ;
    buf_clk cell_3814 ( .C ( clk ), .D ( signal_6173 ), .Q ( signal_6174 ) ) ;
    buf_clk cell_3820 ( .C ( clk ), .D ( signal_6179 ), .Q ( signal_6180 ) ) ;
    buf_clk cell_3826 ( .C ( clk ), .D ( signal_6185 ), .Q ( signal_6186 ) ) ;
    buf_clk cell_3832 ( .C ( clk ), .D ( signal_6191 ), .Q ( signal_6192 ) ) ;
    buf_clk cell_3838 ( .C ( clk ), .D ( signal_6197 ), .Q ( signal_6198 ) ) ;
    buf_clk cell_3842 ( .C ( clk ), .D ( signal_6201 ), .Q ( signal_6202 ) ) ;
    buf_clk cell_3846 ( .C ( clk ), .D ( signal_6205 ), .Q ( signal_6206 ) ) ;
    buf_clk cell_3852 ( .C ( clk ), .D ( signal_6211 ), .Q ( signal_6212 ) ) ;
    buf_clk cell_3858 ( .C ( clk ), .D ( signal_6217 ), .Q ( signal_6218 ) ) ;
    buf_clk cell_3862 ( .C ( clk ), .D ( signal_6221 ), .Q ( signal_6222 ) ) ;
    buf_clk cell_3866 ( .C ( clk ), .D ( signal_6225 ), .Q ( signal_6226 ) ) ;
    buf_clk cell_3870 ( .C ( clk ), .D ( signal_6229 ), .Q ( signal_6230 ) ) ;
    buf_clk cell_3874 ( .C ( clk ), .D ( signal_6233 ), .Q ( signal_6234 ) ) ;
    buf_clk cell_3888 ( .C ( clk ), .D ( signal_6247 ), .Q ( signal_6248 ) ) ;
    buf_clk cell_3894 ( .C ( clk ), .D ( signal_6253 ), .Q ( signal_6254 ) ) ;
    buf_clk cell_3900 ( .C ( clk ), .D ( signal_6259 ), .Q ( signal_6260 ) ) ;
    buf_clk cell_3906 ( .C ( clk ), .D ( signal_6265 ), .Q ( signal_6266 ) ) ;
    buf_clk cell_3912 ( .C ( clk ), .D ( signal_6271 ), .Q ( signal_6272 ) ) ;
    buf_clk cell_3918 ( .C ( clk ), .D ( signal_6277 ), .Q ( signal_6278 ) ) ;
    buf_clk cell_3926 ( .C ( clk ), .D ( signal_6285 ), .Q ( signal_6286 ) ) ;
    buf_clk cell_3930 ( .C ( clk ), .D ( signal_6289 ), .Q ( signal_6290 ) ) ;
    buf_clk cell_3936 ( .C ( clk ), .D ( signal_6295 ), .Q ( signal_6296 ) ) ;
    buf_clk cell_3942 ( .C ( clk ), .D ( signal_6301 ), .Q ( signal_6302 ) ) ;
    buf_clk cell_3952 ( .C ( clk ), .D ( signal_6311 ), .Q ( signal_6312 ) ) ;
    buf_clk cell_3958 ( .C ( clk ), .D ( signal_6317 ), .Q ( signal_6318 ) ) ;
    buf_clk cell_3970 ( .C ( clk ), .D ( signal_6329 ), .Q ( signal_6330 ) ) ;
    buf_clk cell_3978 ( .C ( clk ), .D ( signal_6337 ), .Q ( signal_6338 ) ) ;
    buf_clk cell_3982 ( .C ( clk ), .D ( signal_6341 ), .Q ( signal_6342 ) ) ;
    buf_clk cell_3986 ( .C ( clk ), .D ( signal_6345 ), .Q ( signal_6346 ) ) ;
    buf_clk cell_3990 ( .C ( clk ), .D ( signal_6349 ), .Q ( signal_6350 ) ) ;
    buf_clk cell_3994 ( .C ( clk ), .D ( signal_6353 ), .Q ( signal_6354 ) ) ;
    buf_clk cell_4000 ( .C ( clk ), .D ( signal_6359 ), .Q ( signal_6360 ) ) ;
    buf_clk cell_4006 ( .C ( clk ), .D ( signal_6365 ), .Q ( signal_6366 ) ) ;
    buf_clk cell_4012 ( .C ( clk ), .D ( signal_6371 ), .Q ( signal_6372 ) ) ;
    buf_clk cell_4018 ( .C ( clk ), .D ( signal_6377 ), .Q ( signal_6378 ) ) ;
    buf_clk cell_4022 ( .C ( clk ), .D ( signal_6381 ), .Q ( signal_6382 ) ) ;
    buf_clk cell_4026 ( .C ( clk ), .D ( signal_6385 ), .Q ( signal_6386 ) ) ;
    buf_clk cell_4034 ( .C ( clk ), .D ( signal_6393 ), .Q ( signal_6394 ) ) ;
    buf_clk cell_4042 ( .C ( clk ), .D ( signal_6401 ), .Q ( signal_6402 ) ) ;
    buf_clk cell_4048 ( .C ( clk ), .D ( signal_6407 ), .Q ( signal_6408 ) ) ;
    buf_clk cell_4054 ( .C ( clk ), .D ( signal_6413 ), .Q ( signal_6414 ) ) ;
    buf_clk cell_4060 ( .C ( clk ), .D ( signal_6419 ), .Q ( signal_6420 ) ) ;
    buf_clk cell_4066 ( .C ( clk ), .D ( signal_6425 ), .Q ( signal_6426 ) ) ;
    buf_clk cell_4080 ( .C ( clk ), .D ( signal_6439 ), .Q ( signal_6440 ) ) ;
    buf_clk cell_4086 ( .C ( clk ), .D ( signal_6445 ), .Q ( signal_6446 ) ) ;
    buf_clk cell_4100 ( .C ( clk ), .D ( signal_6459 ), .Q ( signal_6460 ) ) ;
    buf_clk cell_4106 ( .C ( clk ), .D ( signal_6465 ), .Q ( signal_6466 ) ) ;
    buf_clk cell_4112 ( .C ( clk ), .D ( signal_6471 ), .Q ( signal_6472 ) ) ;
    buf_clk cell_4118 ( .C ( clk ), .D ( signal_6477 ), .Q ( signal_6478 ) ) ;
    buf_clk cell_4122 ( .C ( clk ), .D ( signal_6481 ), .Q ( signal_6482 ) ) ;
    buf_clk cell_4126 ( .C ( clk ), .D ( signal_6485 ), .Q ( signal_6486 ) ) ;
    buf_clk cell_4134 ( .C ( clk ), .D ( signal_6493 ), .Q ( signal_6494 ) ) ;
    buf_clk cell_4144 ( .C ( clk ), .D ( signal_6503 ), .Q ( signal_6504 ) ) ;
    buf_clk cell_4150 ( .C ( clk ), .D ( signal_6509 ), .Q ( signal_6510 ) ) ;
    buf_clk cell_4156 ( .C ( clk ), .D ( signal_6515 ), .Q ( signal_6516 ) ) ;
    buf_clk cell_4164 ( .C ( clk ), .D ( signal_6523 ), .Q ( signal_6524 ) ) ;
    buf_clk cell_4172 ( .C ( clk ), .D ( signal_6531 ), .Q ( signal_6532 ) ) ;
    buf_clk cell_4180 ( .C ( clk ), .D ( signal_6539 ), .Q ( signal_6540 ) ) ;
    buf_clk cell_4188 ( .C ( clk ), .D ( signal_6547 ), .Q ( signal_6548 ) ) ;
    buf_clk cell_4230 ( .C ( clk ), .D ( signal_6589 ), .Q ( signal_6590 ) ) ;
    buf_clk cell_4240 ( .C ( clk ), .D ( signal_6599 ), .Q ( signal_6600 ) ) ;
    buf_clk cell_4246 ( .C ( clk ), .D ( signal_6605 ), .Q ( signal_6606 ) ) ;
    buf_clk cell_4252 ( .C ( clk ), .D ( signal_6611 ), .Q ( signal_6612 ) ) ;
    buf_clk cell_4264 ( .C ( clk ), .D ( signal_6623 ), .Q ( signal_6624 ) ) ;
    buf_clk cell_4272 ( .C ( clk ), .D ( signal_6631 ), .Q ( signal_6632 ) ) ;
    buf_clk cell_4278 ( .C ( clk ), .D ( signal_6637 ), .Q ( signal_6638 ) ) ;
    buf_clk cell_4284 ( .C ( clk ), .D ( signal_6643 ), .Q ( signal_6644 ) ) ;
    buf_clk cell_4292 ( .C ( clk ), .D ( signal_6651 ), .Q ( signal_6652 ) ) ;
    buf_clk cell_4300 ( .C ( clk ), .D ( signal_6659 ), .Q ( signal_6660 ) ) ;
    buf_clk cell_4308 ( .C ( clk ), .D ( signal_6667 ), .Q ( signal_6668 ) ) ;
    buf_clk cell_4316 ( .C ( clk ), .D ( signal_6675 ), .Q ( signal_6676 ) ) ;
    buf_clk cell_4324 ( .C ( clk ), .D ( signal_6683 ), .Q ( signal_6684 ) ) ;
    buf_clk cell_4332 ( .C ( clk ), .D ( signal_6691 ), .Q ( signal_6692 ) ) ;
    buf_clk cell_4342 ( .C ( clk ), .D ( signal_6701 ), .Q ( signal_6702 ) ) ;
    buf_clk cell_4352 ( .C ( clk ), .D ( signal_6711 ), .Q ( signal_6712 ) ) ;
    buf_clk cell_4360 ( .C ( clk ), .D ( signal_6719 ), .Q ( signal_6720 ) ) ;
    buf_clk cell_4368 ( .C ( clk ), .D ( signal_6727 ), .Q ( signal_6728 ) ) ;
    buf_clk cell_4376 ( .C ( clk ), .D ( signal_6735 ), .Q ( signal_6736 ) ) ;
    buf_clk cell_4384 ( .C ( clk ), .D ( signal_6743 ), .Q ( signal_6744 ) ) ;
    buf_clk cell_4396 ( .C ( clk ), .D ( signal_6755 ), .Q ( signal_6756 ) ) ;
    buf_clk cell_4404 ( .C ( clk ), .D ( signal_6763 ), .Q ( signal_6764 ) ) ;
    buf_clk cell_4412 ( .C ( clk ), .D ( signal_6771 ), .Q ( signal_6772 ) ) ;
    buf_clk cell_4420 ( .C ( clk ), .D ( signal_6779 ), .Q ( signal_6780 ) ) ;
    buf_clk cell_4428 ( .C ( clk ), .D ( signal_6787 ), .Q ( signal_6788 ) ) ;
    buf_clk cell_4436 ( .C ( clk ), .D ( signal_6795 ), .Q ( signal_6796 ) ) ;
    buf_clk cell_4454 ( .C ( clk ), .D ( signal_6813 ), .Q ( signal_6814 ) ) ;
    buf_clk cell_4462 ( .C ( clk ), .D ( signal_6821 ), .Q ( signal_6822 ) ) ;
    buf_clk cell_4494 ( .C ( clk ), .D ( signal_6853 ), .Q ( signal_6854 ) ) ;
    buf_clk cell_4502 ( .C ( clk ), .D ( signal_6861 ), .Q ( signal_6862 ) ) ;
    buf_clk cell_4512 ( .C ( clk ), .D ( signal_6871 ), .Q ( signal_6872 ) ) ;
    buf_clk cell_4522 ( .C ( clk ), .D ( signal_6881 ), .Q ( signal_6882 ) ) ;
    buf_clk cell_4546 ( .C ( clk ), .D ( signal_6905 ), .Q ( signal_6906 ) ) ;
    buf_clk cell_4554 ( .C ( clk ), .D ( signal_6913 ), .Q ( signal_6914 ) ) ;
    buf_clk cell_4564 ( .C ( clk ), .D ( signal_6923 ), .Q ( signal_6924 ) ) ;
    buf_clk cell_4574 ( .C ( clk ), .D ( signal_6933 ), .Q ( signal_6934 ) ) ;
    buf_clk cell_4582 ( .C ( clk ), .D ( signal_6941 ), .Q ( signal_6942 ) ) ;
    buf_clk cell_4590 ( .C ( clk ), .D ( signal_6949 ), .Q ( signal_6950 ) ) ;
    buf_clk cell_4742 ( .C ( clk ), .D ( signal_7101 ), .Q ( signal_7102 ) ) ;
    buf_clk cell_4752 ( .C ( clk ), .D ( signal_7111 ), .Q ( signal_7112 ) ) ;
    buf_clk cell_4918 ( .C ( clk ), .D ( signal_7277 ), .Q ( signal_7278 ) ) ;
    buf_clk cell_4930 ( .C ( clk ), .D ( signal_7289 ), .Q ( signal_7290 ) ) ;
    buf_clk cell_4968 ( .C ( clk ), .D ( signal_7327 ), .Q ( signal_7328 ) ) ;
    buf_clk cell_4982 ( .C ( clk ), .D ( signal_7341 ), .Q ( signal_7342 ) ) ;
    buf_clk cell_5012 ( .C ( clk ), .D ( signal_7371 ), .Q ( signal_7372 ) ) ;
    buf_clk cell_5026 ( .C ( clk ), .D ( signal_7385 ), .Q ( signal_7386 ) ) ;
    buf_clk cell_5092 ( .C ( clk ), .D ( signal_7451 ), .Q ( signal_7452 ) ) ;
    buf_clk cell_5108 ( .C ( clk ), .D ( signal_7467 ), .Q ( signal_7468 ) ) ;
    buf_clk cell_5132 ( .C ( clk ), .D ( signal_7491 ), .Q ( signal_7492 ) ) ;
    buf_clk cell_5148 ( .C ( clk ), .D ( signal_7507 ), .Q ( signal_7508 ) ) ;
    buf_clk cell_5254 ( .C ( clk ), .D ( signal_7613 ), .Q ( signal_7614 ) ) ;
    buf_clk cell_5270 ( .C ( clk ), .D ( signal_7629 ), .Q ( signal_7630 ) ) ;
    buf_clk cell_5288 ( .C ( clk ), .D ( signal_7647 ), .Q ( signal_7648 ) ) ;
    buf_clk cell_5306 ( .C ( clk ), .D ( signal_7665 ), .Q ( signal_7666 ) ) ;
    buf_clk cell_5388 ( .C ( clk ), .D ( signal_7747 ), .Q ( signal_7748 ) ) ;
    buf_clk cell_5408 ( .C ( clk ), .D ( signal_7767 ), .Q ( signal_7768 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_3799 ( .C ( clk ), .D ( signal_6158 ), .Q ( signal_6159 ) ) ;
    buf_clk cell_3807 ( .C ( clk ), .D ( signal_6166 ), .Q ( signal_6167 ) ) ;
    buf_clk cell_3811 ( .C ( clk ), .D ( signal_6170 ), .Q ( signal_6171 ) ) ;
    buf_clk cell_3815 ( .C ( clk ), .D ( signal_6174 ), .Q ( signal_6175 ) ) ;
    buf_clk cell_3821 ( .C ( clk ), .D ( signal_6180 ), .Q ( signal_6181 ) ) ;
    buf_clk cell_3827 ( .C ( clk ), .D ( signal_6186 ), .Q ( signal_6187 ) ) ;
    buf_clk cell_3833 ( .C ( clk ), .D ( signal_6192 ), .Q ( signal_6193 ) ) ;
    buf_clk cell_3839 ( .C ( clk ), .D ( signal_6198 ), .Q ( signal_6199 ) ) ;
    buf_clk cell_3843 ( .C ( clk ), .D ( signal_6202 ), .Q ( signal_6203 ) ) ;
    buf_clk cell_3847 ( .C ( clk ), .D ( signal_6206 ), .Q ( signal_6207 ) ) ;
    buf_clk cell_3853 ( .C ( clk ), .D ( signal_6212 ), .Q ( signal_6213 ) ) ;
    buf_clk cell_3859 ( .C ( clk ), .D ( signal_6218 ), .Q ( signal_6219 ) ) ;
    buf_clk cell_3863 ( .C ( clk ), .D ( signal_6222 ), .Q ( signal_6223 ) ) ;
    buf_clk cell_3867 ( .C ( clk ), .D ( signal_6226 ), .Q ( signal_6227 ) ) ;
    buf_clk cell_3871 ( .C ( clk ), .D ( signal_6230 ), .Q ( signal_6231 ) ) ;
    buf_clk cell_3875 ( .C ( clk ), .D ( signal_6234 ), .Q ( signal_6235 ) ) ;
    buf_clk cell_3877 ( .C ( clk ), .D ( signal_2071 ), .Q ( signal_6237 ) ) ;
    buf_clk cell_3879 ( .C ( clk ), .D ( signal_3529 ), .Q ( signal_6239 ) ) ;
    buf_clk cell_3881 ( .C ( clk ), .D ( signal_5994 ), .Q ( signal_6241 ) ) ;
    buf_clk cell_3883 ( .C ( clk ), .D ( signal_5996 ), .Q ( signal_6243 ) ) ;
    buf_clk cell_3889 ( .C ( clk ), .D ( signal_6248 ), .Q ( signal_6249 ) ) ;
    buf_clk cell_3895 ( .C ( clk ), .D ( signal_6254 ), .Q ( signal_6255 ) ) ;
    buf_clk cell_3901 ( .C ( clk ), .D ( signal_6260 ), .Q ( signal_6261 ) ) ;
    buf_clk cell_3907 ( .C ( clk ), .D ( signal_6266 ), .Q ( signal_6267 ) ) ;
    buf_clk cell_3913 ( .C ( clk ), .D ( signal_6272 ), .Q ( signal_6273 ) ) ;
    buf_clk cell_3919 ( .C ( clk ), .D ( signal_6278 ), .Q ( signal_6279 ) ) ;
    buf_clk cell_3921 ( .C ( clk ), .D ( signal_5864 ), .Q ( signal_6281 ) ) ;
    buf_clk cell_3923 ( .C ( clk ), .D ( signal_5868 ), .Q ( signal_6283 ) ) ;
    buf_clk cell_3927 ( .C ( clk ), .D ( signal_6286 ), .Q ( signal_6287 ) ) ;
    buf_clk cell_3931 ( .C ( clk ), .D ( signal_6290 ), .Q ( signal_6291 ) ) ;
    buf_clk cell_3937 ( .C ( clk ), .D ( signal_6296 ), .Q ( signal_6297 ) ) ;
    buf_clk cell_3943 ( .C ( clk ), .D ( signal_6302 ), .Q ( signal_6303 ) ) ;
    buf_clk cell_3945 ( .C ( clk ), .D ( signal_2081 ), .Q ( signal_6305 ) ) ;
    buf_clk cell_3947 ( .C ( clk ), .D ( signal_3539 ), .Q ( signal_6307 ) ) ;
    buf_clk cell_3953 ( .C ( clk ), .D ( signal_6312 ), .Q ( signal_6313 ) ) ;
    buf_clk cell_3959 ( .C ( clk ), .D ( signal_6318 ), .Q ( signal_6319 ) ) ;
    buf_clk cell_3961 ( .C ( clk ), .D ( signal_2069 ), .Q ( signal_6321 ) ) ;
    buf_clk cell_3963 ( .C ( clk ), .D ( signal_3527 ), .Q ( signal_6323 ) ) ;
    buf_clk cell_3971 ( .C ( clk ), .D ( signal_6330 ), .Q ( signal_6331 ) ) ;
    buf_clk cell_3979 ( .C ( clk ), .D ( signal_6338 ), .Q ( signal_6339 ) ) ;
    buf_clk cell_3983 ( .C ( clk ), .D ( signal_6342 ), .Q ( signal_6343 ) ) ;
    buf_clk cell_3987 ( .C ( clk ), .D ( signal_6346 ), .Q ( signal_6347 ) ) ;
    buf_clk cell_3991 ( .C ( clk ), .D ( signal_6350 ), .Q ( signal_6351 ) ) ;
    buf_clk cell_3995 ( .C ( clk ), .D ( signal_6354 ), .Q ( signal_6355 ) ) ;
    buf_clk cell_4001 ( .C ( clk ), .D ( signal_6360 ), .Q ( signal_6361 ) ) ;
    buf_clk cell_4007 ( .C ( clk ), .D ( signal_6366 ), .Q ( signal_6367 ) ) ;
    buf_clk cell_4013 ( .C ( clk ), .D ( signal_6372 ), .Q ( signal_6373 ) ) ;
    buf_clk cell_4019 ( .C ( clk ), .D ( signal_6378 ), .Q ( signal_6379 ) ) ;
    buf_clk cell_4023 ( .C ( clk ), .D ( signal_6382 ), .Q ( signal_6383 ) ) ;
    buf_clk cell_4027 ( .C ( clk ), .D ( signal_6386 ), .Q ( signal_6387 ) ) ;
    buf_clk cell_4035 ( .C ( clk ), .D ( signal_6394 ), .Q ( signal_6395 ) ) ;
    buf_clk cell_4043 ( .C ( clk ), .D ( signal_6402 ), .Q ( signal_6403 ) ) ;
    buf_clk cell_4049 ( .C ( clk ), .D ( signal_6408 ), .Q ( signal_6409 ) ) ;
    buf_clk cell_4055 ( .C ( clk ), .D ( signal_6414 ), .Q ( signal_6415 ) ) ;
    buf_clk cell_4061 ( .C ( clk ), .D ( signal_6420 ), .Q ( signal_6421 ) ) ;
    buf_clk cell_4067 ( .C ( clk ), .D ( signal_6426 ), .Q ( signal_6427 ) ) ;
    buf_clk cell_4069 ( .C ( clk ), .D ( signal_2201 ), .Q ( signal_6429 ) ) ;
    buf_clk cell_4071 ( .C ( clk ), .D ( signal_3659 ), .Q ( signal_6431 ) ) ;
    buf_clk cell_4073 ( .C ( clk ), .D ( signal_5938 ), .Q ( signal_6433 ) ) ;
    buf_clk cell_4075 ( .C ( clk ), .D ( signal_5940 ), .Q ( signal_6435 ) ) ;
    buf_clk cell_4081 ( .C ( clk ), .D ( signal_6440 ), .Q ( signal_6441 ) ) ;
    buf_clk cell_4087 ( .C ( clk ), .D ( signal_6446 ), .Q ( signal_6447 ) ) ;
    buf_clk cell_4089 ( .C ( clk ), .D ( signal_5934 ), .Q ( signal_6449 ) ) ;
    buf_clk cell_4091 ( .C ( clk ), .D ( signal_5936 ), .Q ( signal_6451 ) ) ;
    buf_clk cell_4093 ( .C ( clk ), .D ( signal_5758 ), .Q ( signal_6453 ) ) ;
    buf_clk cell_4095 ( .C ( clk ), .D ( signal_5764 ), .Q ( signal_6455 ) ) ;
    buf_clk cell_4101 ( .C ( clk ), .D ( signal_6460 ), .Q ( signal_6461 ) ) ;
    buf_clk cell_4107 ( .C ( clk ), .D ( signal_6466 ), .Q ( signal_6467 ) ) ;
    buf_clk cell_4113 ( .C ( clk ), .D ( signal_6472 ), .Q ( signal_6473 ) ) ;
    buf_clk cell_4119 ( .C ( clk ), .D ( signal_6478 ), .Q ( signal_6479 ) ) ;
    buf_clk cell_4123 ( .C ( clk ), .D ( signal_6482 ), .Q ( signal_6483 ) ) ;
    buf_clk cell_4127 ( .C ( clk ), .D ( signal_6486 ), .Q ( signal_6487 ) ) ;
    buf_clk cell_4135 ( .C ( clk ), .D ( signal_6494 ), .Q ( signal_6495 ) ) ;
    buf_clk cell_4145 ( .C ( clk ), .D ( signal_6504 ), .Q ( signal_6505 ) ) ;
    buf_clk cell_4151 ( .C ( clk ), .D ( signal_6510 ), .Q ( signal_6511 ) ) ;
    buf_clk cell_4157 ( .C ( clk ), .D ( signal_6516 ), .Q ( signal_6517 ) ) ;
    buf_clk cell_4165 ( .C ( clk ), .D ( signal_6524 ), .Q ( signal_6525 ) ) ;
    buf_clk cell_4173 ( .C ( clk ), .D ( signal_6532 ), .Q ( signal_6533 ) ) ;
    buf_clk cell_4181 ( .C ( clk ), .D ( signal_6540 ), .Q ( signal_6541 ) ) ;
    buf_clk cell_4189 ( .C ( clk ), .D ( signal_6548 ), .Q ( signal_6549 ) ) ;
    buf_clk cell_4193 ( .C ( clk ), .D ( signal_5906 ), .Q ( signal_6553 ) ) ;
    buf_clk cell_4197 ( .C ( clk ), .D ( signal_5908 ), .Q ( signal_6557 ) ) ;
    buf_clk cell_4201 ( .C ( clk ), .D ( signal_2116 ), .Q ( signal_6561 ) ) ;
    buf_clk cell_4205 ( .C ( clk ), .D ( signal_3574 ), .Q ( signal_6565 ) ) ;
    buf_clk cell_4217 ( .C ( clk ), .D ( signal_2109 ), .Q ( signal_6577 ) ) ;
    buf_clk cell_4221 ( .C ( clk ), .D ( signal_3567 ), .Q ( signal_6581 ) ) ;
    buf_clk cell_4231 ( .C ( clk ), .D ( signal_6590 ), .Q ( signal_6591 ) ) ;
    buf_clk cell_4241 ( .C ( clk ), .D ( signal_6600 ), .Q ( signal_6601 ) ) ;
    buf_clk cell_4247 ( .C ( clk ), .D ( signal_6606 ), .Q ( signal_6607 ) ) ;
    buf_clk cell_4253 ( .C ( clk ), .D ( signal_6612 ), .Q ( signal_6613 ) ) ;
    buf_clk cell_4265 ( .C ( clk ), .D ( signal_6624 ), .Q ( signal_6625 ) ) ;
    buf_clk cell_4273 ( .C ( clk ), .D ( signal_6632 ), .Q ( signal_6633 ) ) ;
    buf_clk cell_4279 ( .C ( clk ), .D ( signal_6638 ), .Q ( signal_6639 ) ) ;
    buf_clk cell_4285 ( .C ( clk ), .D ( signal_6644 ), .Q ( signal_6645 ) ) ;
    buf_clk cell_4293 ( .C ( clk ), .D ( signal_6652 ), .Q ( signal_6653 ) ) ;
    buf_clk cell_4301 ( .C ( clk ), .D ( signal_6660 ), .Q ( signal_6661 ) ) ;
    buf_clk cell_4309 ( .C ( clk ), .D ( signal_6668 ), .Q ( signal_6669 ) ) ;
    buf_clk cell_4317 ( .C ( clk ), .D ( signal_6676 ), .Q ( signal_6677 ) ) ;
    buf_clk cell_4325 ( .C ( clk ), .D ( signal_6684 ), .Q ( signal_6685 ) ) ;
    buf_clk cell_4333 ( .C ( clk ), .D ( signal_6692 ), .Q ( signal_6693 ) ) ;
    buf_clk cell_4343 ( .C ( clk ), .D ( signal_6702 ), .Q ( signal_6703 ) ) ;
    buf_clk cell_4353 ( .C ( clk ), .D ( signal_6712 ), .Q ( signal_6713 ) ) ;
    buf_clk cell_4361 ( .C ( clk ), .D ( signal_6720 ), .Q ( signal_6721 ) ) ;
    buf_clk cell_4369 ( .C ( clk ), .D ( signal_6728 ), .Q ( signal_6729 ) ) ;
    buf_clk cell_4377 ( .C ( clk ), .D ( signal_6736 ), .Q ( signal_6737 ) ) ;
    buf_clk cell_4385 ( .C ( clk ), .D ( signal_6744 ), .Q ( signal_6745 ) ) ;
    buf_clk cell_4397 ( .C ( clk ), .D ( signal_6756 ), .Q ( signal_6757 ) ) ;
    buf_clk cell_4405 ( .C ( clk ), .D ( signal_6764 ), .Q ( signal_6765 ) ) ;
    buf_clk cell_4413 ( .C ( clk ), .D ( signal_6772 ), .Q ( signal_6773 ) ) ;
    buf_clk cell_4421 ( .C ( clk ), .D ( signal_6780 ), .Q ( signal_6781 ) ) ;
    buf_clk cell_4429 ( .C ( clk ), .D ( signal_6788 ), .Q ( signal_6789 ) ) ;
    buf_clk cell_4437 ( .C ( clk ), .D ( signal_6796 ), .Q ( signal_6797 ) ) ;
    buf_clk cell_4441 ( .C ( clk ), .D ( signal_1945 ), .Q ( signal_6801 ) ) ;
    buf_clk cell_4447 ( .C ( clk ), .D ( signal_3403 ), .Q ( signal_6807 ) ) ;
    buf_clk cell_4455 ( .C ( clk ), .D ( signal_6814 ), .Q ( signal_6815 ) ) ;
    buf_clk cell_4463 ( .C ( clk ), .D ( signal_6822 ), .Q ( signal_6823 ) ) ;
    buf_clk cell_4469 ( .C ( clk ), .D ( signal_2111 ), .Q ( signal_6829 ) ) ;
    buf_clk cell_4475 ( .C ( clk ), .D ( signal_3569 ), .Q ( signal_6835 ) ) ;
    buf_clk cell_4481 ( .C ( clk ), .D ( signal_1976 ), .Q ( signal_6841 ) ) ;
    buf_clk cell_4487 ( .C ( clk ), .D ( signal_3434 ), .Q ( signal_6847 ) ) ;
    buf_clk cell_4495 ( .C ( clk ), .D ( signal_6854 ), .Q ( signal_6855 ) ) ;
    buf_clk cell_4503 ( .C ( clk ), .D ( signal_6862 ), .Q ( signal_6863 ) ) ;
    buf_clk cell_4513 ( .C ( clk ), .D ( signal_6872 ), .Q ( signal_6873 ) ) ;
    buf_clk cell_4523 ( .C ( clk ), .D ( signal_6882 ), .Q ( signal_6883 ) ) ;
    buf_clk cell_4533 ( .C ( clk ), .D ( signal_2070 ), .Q ( signal_6893 ) ) ;
    buf_clk cell_4539 ( .C ( clk ), .D ( signal_3528 ), .Q ( signal_6899 ) ) ;
    buf_clk cell_4547 ( .C ( clk ), .D ( signal_6906 ), .Q ( signal_6907 ) ) ;
    buf_clk cell_4555 ( .C ( clk ), .D ( signal_6914 ), .Q ( signal_6915 ) ) ;
    buf_clk cell_4565 ( .C ( clk ), .D ( signal_6924 ), .Q ( signal_6925 ) ) ;
    buf_clk cell_4575 ( .C ( clk ), .D ( signal_6934 ), .Q ( signal_6935 ) ) ;
    buf_clk cell_4583 ( .C ( clk ), .D ( signal_6942 ), .Q ( signal_6943 ) ) ;
    buf_clk cell_4591 ( .C ( clk ), .D ( signal_6950 ), .Q ( signal_6951 ) ) ;
    buf_clk cell_4597 ( .C ( clk ), .D ( signal_1890 ), .Q ( signal_6957 ) ) ;
    buf_clk cell_4603 ( .C ( clk ), .D ( signal_3348 ), .Q ( signal_6963 ) ) ;
    buf_clk cell_4609 ( .C ( clk ), .D ( signal_2002 ), .Q ( signal_6969 ) ) ;
    buf_clk cell_4615 ( .C ( clk ), .D ( signal_3460 ), .Q ( signal_6975 ) ) ;
    buf_clk cell_4641 ( .C ( clk ), .D ( signal_2106 ), .Q ( signal_7001 ) ) ;
    buf_clk cell_4647 ( .C ( clk ), .D ( signal_3564 ), .Q ( signal_7007 ) ) ;
    buf_clk cell_4657 ( .C ( clk ), .D ( signal_2068 ), .Q ( signal_7017 ) ) ;
    buf_clk cell_4663 ( .C ( clk ), .D ( signal_3526 ), .Q ( signal_7023 ) ) ;
    buf_clk cell_4677 ( .C ( clk ), .D ( signal_2073 ), .Q ( signal_7037 ) ) ;
    buf_clk cell_4683 ( .C ( clk ), .D ( signal_3531 ), .Q ( signal_7043 ) ) ;
    buf_clk cell_4713 ( .C ( clk ), .D ( signal_2110 ), .Q ( signal_7073 ) ) ;
    buf_clk cell_4721 ( .C ( clk ), .D ( signal_3568 ), .Q ( signal_7081 ) ) ;
    buf_clk cell_4743 ( .C ( clk ), .D ( signal_7102 ), .Q ( signal_7103 ) ) ;
    buf_clk cell_4753 ( .C ( clk ), .D ( signal_7112 ), .Q ( signal_7113 ) ) ;
    buf_clk cell_4781 ( .C ( clk ), .D ( signal_5956 ), .Q ( signal_7141 ) ) ;
    buf_clk cell_4789 ( .C ( clk ), .D ( signal_5960 ), .Q ( signal_7149 ) ) ;
    buf_clk cell_4809 ( .C ( clk ), .D ( signal_1986 ), .Q ( signal_7169 ) ) ;
    buf_clk cell_4817 ( .C ( clk ), .D ( signal_3444 ), .Q ( signal_7177 ) ) ;
    buf_clk cell_4837 ( .C ( clk ), .D ( signal_2082 ), .Q ( signal_7197 ) ) ;
    buf_clk cell_4845 ( .C ( clk ), .D ( signal_3540 ), .Q ( signal_7205 ) ) ;
    buf_clk cell_4919 ( .C ( clk ), .D ( signal_7278 ), .Q ( signal_7279 ) ) ;
    buf_clk cell_4931 ( .C ( clk ), .D ( signal_7290 ), .Q ( signal_7291 ) ) ;
    buf_clk cell_4969 ( .C ( clk ), .D ( signal_7328 ), .Q ( signal_7329 ) ) ;
    buf_clk cell_4983 ( .C ( clk ), .D ( signal_7342 ), .Q ( signal_7343 ) ) ;
    buf_clk cell_5013 ( .C ( clk ), .D ( signal_7372 ), .Q ( signal_7373 ) ) ;
    buf_clk cell_5027 ( .C ( clk ), .D ( signal_7386 ), .Q ( signal_7387 ) ) ;
    buf_clk cell_5093 ( .C ( clk ), .D ( signal_7452 ), .Q ( signal_7453 ) ) ;
    buf_clk cell_5109 ( .C ( clk ), .D ( signal_7468 ), .Q ( signal_7469 ) ) ;
    buf_clk cell_5133 ( .C ( clk ), .D ( signal_7492 ), .Q ( signal_7493 ) ) ;
    buf_clk cell_5149 ( .C ( clk ), .D ( signal_7508 ), .Q ( signal_7509 ) ) ;
    buf_clk cell_5255 ( .C ( clk ), .D ( signal_7614 ), .Q ( signal_7615 ) ) ;
    buf_clk cell_5271 ( .C ( clk ), .D ( signal_7630 ), .Q ( signal_7631 ) ) ;
    buf_clk cell_5289 ( .C ( clk ), .D ( signal_7648 ), .Q ( signal_7649 ) ) ;
    buf_clk cell_5307 ( .C ( clk ), .D ( signal_7666 ), .Q ( signal_7667 ) ) ;
    buf_clk cell_5389 ( .C ( clk ), .D ( signal_7748 ), .Q ( signal_7749 ) ) ;
    buf_clk cell_5409 ( .C ( clk ), .D ( signal_7768 ), .Q ( signal_7769 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2027 ( .a ({signal_5752, signal_5750}), .b ({signal_3384, signal_1926}), .clk ( clk ), .r ( Fresh[665] ), .c ({signal_3500, signal_2042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2032 ( .a ({signal_5764, signal_5758}), .b ({signal_3345, signal_1887}), .clk ( clk ), .r ( Fresh[666] ), .c ({signal_3505, signal_2047}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2037 ( .a ({signal_5776, signal_5770}), .b ({signal_3398, signal_1940}), .clk ( clk ), .r ( Fresh[667] ), .c ({signal_3510, signal_2052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2038 ( .a ({signal_5788, signal_5782}), .b ({signal_3401, signal_1943}), .clk ( clk ), .r ( Fresh[668] ), .c ({signal_3511, signal_2053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2039 ( .a ({signal_5796, signal_5792}), .b ({signal_3404, signal_1946}), .clk ( clk ), .r ( Fresh[669] ), .c ({signal_3512, signal_2054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2040 ( .a ({signal_5808, signal_5802}), .b ({signal_3406, signal_1948}), .clk ( clk ), .r ( Fresh[670] ), .c ({signal_3513, signal_2055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2041 ( .a ({signal_5816, signal_5812}), .b ({signal_3408, signal_1950}), .clk ( clk ), .r ( Fresh[671] ), .c ({signal_3514, signal_2056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2042 ( .a ({signal_5824, signal_5820}), .b ({signal_3412, signal_1954}), .clk ( clk ), .r ( Fresh[672] ), .c ({signal_3515, signal_2057}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2043 ( .a ({signal_5832, signal_5828}), .b ({signal_3413, signal_1955}), .clk ( clk ), .r ( Fresh[673] ), .c ({signal_3516, signal_2058}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2044 ( .a ({signal_5840, signal_5836}), .b ({signal_3414, signal_1956}), .clk ( clk ), .r ( Fresh[674] ), .c ({signal_3517, signal_2059}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2045 ( .a ({signal_5848, signal_5844}), .b ({signal_3419, signal_1961}), .clk ( clk ), .r ( Fresh[675] ), .c ({signal_3518, signal_2060}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2064 ( .a ({signal_3500, signal_2042}), .b ({signal_3537, signal_2079}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2068 ( .a ({signal_3505, signal_2047}), .b ({signal_3541, signal_2083}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2072 ( .a ({signal_3510, signal_2052}), .b ({signal_3545, signal_2087}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2073 ( .a ({signal_3516, signal_2058}), .b ({signal_3546, signal_2088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2084 ( .a ({signal_5860, signal_5854}), .b ({signal_3442, signal_1984}), .clk ( clk ), .r ( Fresh[676] ), .c ({signal_3557, signal_2099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2090 ( .a ({signal_5868, signal_5864}), .b ({signal_3451, signal_1993}), .clk ( clk ), .r ( Fresh[677] ), .c ({signal_3563, signal_2105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2098 ( .a ({signal_3391, signal_1933}), .b ({signal_5872, signal_5870}), .clk ( clk ), .r ( Fresh[678] ), .c ({signal_3571, signal_2113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2100 ( .a ({signal_5876, signal_5874}), .b ({signal_3459, signal_2001}), .clk ( clk ), .r ( Fresh[679] ), .c ({signal_3573, signal_2115}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2102 ( .a ({signal_5880, signal_5878}), .b ({signal_3462, signal_2004}), .clk ( clk ), .r ( Fresh[680] ), .c ({signal_3575, signal_2117}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2103 ( .a ({signal_5884, signal_5882}), .b ({signal_3399, signal_1941}), .clk ( clk ), .r ( Fresh[681] ), .c ({signal_3576, signal_2118}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2105 ( .a ({signal_5888, signal_5886}), .b ({signal_3399, signal_1941}), .clk ( clk ), .r ( Fresh[682] ), .c ({signal_3578, signal_2120}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2106 ( .a ({signal_5896, signal_5892}), .b ({signal_3498, signal_2040}), .clk ( clk ), .r ( Fresh[683] ), .c ({signal_3579, signal_2121}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2107 ( .a ({signal_5900, signal_5898}), .b ({signal_3402, signal_1944}), .clk ( clk ), .r ( Fresh[684] ), .c ({signal_3580, signal_2122}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2108 ( .a ({signal_5904, signal_5902}), .b ({signal_3503, signal_2045}), .clk ( clk ), .r ( Fresh[685] ), .c ({signal_3581, signal_2123}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2109 ( .a ({signal_5908, signal_5906}), .b ({signal_3465, signal_2007}), .clk ( clk ), .r ( Fresh[686] ), .c ({signal_3582, signal_2124}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2111 ( .a ({signal_5920, signal_5914}), .b ({signal_3466, signal_2008}), .clk ( clk ), .r ( Fresh[687] ), .c ({signal_3584, signal_2126}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2112 ( .a ({signal_5924, signal_5922}), .b ({signal_3410, signal_1952}), .clk ( clk ), .r ( Fresh[688] ), .c ({signal_3585, signal_2127}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2113 ( .a ({signal_5932, signal_5928}), .b ({signal_3507, signal_2049}), .clk ( clk ), .r ( Fresh[689] ), .c ({signal_3586, signal_2128}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2114 ( .a ({signal_5936, signal_5934}), .b ({signal_3467, signal_2009}), .clk ( clk ), .r ( Fresh[690] ), .c ({signal_3587, signal_2129}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2115 ( .a ({signal_5860, signal_5854}), .b ({signal_3468, signal_2010}), .clk ( clk ), .r ( Fresh[691] ), .c ({signal_3588, signal_2130}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2117 ( .a ({signal_5940, signal_5938}), .b ({signal_3470, signal_2012}), .clk ( clk ), .r ( Fresh[692] ), .c ({signal_3590, signal_2132}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2120 ( .a ({signal_5868, signal_5864}), .b ({signal_3471, signal_2013}), .clk ( clk ), .r ( Fresh[693] ), .c ({signal_3593, signal_2135}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2129 ( .a ({signal_3557, signal_2099}), .b ({signal_3602, signal_2144}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2131 ( .a ({signal_3563, signal_2105}), .b ({signal_3604, signal_2146}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2132 ( .a ({signal_3573, signal_2115}), .b ({signal_3605, signal_2147}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2134 ( .a ({signal_3582, signal_2124}), .b ({signal_3607, signal_2149}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2136 ( .a ({signal_3584, signal_2126}), .b ({signal_3609, signal_2151}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2137 ( .a ({signal_3587, signal_2129}), .b ({signal_3610, signal_2152}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2138 ( .a ({signal_3588, signal_2130}), .b ({signal_3611, signal_2153}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2139 ( .a ({signal_3590, signal_2132}), .b ({signal_3612, signal_2154}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2141 ( .a ({signal_3593, signal_2135}), .b ({signal_3614, signal_2156}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2142 ( .a ({signal_5952, signal_5946}), .b ({signal_3519, signal_2061}), .clk ( clk ), .r ( Fresh[694] ), .c ({signal_3615, signal_2157}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2143 ( .a ({signal_5960, signal_5956}), .b ({signal_3520, signal_2062}), .clk ( clk ), .r ( Fresh[695] ), .c ({signal_3616, signal_2158}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2145 ( .a ({signal_5964, signal_5962}), .b ({signal_3548, signal_2090}), .clk ( clk ), .r ( Fresh[696] ), .c ({signal_3618, signal_2160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2146 ( .a ({signal_3523, signal_2065}), .b ({signal_5968, signal_5966}), .clk ( clk ), .r ( Fresh[697] ), .c ({signal_3619, signal_2161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2147 ( .a ({signal_5976, signal_5972}), .b ({signal_3524, signal_2066}), .clk ( clk ), .r ( Fresh[698] ), .c ({signal_3620, signal_2162}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2149 ( .a ({signal_5984, signal_5980}), .b ({signal_3551, signal_2093}), .clk ( clk ), .r ( Fresh[699] ), .c ({signal_3622, signal_2164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2150 ( .a ({signal_5992, signal_5988}), .b ({signal_3552, signal_2094}), .clk ( clk ), .r ( Fresh[700] ), .c ({signal_3623, signal_2165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2151 ( .a ({signal_5996, signal_5994}), .b ({signal_3530, signal_2072}), .clk ( clk ), .r ( Fresh[701] ), .c ({signal_3624, signal_2166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2152 ( .a ({signal_6008, signal_6002}), .b ({signal_3553, signal_2095}), .clk ( clk ), .r ( Fresh[702] ), .c ({signal_3625, signal_2167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2153 ( .a ({signal_6016, signal_6012}), .b ({signal_3556, signal_2098}), .clk ( clk ), .r ( Fresh[703] ), .c ({signal_3626, signal_2168}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2154 ( .a ({signal_6028, signal_6022}), .b ({signal_3533, signal_2075}), .clk ( clk ), .r ( Fresh[704] ), .c ({signal_3627, signal_2169}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2155 ( .a ({signal_3522, signal_2064}), .b ({signal_3534, signal_2076}), .clk ( clk ), .r ( Fresh[705] ), .c ({signal_3628, signal_2170}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2156 ( .a ({signal_6036, signal_6032}), .b ({signal_3535, signal_2077}), .clk ( clk ), .r ( Fresh[706] ), .c ({signal_3629, signal_2171}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2157 ( .a ({signal_5764, signal_5758}), .b ({signal_3536, signal_2078}), .clk ( clk ), .r ( Fresh[707] ), .c ({signal_3630, signal_2172}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2158 ( .a ({signal_6044, signal_6040}), .b ({signal_3558, signal_2100}), .clk ( clk ), .r ( Fresh[708] ), .c ({signal_3631, signal_2173}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2159 ( .a ({signal_6052, signal_6048}), .b ({signal_3560, signal_2102}), .clk ( clk ), .r ( Fresh[709] ), .c ({signal_3632, signal_2174}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2160 ( .a ({signal_6056, signal_6054}), .b ({signal_3561, signal_2103}), .clk ( clk ), .r ( Fresh[710] ), .c ({signal_3633, signal_2175}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2161 ( .a ({signal_6064, signal_6060}), .b ({signal_3562, signal_2104}), .clk ( clk ), .r ( Fresh[711] ), .c ({signal_3634, signal_2176}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2163 ( .a ({signal_6072, signal_6068}), .b ({signal_3538, signal_2080}), .clk ( clk ), .r ( Fresh[712] ), .c ({signal_3636, signal_2178}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2164 ( .a ({signal_6084, signal_6078}), .b ({signal_3565, signal_2107}), .clk ( clk ), .r ( Fresh[713] ), .c ({signal_3637, signal_2179}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2165 ( .a ({signal_3566, signal_2108}), .b ({signal_3411, signal_1953}), .clk ( clk ), .r ( Fresh[714] ), .c ({signal_3638, signal_2180}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2166 ( .a ({signal_5764, signal_5758}), .b ({signal_3542, signal_2084}), .clk ( clk ), .r ( Fresh[715] ), .c ({signal_3639, signal_2181}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2167 ( .a ({signal_3543, signal_2085}), .b ({signal_6088, signal_6086}), .clk ( clk ), .r ( Fresh[716] ), .c ({signal_3640, signal_2182}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2168 ( .a ({signal_6092, signal_6090}), .b ({signal_3570, signal_2112}), .clk ( clk ), .r ( Fresh[717] ), .c ({signal_3641, signal_2183}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2169 ( .a ({signal_6100, signal_6096}), .b ({signal_3544, signal_2086}), .clk ( clk ), .r ( Fresh[718] ), .c ({signal_3642, signal_2184}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2171 ( .a ({signal_6112, signal_6106}), .b ({signal_3572, signal_2114}), .clk ( clk ), .r ( Fresh[719] ), .c ({signal_3644, signal_2186}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2184 ( .a ({signal_3616, signal_2158}), .b ({signal_3657, signal_2199}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2187 ( .a ({signal_3624, signal_2166}), .b ({signal_3660, signal_2202}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2188 ( .a ({signal_3630, signal_2172}), .b ({signal_3661, signal_2203}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2189 ( .a ({signal_3632, signal_2174}), .b ({signal_3662, signal_2204}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2191 ( .a ({signal_3637, signal_2179}), .b ({signal_3664, signal_2206}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2192 ( .a ({signal_3638, signal_2180}), .b ({signal_3665, signal_2207}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2193 ( .a ({signal_3639, signal_2181}), .b ({signal_3666, signal_2208}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2194 ( .a ({signal_3644, signal_2186}), .b ({signal_3667, signal_2209}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2201 ( .a ({signal_6124, signal_6118}), .b ({signal_3597, signal_2139}), .clk ( clk ), .r ( Fresh[720] ), .c ({signal_3674, signal_2216}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2202 ( .a ({signal_6136, signal_6130}), .b ({signal_3598, signal_2140}), .clk ( clk ), .r ( Fresh[721] ), .c ({signal_3675, signal_2217}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2203 ( .a ({signal_6144, signal_6140}), .b ({signal_3599, signal_2141}), .clk ( clk ), .r ( Fresh[722] ), .c ({signal_3676, signal_2218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2204 ( .a ({signal_5764, signal_5758}), .b ({signal_3600, signal_2142}), .clk ( clk ), .r ( Fresh[723] ), .c ({signal_3677, signal_2219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2205 ( .a ({signal_6148, signal_6146}), .b ({signal_3601, signal_2143}), .clk ( clk ), .r ( Fresh[724] ), .c ({signal_3678, signal_2220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2206 ( .a ({signal_5936, signal_5934}), .b ({signal_3603, signal_2145}), .clk ( clk ), .r ( Fresh[725] ), .c ({signal_3679, signal_2221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2213 ( .a ({signal_6152, signal_6150}), .b ({signal_3606, signal_2148}), .clk ( clk ), .r ( Fresh[726] ), .c ({signal_3686, signal_2228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2221 ( .a ({signal_6136, signal_6130}), .b ({signal_3608, signal_2150}), .clk ( clk ), .r ( Fresh[727] ), .c ({signal_3694, signal_2236}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2233 ( .a ({signal_3674, signal_2216}), .b ({signal_3706, signal_2248}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2234 ( .a ({signal_3675, signal_2217}), .b ({signal_3707, signal_2249}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2235 ( .a ({signal_3676, signal_2218}), .b ({signal_3708, signal_2250}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2236 ( .a ({signal_3677, signal_2219}), .b ({signal_3709, signal_2251}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2237 ( .a ({signal_3678, signal_2220}), .b ({signal_3710, signal_2252}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2238 ( .a ({signal_3679, signal_2221}), .b ({signal_3711, signal_2253}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2240 ( .a ({signal_3686, signal_2228}), .b ({signal_3713, signal_2255}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2242 ( .a ({signal_3694, signal_2236}), .b ({signal_3715, signal_2257}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2248 ( .a ({signal_3532, signal_2074}), .b ({signal_3658, signal_2200}), .clk ( clk ), .r ( Fresh[728] ), .c ({signal_3721, signal_2263}) ) ;
    buf_clk cell_3800 ( .C ( clk ), .D ( signal_6159 ), .Q ( signal_6160 ) ) ;
    buf_clk cell_3808 ( .C ( clk ), .D ( signal_6167 ), .Q ( signal_6168 ) ) ;
    buf_clk cell_3812 ( .C ( clk ), .D ( signal_6171 ), .Q ( signal_6172 ) ) ;
    buf_clk cell_3816 ( .C ( clk ), .D ( signal_6175 ), .Q ( signal_6176 ) ) ;
    buf_clk cell_3822 ( .C ( clk ), .D ( signal_6181 ), .Q ( signal_6182 ) ) ;
    buf_clk cell_3828 ( .C ( clk ), .D ( signal_6187 ), .Q ( signal_6188 ) ) ;
    buf_clk cell_3834 ( .C ( clk ), .D ( signal_6193 ), .Q ( signal_6194 ) ) ;
    buf_clk cell_3840 ( .C ( clk ), .D ( signal_6199 ), .Q ( signal_6200 ) ) ;
    buf_clk cell_3844 ( .C ( clk ), .D ( signal_6203 ), .Q ( signal_6204 ) ) ;
    buf_clk cell_3848 ( .C ( clk ), .D ( signal_6207 ), .Q ( signal_6208 ) ) ;
    buf_clk cell_3854 ( .C ( clk ), .D ( signal_6213 ), .Q ( signal_6214 ) ) ;
    buf_clk cell_3860 ( .C ( clk ), .D ( signal_6219 ), .Q ( signal_6220 ) ) ;
    buf_clk cell_3864 ( .C ( clk ), .D ( signal_6223 ), .Q ( signal_6224 ) ) ;
    buf_clk cell_3868 ( .C ( clk ), .D ( signal_6227 ), .Q ( signal_6228 ) ) ;
    buf_clk cell_3872 ( .C ( clk ), .D ( signal_6231 ), .Q ( signal_6232 ) ) ;
    buf_clk cell_3876 ( .C ( clk ), .D ( signal_6235 ), .Q ( signal_6236 ) ) ;
    buf_clk cell_3878 ( .C ( clk ), .D ( signal_6237 ), .Q ( signal_6238 ) ) ;
    buf_clk cell_3880 ( .C ( clk ), .D ( signal_6239 ), .Q ( signal_6240 ) ) ;
    buf_clk cell_3882 ( .C ( clk ), .D ( signal_6241 ), .Q ( signal_6242 ) ) ;
    buf_clk cell_3884 ( .C ( clk ), .D ( signal_6243 ), .Q ( signal_6244 ) ) ;
    buf_clk cell_3890 ( .C ( clk ), .D ( signal_6249 ), .Q ( signal_6250 ) ) ;
    buf_clk cell_3896 ( .C ( clk ), .D ( signal_6255 ), .Q ( signal_6256 ) ) ;
    buf_clk cell_3902 ( .C ( clk ), .D ( signal_6261 ), .Q ( signal_6262 ) ) ;
    buf_clk cell_3908 ( .C ( clk ), .D ( signal_6267 ), .Q ( signal_6268 ) ) ;
    buf_clk cell_3914 ( .C ( clk ), .D ( signal_6273 ), .Q ( signal_6274 ) ) ;
    buf_clk cell_3920 ( .C ( clk ), .D ( signal_6279 ), .Q ( signal_6280 ) ) ;
    buf_clk cell_3922 ( .C ( clk ), .D ( signal_6281 ), .Q ( signal_6282 ) ) ;
    buf_clk cell_3924 ( .C ( clk ), .D ( signal_6283 ), .Q ( signal_6284 ) ) ;
    buf_clk cell_3928 ( .C ( clk ), .D ( signal_6287 ), .Q ( signal_6288 ) ) ;
    buf_clk cell_3932 ( .C ( clk ), .D ( signal_6291 ), .Q ( signal_6292 ) ) ;
    buf_clk cell_3938 ( .C ( clk ), .D ( signal_6297 ), .Q ( signal_6298 ) ) ;
    buf_clk cell_3944 ( .C ( clk ), .D ( signal_6303 ), .Q ( signal_6304 ) ) ;
    buf_clk cell_3946 ( .C ( clk ), .D ( signal_6305 ), .Q ( signal_6306 ) ) ;
    buf_clk cell_3948 ( .C ( clk ), .D ( signal_6307 ), .Q ( signal_6308 ) ) ;
    buf_clk cell_3954 ( .C ( clk ), .D ( signal_6313 ), .Q ( signal_6314 ) ) ;
    buf_clk cell_3960 ( .C ( clk ), .D ( signal_6319 ), .Q ( signal_6320 ) ) ;
    buf_clk cell_3962 ( .C ( clk ), .D ( signal_6321 ), .Q ( signal_6322 ) ) ;
    buf_clk cell_3964 ( .C ( clk ), .D ( signal_6323 ), .Q ( signal_6324 ) ) ;
    buf_clk cell_3972 ( .C ( clk ), .D ( signal_6331 ), .Q ( signal_6332 ) ) ;
    buf_clk cell_3980 ( .C ( clk ), .D ( signal_6339 ), .Q ( signal_6340 ) ) ;
    buf_clk cell_3984 ( .C ( clk ), .D ( signal_6343 ), .Q ( signal_6344 ) ) ;
    buf_clk cell_3988 ( .C ( clk ), .D ( signal_6347 ), .Q ( signal_6348 ) ) ;
    buf_clk cell_3992 ( .C ( clk ), .D ( signal_6351 ), .Q ( signal_6352 ) ) ;
    buf_clk cell_3996 ( .C ( clk ), .D ( signal_6355 ), .Q ( signal_6356 ) ) ;
    buf_clk cell_4002 ( .C ( clk ), .D ( signal_6361 ), .Q ( signal_6362 ) ) ;
    buf_clk cell_4008 ( .C ( clk ), .D ( signal_6367 ), .Q ( signal_6368 ) ) ;
    buf_clk cell_4014 ( .C ( clk ), .D ( signal_6373 ), .Q ( signal_6374 ) ) ;
    buf_clk cell_4020 ( .C ( clk ), .D ( signal_6379 ), .Q ( signal_6380 ) ) ;
    buf_clk cell_4024 ( .C ( clk ), .D ( signal_6383 ), .Q ( signal_6384 ) ) ;
    buf_clk cell_4028 ( .C ( clk ), .D ( signal_6387 ), .Q ( signal_6388 ) ) ;
    buf_clk cell_4036 ( .C ( clk ), .D ( signal_6395 ), .Q ( signal_6396 ) ) ;
    buf_clk cell_4044 ( .C ( clk ), .D ( signal_6403 ), .Q ( signal_6404 ) ) ;
    buf_clk cell_4050 ( .C ( clk ), .D ( signal_6409 ), .Q ( signal_6410 ) ) ;
    buf_clk cell_4056 ( .C ( clk ), .D ( signal_6415 ), .Q ( signal_6416 ) ) ;
    buf_clk cell_4062 ( .C ( clk ), .D ( signal_6421 ), .Q ( signal_6422 ) ) ;
    buf_clk cell_4068 ( .C ( clk ), .D ( signal_6427 ), .Q ( signal_6428 ) ) ;
    buf_clk cell_4070 ( .C ( clk ), .D ( signal_6429 ), .Q ( signal_6430 ) ) ;
    buf_clk cell_4072 ( .C ( clk ), .D ( signal_6431 ), .Q ( signal_6432 ) ) ;
    buf_clk cell_4074 ( .C ( clk ), .D ( signal_6433 ), .Q ( signal_6434 ) ) ;
    buf_clk cell_4076 ( .C ( clk ), .D ( signal_6435 ), .Q ( signal_6436 ) ) ;
    buf_clk cell_4082 ( .C ( clk ), .D ( signal_6441 ), .Q ( signal_6442 ) ) ;
    buf_clk cell_4088 ( .C ( clk ), .D ( signal_6447 ), .Q ( signal_6448 ) ) ;
    buf_clk cell_4090 ( .C ( clk ), .D ( signal_6449 ), .Q ( signal_6450 ) ) ;
    buf_clk cell_4092 ( .C ( clk ), .D ( signal_6451 ), .Q ( signal_6452 ) ) ;
    buf_clk cell_4094 ( .C ( clk ), .D ( signal_6453 ), .Q ( signal_6454 ) ) ;
    buf_clk cell_4096 ( .C ( clk ), .D ( signal_6455 ), .Q ( signal_6456 ) ) ;
    buf_clk cell_4102 ( .C ( clk ), .D ( signal_6461 ), .Q ( signal_6462 ) ) ;
    buf_clk cell_4108 ( .C ( clk ), .D ( signal_6467 ), .Q ( signal_6468 ) ) ;
    buf_clk cell_4114 ( .C ( clk ), .D ( signal_6473 ), .Q ( signal_6474 ) ) ;
    buf_clk cell_4120 ( .C ( clk ), .D ( signal_6479 ), .Q ( signal_6480 ) ) ;
    buf_clk cell_4124 ( .C ( clk ), .D ( signal_6483 ), .Q ( signal_6484 ) ) ;
    buf_clk cell_4128 ( .C ( clk ), .D ( signal_6487 ), .Q ( signal_6488 ) ) ;
    buf_clk cell_4136 ( .C ( clk ), .D ( signal_6495 ), .Q ( signal_6496 ) ) ;
    buf_clk cell_4146 ( .C ( clk ), .D ( signal_6505 ), .Q ( signal_6506 ) ) ;
    buf_clk cell_4152 ( .C ( clk ), .D ( signal_6511 ), .Q ( signal_6512 ) ) ;
    buf_clk cell_4158 ( .C ( clk ), .D ( signal_6517 ), .Q ( signal_6518 ) ) ;
    buf_clk cell_4166 ( .C ( clk ), .D ( signal_6525 ), .Q ( signal_6526 ) ) ;
    buf_clk cell_4174 ( .C ( clk ), .D ( signal_6533 ), .Q ( signal_6534 ) ) ;
    buf_clk cell_4182 ( .C ( clk ), .D ( signal_6541 ), .Q ( signal_6542 ) ) ;
    buf_clk cell_4190 ( .C ( clk ), .D ( signal_6549 ), .Q ( signal_6550 ) ) ;
    buf_clk cell_4194 ( .C ( clk ), .D ( signal_6553 ), .Q ( signal_6554 ) ) ;
    buf_clk cell_4198 ( .C ( clk ), .D ( signal_6557 ), .Q ( signal_6558 ) ) ;
    buf_clk cell_4202 ( .C ( clk ), .D ( signal_6561 ), .Q ( signal_6562 ) ) ;
    buf_clk cell_4206 ( .C ( clk ), .D ( signal_6565 ), .Q ( signal_6566 ) ) ;
    buf_clk cell_4218 ( .C ( clk ), .D ( signal_6577 ), .Q ( signal_6578 ) ) ;
    buf_clk cell_4222 ( .C ( clk ), .D ( signal_6581 ), .Q ( signal_6582 ) ) ;
    buf_clk cell_4232 ( .C ( clk ), .D ( signal_6591 ), .Q ( signal_6592 ) ) ;
    buf_clk cell_4242 ( .C ( clk ), .D ( signal_6601 ), .Q ( signal_6602 ) ) ;
    buf_clk cell_4248 ( .C ( clk ), .D ( signal_6607 ), .Q ( signal_6608 ) ) ;
    buf_clk cell_4254 ( .C ( clk ), .D ( signal_6613 ), .Q ( signal_6614 ) ) ;
    buf_clk cell_4266 ( .C ( clk ), .D ( signal_6625 ), .Q ( signal_6626 ) ) ;
    buf_clk cell_4274 ( .C ( clk ), .D ( signal_6633 ), .Q ( signal_6634 ) ) ;
    buf_clk cell_4280 ( .C ( clk ), .D ( signal_6639 ), .Q ( signal_6640 ) ) ;
    buf_clk cell_4286 ( .C ( clk ), .D ( signal_6645 ), .Q ( signal_6646 ) ) ;
    buf_clk cell_4294 ( .C ( clk ), .D ( signal_6653 ), .Q ( signal_6654 ) ) ;
    buf_clk cell_4302 ( .C ( clk ), .D ( signal_6661 ), .Q ( signal_6662 ) ) ;
    buf_clk cell_4310 ( .C ( clk ), .D ( signal_6669 ), .Q ( signal_6670 ) ) ;
    buf_clk cell_4318 ( .C ( clk ), .D ( signal_6677 ), .Q ( signal_6678 ) ) ;
    buf_clk cell_4326 ( .C ( clk ), .D ( signal_6685 ), .Q ( signal_6686 ) ) ;
    buf_clk cell_4334 ( .C ( clk ), .D ( signal_6693 ), .Q ( signal_6694 ) ) ;
    buf_clk cell_4344 ( .C ( clk ), .D ( signal_6703 ), .Q ( signal_6704 ) ) ;
    buf_clk cell_4354 ( .C ( clk ), .D ( signal_6713 ), .Q ( signal_6714 ) ) ;
    buf_clk cell_4362 ( .C ( clk ), .D ( signal_6721 ), .Q ( signal_6722 ) ) ;
    buf_clk cell_4370 ( .C ( clk ), .D ( signal_6729 ), .Q ( signal_6730 ) ) ;
    buf_clk cell_4378 ( .C ( clk ), .D ( signal_6737 ), .Q ( signal_6738 ) ) ;
    buf_clk cell_4386 ( .C ( clk ), .D ( signal_6745 ), .Q ( signal_6746 ) ) ;
    buf_clk cell_4398 ( .C ( clk ), .D ( signal_6757 ), .Q ( signal_6758 ) ) ;
    buf_clk cell_4406 ( .C ( clk ), .D ( signal_6765 ), .Q ( signal_6766 ) ) ;
    buf_clk cell_4414 ( .C ( clk ), .D ( signal_6773 ), .Q ( signal_6774 ) ) ;
    buf_clk cell_4422 ( .C ( clk ), .D ( signal_6781 ), .Q ( signal_6782 ) ) ;
    buf_clk cell_4430 ( .C ( clk ), .D ( signal_6789 ), .Q ( signal_6790 ) ) ;
    buf_clk cell_4438 ( .C ( clk ), .D ( signal_6797 ), .Q ( signal_6798 ) ) ;
    buf_clk cell_4442 ( .C ( clk ), .D ( signal_6801 ), .Q ( signal_6802 ) ) ;
    buf_clk cell_4448 ( .C ( clk ), .D ( signal_6807 ), .Q ( signal_6808 ) ) ;
    buf_clk cell_4456 ( .C ( clk ), .D ( signal_6815 ), .Q ( signal_6816 ) ) ;
    buf_clk cell_4464 ( .C ( clk ), .D ( signal_6823 ), .Q ( signal_6824 ) ) ;
    buf_clk cell_4470 ( .C ( clk ), .D ( signal_6829 ), .Q ( signal_6830 ) ) ;
    buf_clk cell_4476 ( .C ( clk ), .D ( signal_6835 ), .Q ( signal_6836 ) ) ;
    buf_clk cell_4482 ( .C ( clk ), .D ( signal_6841 ), .Q ( signal_6842 ) ) ;
    buf_clk cell_4488 ( .C ( clk ), .D ( signal_6847 ), .Q ( signal_6848 ) ) ;
    buf_clk cell_4496 ( .C ( clk ), .D ( signal_6855 ), .Q ( signal_6856 ) ) ;
    buf_clk cell_4504 ( .C ( clk ), .D ( signal_6863 ), .Q ( signal_6864 ) ) ;
    buf_clk cell_4514 ( .C ( clk ), .D ( signal_6873 ), .Q ( signal_6874 ) ) ;
    buf_clk cell_4524 ( .C ( clk ), .D ( signal_6883 ), .Q ( signal_6884 ) ) ;
    buf_clk cell_4534 ( .C ( clk ), .D ( signal_6893 ), .Q ( signal_6894 ) ) ;
    buf_clk cell_4540 ( .C ( clk ), .D ( signal_6899 ), .Q ( signal_6900 ) ) ;
    buf_clk cell_4548 ( .C ( clk ), .D ( signal_6907 ), .Q ( signal_6908 ) ) ;
    buf_clk cell_4556 ( .C ( clk ), .D ( signal_6915 ), .Q ( signal_6916 ) ) ;
    buf_clk cell_4566 ( .C ( clk ), .D ( signal_6925 ), .Q ( signal_6926 ) ) ;
    buf_clk cell_4576 ( .C ( clk ), .D ( signal_6935 ), .Q ( signal_6936 ) ) ;
    buf_clk cell_4584 ( .C ( clk ), .D ( signal_6943 ), .Q ( signal_6944 ) ) ;
    buf_clk cell_4592 ( .C ( clk ), .D ( signal_6951 ), .Q ( signal_6952 ) ) ;
    buf_clk cell_4598 ( .C ( clk ), .D ( signal_6957 ), .Q ( signal_6958 ) ) ;
    buf_clk cell_4604 ( .C ( clk ), .D ( signal_6963 ), .Q ( signal_6964 ) ) ;
    buf_clk cell_4610 ( .C ( clk ), .D ( signal_6969 ), .Q ( signal_6970 ) ) ;
    buf_clk cell_4616 ( .C ( clk ), .D ( signal_6975 ), .Q ( signal_6976 ) ) ;
    buf_clk cell_4642 ( .C ( clk ), .D ( signal_7001 ), .Q ( signal_7002 ) ) ;
    buf_clk cell_4648 ( .C ( clk ), .D ( signal_7007 ), .Q ( signal_7008 ) ) ;
    buf_clk cell_4658 ( .C ( clk ), .D ( signal_7017 ), .Q ( signal_7018 ) ) ;
    buf_clk cell_4664 ( .C ( clk ), .D ( signal_7023 ), .Q ( signal_7024 ) ) ;
    buf_clk cell_4678 ( .C ( clk ), .D ( signal_7037 ), .Q ( signal_7038 ) ) ;
    buf_clk cell_4684 ( .C ( clk ), .D ( signal_7043 ), .Q ( signal_7044 ) ) ;
    buf_clk cell_4714 ( .C ( clk ), .D ( signal_7073 ), .Q ( signal_7074 ) ) ;
    buf_clk cell_4722 ( .C ( clk ), .D ( signal_7081 ), .Q ( signal_7082 ) ) ;
    buf_clk cell_4744 ( .C ( clk ), .D ( signal_7103 ), .Q ( signal_7104 ) ) ;
    buf_clk cell_4754 ( .C ( clk ), .D ( signal_7113 ), .Q ( signal_7114 ) ) ;
    buf_clk cell_4782 ( .C ( clk ), .D ( signal_7141 ), .Q ( signal_7142 ) ) ;
    buf_clk cell_4790 ( .C ( clk ), .D ( signal_7149 ), .Q ( signal_7150 ) ) ;
    buf_clk cell_4810 ( .C ( clk ), .D ( signal_7169 ), .Q ( signal_7170 ) ) ;
    buf_clk cell_4818 ( .C ( clk ), .D ( signal_7177 ), .Q ( signal_7178 ) ) ;
    buf_clk cell_4838 ( .C ( clk ), .D ( signal_7197 ), .Q ( signal_7198 ) ) ;
    buf_clk cell_4846 ( .C ( clk ), .D ( signal_7205 ), .Q ( signal_7206 ) ) ;
    buf_clk cell_4920 ( .C ( clk ), .D ( signal_7279 ), .Q ( signal_7280 ) ) ;
    buf_clk cell_4932 ( .C ( clk ), .D ( signal_7291 ), .Q ( signal_7292 ) ) ;
    buf_clk cell_4970 ( .C ( clk ), .D ( signal_7329 ), .Q ( signal_7330 ) ) ;
    buf_clk cell_4984 ( .C ( clk ), .D ( signal_7343 ), .Q ( signal_7344 ) ) ;
    buf_clk cell_5014 ( .C ( clk ), .D ( signal_7373 ), .Q ( signal_7374 ) ) ;
    buf_clk cell_5028 ( .C ( clk ), .D ( signal_7387 ), .Q ( signal_7388 ) ) ;
    buf_clk cell_5094 ( .C ( clk ), .D ( signal_7453 ), .Q ( signal_7454 ) ) ;
    buf_clk cell_5110 ( .C ( clk ), .D ( signal_7469 ), .Q ( signal_7470 ) ) ;
    buf_clk cell_5134 ( .C ( clk ), .D ( signal_7493 ), .Q ( signal_7494 ) ) ;
    buf_clk cell_5150 ( .C ( clk ), .D ( signal_7509 ), .Q ( signal_7510 ) ) ;
    buf_clk cell_5256 ( .C ( clk ), .D ( signal_7615 ), .Q ( signal_7616 ) ) ;
    buf_clk cell_5272 ( .C ( clk ), .D ( signal_7631 ), .Q ( signal_7632 ) ) ;
    buf_clk cell_5290 ( .C ( clk ), .D ( signal_7649 ), .Q ( signal_7650 ) ) ;
    buf_clk cell_5308 ( .C ( clk ), .D ( signal_7667 ), .Q ( signal_7668 ) ) ;
    buf_clk cell_5390 ( .C ( clk ), .D ( signal_7749 ), .Q ( signal_7750 ) ) ;
    buf_clk cell_5410 ( .C ( clk ), .D ( signal_7769 ), .Q ( signal_7770 ) ) ;

    /* cells in depth 13 */
    buf_clk cell_4137 ( .C ( clk ), .D ( signal_6496 ), .Q ( signal_6497 ) ) ;
    buf_clk cell_4147 ( .C ( clk ), .D ( signal_6506 ), .Q ( signal_6507 ) ) ;
    buf_clk cell_4153 ( .C ( clk ), .D ( signal_6512 ), .Q ( signal_6513 ) ) ;
    buf_clk cell_4159 ( .C ( clk ), .D ( signal_6518 ), .Q ( signal_6519 ) ) ;
    buf_clk cell_4167 ( .C ( clk ), .D ( signal_6526 ), .Q ( signal_6527 ) ) ;
    buf_clk cell_4175 ( .C ( clk ), .D ( signal_6534 ), .Q ( signal_6535 ) ) ;
    buf_clk cell_4183 ( .C ( clk ), .D ( signal_6542 ), .Q ( signal_6543 ) ) ;
    buf_clk cell_4191 ( .C ( clk ), .D ( signal_6550 ), .Q ( signal_6551 ) ) ;
    buf_clk cell_4195 ( .C ( clk ), .D ( signal_6554 ), .Q ( signal_6555 ) ) ;
    buf_clk cell_4199 ( .C ( clk ), .D ( signal_6558 ), .Q ( signal_6559 ) ) ;
    buf_clk cell_4203 ( .C ( clk ), .D ( signal_6562 ), .Q ( signal_6563 ) ) ;
    buf_clk cell_4207 ( .C ( clk ), .D ( signal_6566 ), .Q ( signal_6567 ) ) ;
    buf_clk cell_4209 ( .C ( clk ), .D ( signal_6454 ), .Q ( signal_6569 ) ) ;
    buf_clk cell_4211 ( .C ( clk ), .D ( signal_6456 ), .Q ( signal_6571 ) ) ;
    buf_clk cell_4213 ( .C ( clk ), .D ( signal_2156 ), .Q ( signal_6573 ) ) ;
    buf_clk cell_4215 ( .C ( clk ), .D ( signal_3614 ), .Q ( signal_6575 ) ) ;
    buf_clk cell_4219 ( .C ( clk ), .D ( signal_6578 ), .Q ( signal_6579 ) ) ;
    buf_clk cell_4223 ( .C ( clk ), .D ( signal_6582 ), .Q ( signal_6583 ) ) ;
    buf_clk cell_4233 ( .C ( clk ), .D ( signal_6592 ), .Q ( signal_6593 ) ) ;
    buf_clk cell_4243 ( .C ( clk ), .D ( signal_6602 ), .Q ( signal_6603 ) ) ;
    buf_clk cell_4249 ( .C ( clk ), .D ( signal_6608 ), .Q ( signal_6609 ) ) ;
    buf_clk cell_4255 ( .C ( clk ), .D ( signal_6614 ), .Q ( signal_6615 ) ) ;
    buf_clk cell_4257 ( .C ( clk ), .D ( signal_6288 ), .Q ( signal_6617 ) ) ;
    buf_clk cell_4259 ( .C ( clk ), .D ( signal_6292 ), .Q ( signal_6619 ) ) ;
    buf_clk cell_4267 ( .C ( clk ), .D ( signal_6626 ), .Q ( signal_6627 ) ) ;
    buf_clk cell_4275 ( .C ( clk ), .D ( signal_6634 ), .Q ( signal_6635 ) ) ;
    buf_clk cell_4281 ( .C ( clk ), .D ( signal_6640 ), .Q ( signal_6641 ) ) ;
    buf_clk cell_4287 ( .C ( clk ), .D ( signal_6646 ), .Q ( signal_6647 ) ) ;
    buf_clk cell_4295 ( .C ( clk ), .D ( signal_6654 ), .Q ( signal_6655 ) ) ;
    buf_clk cell_4303 ( .C ( clk ), .D ( signal_6662 ), .Q ( signal_6663 ) ) ;
    buf_clk cell_4311 ( .C ( clk ), .D ( signal_6670 ), .Q ( signal_6671 ) ) ;
    buf_clk cell_4319 ( .C ( clk ), .D ( signal_6678 ), .Q ( signal_6679 ) ) ;
    buf_clk cell_4327 ( .C ( clk ), .D ( signal_6686 ), .Q ( signal_6687 ) ) ;
    buf_clk cell_4335 ( .C ( clk ), .D ( signal_6694 ), .Q ( signal_6695 ) ) ;
    buf_clk cell_4345 ( .C ( clk ), .D ( signal_6704 ), .Q ( signal_6705 ) ) ;
    buf_clk cell_4355 ( .C ( clk ), .D ( signal_6714 ), .Q ( signal_6715 ) ) ;
    buf_clk cell_4363 ( .C ( clk ), .D ( signal_6722 ), .Q ( signal_6723 ) ) ;
    buf_clk cell_4371 ( .C ( clk ), .D ( signal_6730 ), .Q ( signal_6731 ) ) ;
    buf_clk cell_4379 ( .C ( clk ), .D ( signal_6738 ), .Q ( signal_6739 ) ) ;
    buf_clk cell_4387 ( .C ( clk ), .D ( signal_6746 ), .Q ( signal_6747 ) ) ;
    buf_clk cell_4389 ( .C ( clk ), .D ( signal_6242 ), .Q ( signal_6749 ) ) ;
    buf_clk cell_4391 ( .C ( clk ), .D ( signal_6244 ), .Q ( signal_6751 ) ) ;
    buf_clk cell_4399 ( .C ( clk ), .D ( signal_6758 ), .Q ( signal_6759 ) ) ;
    buf_clk cell_4407 ( .C ( clk ), .D ( signal_6766 ), .Q ( signal_6767 ) ) ;
    buf_clk cell_4415 ( .C ( clk ), .D ( signal_6774 ), .Q ( signal_6775 ) ) ;
    buf_clk cell_4423 ( .C ( clk ), .D ( signal_6782 ), .Q ( signal_6783 ) ) ;
    buf_clk cell_4431 ( .C ( clk ), .D ( signal_6790 ), .Q ( signal_6791 ) ) ;
    buf_clk cell_4439 ( .C ( clk ), .D ( signal_6798 ), .Q ( signal_6799 ) ) ;
    buf_clk cell_4443 ( .C ( clk ), .D ( signal_6802 ), .Q ( signal_6803 ) ) ;
    buf_clk cell_4449 ( .C ( clk ), .D ( signal_6808 ), .Q ( signal_6809 ) ) ;
    buf_clk cell_4457 ( .C ( clk ), .D ( signal_6816 ), .Q ( signal_6817 ) ) ;
    buf_clk cell_4465 ( .C ( clk ), .D ( signal_6824 ), .Q ( signal_6825 ) ) ;
    buf_clk cell_4471 ( .C ( clk ), .D ( signal_6830 ), .Q ( signal_6831 ) ) ;
    buf_clk cell_4477 ( .C ( clk ), .D ( signal_6836 ), .Q ( signal_6837 ) ) ;
    buf_clk cell_4483 ( .C ( clk ), .D ( signal_6842 ), .Q ( signal_6843 ) ) ;
    buf_clk cell_4489 ( .C ( clk ), .D ( signal_6848 ), .Q ( signal_6849 ) ) ;
    buf_clk cell_4497 ( .C ( clk ), .D ( signal_6856 ), .Q ( signal_6857 ) ) ;
    buf_clk cell_4505 ( .C ( clk ), .D ( signal_6864 ), .Q ( signal_6865 ) ) ;
    buf_clk cell_4515 ( .C ( clk ), .D ( signal_6874 ), .Q ( signal_6875 ) ) ;
    buf_clk cell_4525 ( .C ( clk ), .D ( signal_6884 ), .Q ( signal_6885 ) ) ;
    buf_clk cell_4535 ( .C ( clk ), .D ( signal_6894 ), .Q ( signal_6895 ) ) ;
    buf_clk cell_4541 ( .C ( clk ), .D ( signal_6900 ), .Q ( signal_6901 ) ) ;
    buf_clk cell_4549 ( .C ( clk ), .D ( signal_6908 ), .Q ( signal_6909 ) ) ;
    buf_clk cell_4557 ( .C ( clk ), .D ( signal_6916 ), .Q ( signal_6917 ) ) ;
    buf_clk cell_4567 ( .C ( clk ), .D ( signal_6926 ), .Q ( signal_6927 ) ) ;
    buf_clk cell_4577 ( .C ( clk ), .D ( signal_6936 ), .Q ( signal_6937 ) ) ;
    buf_clk cell_4585 ( .C ( clk ), .D ( signal_6944 ), .Q ( signal_6945 ) ) ;
    buf_clk cell_4593 ( .C ( clk ), .D ( signal_6952 ), .Q ( signal_6953 ) ) ;
    buf_clk cell_4599 ( .C ( clk ), .D ( signal_6958 ), .Q ( signal_6959 ) ) ;
    buf_clk cell_4605 ( .C ( clk ), .D ( signal_6964 ), .Q ( signal_6965 ) ) ;
    buf_clk cell_4611 ( .C ( clk ), .D ( signal_6970 ), .Q ( signal_6971 ) ) ;
    buf_clk cell_4617 ( .C ( clk ), .D ( signal_6976 ), .Q ( signal_6977 ) ) ;
    buf_clk cell_4625 ( .C ( clk ), .D ( signal_6422 ), .Q ( signal_6985 ) ) ;
    buf_clk cell_4629 ( .C ( clk ), .D ( signal_6428 ), .Q ( signal_6989 ) ) ;
    buf_clk cell_4633 ( .C ( clk ), .D ( signal_2253 ), .Q ( signal_6993 ) ) ;
    buf_clk cell_4637 ( .C ( clk ), .D ( signal_3711 ), .Q ( signal_6997 ) ) ;
    buf_clk cell_4643 ( .C ( clk ), .D ( signal_7002 ), .Q ( signal_7003 ) ) ;
    buf_clk cell_4649 ( .C ( clk ), .D ( signal_7008 ), .Q ( signal_7009 ) ) ;
    buf_clk cell_4659 ( .C ( clk ), .D ( signal_7018 ), .Q ( signal_7019 ) ) ;
    buf_clk cell_4665 ( .C ( clk ), .D ( signal_7024 ), .Q ( signal_7025 ) ) ;
    buf_clk cell_4669 ( .C ( clk ), .D ( signal_2208 ), .Q ( signal_7029 ) ) ;
    buf_clk cell_4673 ( .C ( clk ), .D ( signal_3666 ), .Q ( signal_7033 ) ) ;
    buf_clk cell_4679 ( .C ( clk ), .D ( signal_7038 ), .Q ( signal_7039 ) ) ;
    buf_clk cell_4685 ( .C ( clk ), .D ( signal_7044 ), .Q ( signal_7045 ) ) ;
    buf_clk cell_4693 ( .C ( clk ), .D ( signal_2249 ), .Q ( signal_7053 ) ) ;
    buf_clk cell_4697 ( .C ( clk ), .D ( signal_3707 ), .Q ( signal_7057 ) ) ;
    buf_clk cell_4701 ( .C ( clk ), .D ( signal_2161 ), .Q ( signal_7061 ) ) ;
    buf_clk cell_4707 ( .C ( clk ), .D ( signal_3619 ), .Q ( signal_7067 ) ) ;
    buf_clk cell_4715 ( .C ( clk ), .D ( signal_7074 ), .Q ( signal_7075 ) ) ;
    buf_clk cell_4723 ( .C ( clk ), .D ( signal_7082 ), .Q ( signal_7083 ) ) ;
    buf_clk cell_4729 ( .C ( clk ), .D ( signal_2199 ), .Q ( signal_7089 ) ) ;
    buf_clk cell_4735 ( .C ( clk ), .D ( signal_3657 ), .Q ( signal_7095 ) ) ;
    buf_clk cell_4745 ( .C ( clk ), .D ( signal_7104 ), .Q ( signal_7105 ) ) ;
    buf_clk cell_4755 ( .C ( clk ), .D ( signal_7114 ), .Q ( signal_7115 ) ) ;
    buf_clk cell_4761 ( .C ( clk ), .D ( signal_2255 ), .Q ( signal_7121 ) ) ;
    buf_clk cell_4767 ( .C ( clk ), .D ( signal_3713 ), .Q ( signal_7127 ) ) ;
    buf_clk cell_4783 ( .C ( clk ), .D ( signal_7142 ), .Q ( signal_7143 ) ) ;
    buf_clk cell_4791 ( .C ( clk ), .D ( signal_7150 ), .Q ( signal_7151 ) ) ;
    buf_clk cell_4797 ( .C ( clk ), .D ( signal_2183 ), .Q ( signal_7157 ) ) ;
    buf_clk cell_4803 ( .C ( clk ), .D ( signal_3641 ), .Q ( signal_7163 ) ) ;
    buf_clk cell_4811 ( .C ( clk ), .D ( signal_7170 ), .Q ( signal_7171 ) ) ;
    buf_clk cell_4819 ( .C ( clk ), .D ( signal_7178 ), .Q ( signal_7179 ) ) ;
    buf_clk cell_4825 ( .C ( clk ), .D ( signal_6450 ), .Q ( signal_7185 ) ) ;
    buf_clk cell_4831 ( .C ( clk ), .D ( signal_6452 ), .Q ( signal_7191 ) ) ;
    buf_clk cell_4839 ( .C ( clk ), .D ( signal_7198 ), .Q ( signal_7199 ) ) ;
    buf_clk cell_4847 ( .C ( clk ), .D ( signal_7206 ), .Q ( signal_7207 ) ) ;
    buf_clk cell_4861 ( .C ( clk ), .D ( signal_2252 ), .Q ( signal_7221 ) ) ;
    buf_clk cell_4867 ( .C ( clk ), .D ( signal_3710 ), .Q ( signal_7227 ) ) ;
    buf_clk cell_4873 ( .C ( clk ), .D ( signal_2160 ), .Q ( signal_7233 ) ) ;
    buf_clk cell_4879 ( .C ( clk ), .D ( signal_3618 ), .Q ( signal_7239 ) ) ;
    buf_clk cell_4901 ( .C ( clk ), .D ( signal_2202 ), .Q ( signal_7261 ) ) ;
    buf_clk cell_4909 ( .C ( clk ), .D ( signal_3660 ), .Q ( signal_7269 ) ) ;
    buf_clk cell_4921 ( .C ( clk ), .D ( signal_7280 ), .Q ( signal_7281 ) ) ;
    buf_clk cell_4933 ( .C ( clk ), .D ( signal_7292 ), .Q ( signal_7293 ) ) ;
    buf_clk cell_4971 ( .C ( clk ), .D ( signal_7330 ), .Q ( signal_7331 ) ) ;
    buf_clk cell_4985 ( .C ( clk ), .D ( signal_7344 ), .Q ( signal_7345 ) ) ;
    buf_clk cell_4993 ( .C ( clk ), .D ( signal_2154 ), .Q ( signal_7353 ) ) ;
    buf_clk cell_5001 ( .C ( clk ), .D ( signal_3612 ), .Q ( signal_7361 ) ) ;
    buf_clk cell_5015 ( .C ( clk ), .D ( signal_7374 ), .Q ( signal_7375 ) ) ;
    buf_clk cell_5029 ( .C ( clk ), .D ( signal_7388 ), .Q ( signal_7389 ) ) ;
    buf_clk cell_5037 ( .C ( clk ), .D ( signal_2149 ), .Q ( signal_7397 ) ) ;
    buf_clk cell_5045 ( .C ( clk ), .D ( signal_3607 ), .Q ( signal_7405 ) ) ;
    buf_clk cell_5061 ( .C ( clk ), .D ( signal_2152 ), .Q ( signal_7421 ) ) ;
    buf_clk cell_5071 ( .C ( clk ), .D ( signal_3610 ), .Q ( signal_7431 ) ) ;
    buf_clk cell_5095 ( .C ( clk ), .D ( signal_7454 ), .Q ( signal_7455 ) ) ;
    buf_clk cell_5111 ( .C ( clk ), .D ( signal_7470 ), .Q ( signal_7471 ) ) ;
    buf_clk cell_5135 ( .C ( clk ), .D ( signal_7494 ), .Q ( signal_7495 ) ) ;
    buf_clk cell_5151 ( .C ( clk ), .D ( signal_7510 ), .Q ( signal_7511 ) ) ;
    buf_clk cell_5161 ( .C ( clk ), .D ( signal_2257 ), .Q ( signal_7521 ) ) ;
    buf_clk cell_5171 ( .C ( clk ), .D ( signal_3715 ), .Q ( signal_7531 ) ) ;
    buf_clk cell_5257 ( .C ( clk ), .D ( signal_7616 ), .Q ( signal_7617 ) ) ;
    buf_clk cell_5273 ( .C ( clk ), .D ( signal_7632 ), .Q ( signal_7633 ) ) ;
    buf_clk cell_5291 ( .C ( clk ), .D ( signal_7650 ), .Q ( signal_7651 ) ) ;
    buf_clk cell_5309 ( .C ( clk ), .D ( signal_7668 ), .Q ( signal_7669 ) ) ;
    buf_clk cell_5391 ( .C ( clk ), .D ( signal_7750 ), .Q ( signal_7751 ) ) ;
    buf_clk cell_5411 ( .C ( clk ), .D ( signal_7770 ), .Q ( signal_7771 ) ) ;

    /* cells in depth 14 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2116 ( .a ({signal_6168, signal_6160}), .b ({signal_3511, signal_2053}), .clk ( clk ), .r ( Fresh[729] ), .c ({signal_3589, signal_2131}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2118 ( .a ({signal_6176, signal_6172}), .b ({signal_3512, signal_2054}), .clk ( clk ), .r ( Fresh[730] ), .c ({signal_3591, signal_2133}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2119 ( .a ({signal_6188, signal_6182}), .b ({signal_3513, signal_2055}), .clk ( clk ), .r ( Fresh[731] ), .c ({signal_3592, signal_2134}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2121 ( .a ({signal_6200, signal_6194}), .b ({signal_3515, signal_2057}), .clk ( clk ), .r ( Fresh[732] ), .c ({signal_3594, signal_2136}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2122 ( .a ({signal_6208, signal_6204}), .b ({signal_3517, signal_2059}), .clk ( clk ), .r ( Fresh[733] ), .c ({signal_3595, signal_2137}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2123 ( .a ({signal_6220, signal_6214}), .b ({signal_3518, signal_2060}), .clk ( clk ), .r ( Fresh[734] ), .c ({signal_3596, signal_2138}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2140 ( .a ({signal_3592, signal_2134}), .b ({signal_3613, signal_2155}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2162 ( .a ({signal_6228, signal_6224}), .b ({signal_3537, signal_2079}), .clk ( clk ), .r ( Fresh[735] ), .c ({signal_3635, signal_2177}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2170 ( .a ({signal_6236, signal_6232}), .b ({signal_3571, signal_2113}), .clk ( clk ), .r ( Fresh[736] ), .c ({signal_3643, signal_2185}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2172 ( .a ({signal_6240, signal_6238}), .b ({signal_3575, signal_2117}), .clk ( clk ), .r ( Fresh[737] ), .c ({signal_3645, signal_2187}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2173 ( .a ({signal_6244, signal_6242}), .b ({signal_3545, signal_2087}), .clk ( clk ), .r ( Fresh[738] ), .c ({signal_3646, signal_2188}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2174 ( .a ({signal_6256, signal_6250}), .b ({signal_3579, signal_2121}), .clk ( clk ), .r ( Fresh[739] ), .c ({signal_3647, signal_2189}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2175 ( .a ({signal_6268, signal_6262}), .b ({signal_3580, signal_2122}), .clk ( clk ), .r ( Fresh[740] ), .c ({signal_3648, signal_2190}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2176 ( .a ({signal_6280, signal_6274}), .b ({signal_3581, signal_2123}), .clk ( clk ), .r ( Fresh[741] ), .c ({signal_3649, signal_2191}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2177 ( .a ({signal_3541, signal_2083}), .b ({signal_3514, signal_2056}), .clk ( clk ), .r ( Fresh[742] ), .c ({signal_3650, signal_2192}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2178 ( .a ({signal_6284, signal_6282}), .b ({signal_3546, signal_2088}), .clk ( clk ), .r ( Fresh[743] ), .c ({signal_3651, signal_2193}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2179 ( .a ({signal_6292, signal_6288}), .b ({signal_3586, signal_2128}), .clk ( clk ), .r ( Fresh[744] ), .c ({signal_3652, signal_2194}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2190 ( .a ({signal_3635, signal_2177}), .b ({signal_3663, signal_2205}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2195 ( .a ({signal_3646, signal_2188}), .b ({signal_3668, signal_2210}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2196 ( .a ({signal_3648, signal_2190}), .b ({signal_3669, signal_2211}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2197 ( .a ({signal_3649, signal_2191}), .b ({signal_3670, signal_2212}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2198 ( .a ({signal_3651, signal_2193}), .b ({signal_3671, signal_2213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2200 ( .a ({signal_6304, signal_6298}), .b ({signal_3615, signal_2157}), .clk ( clk ), .r ( Fresh[745] ), .c ({signal_3673, signal_2215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2207 ( .a ({signal_6308, signal_6306}), .b ({signal_3604, signal_2146}), .clk ( clk ), .r ( Fresh[746] ), .c ({signal_3680, signal_2222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2208 ( .a ({signal_6320, signal_6314}), .b ({signal_3622, signal_2164}), .clk ( clk ), .r ( Fresh[747] ), .c ({signal_3681, signal_2223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2209 ( .a ({signal_6324, signal_6322}), .b ({signal_3605, signal_2147}), .clk ( clk ), .r ( Fresh[748] ), .c ({signal_3682, signal_2224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2210 ( .a ({signal_6340, signal_6332}), .b ({signal_3623, signal_2165}), .clk ( clk ), .r ( Fresh[749] ), .c ({signal_3683, signal_2225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2211 ( .a ({signal_6348, signal_6344}), .b ({signal_3625, signal_2167}), .clk ( clk ), .r ( Fresh[750] ), .c ({signal_3684, signal_2226}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2212 ( .a ({signal_3576, signal_2118}), .b ({signal_3626, signal_2168}), .clk ( clk ), .r ( Fresh[751] ), .c ({signal_3685, signal_2227}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2214 ( .a ({signal_6356, signal_6352}), .b ({signal_3627, signal_2169}), .clk ( clk ), .r ( Fresh[752] ), .c ({signal_3687, signal_2229}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2215 ( .a ({signal_3578, signal_2120}), .b ({signal_3628, signal_2170}), .clk ( clk ), .r ( Fresh[753] ), .c ({signal_3688, signal_2230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2216 ( .a ({signal_6368, signal_6362}), .b ({signal_3629, signal_2171}), .clk ( clk ), .r ( Fresh[754] ), .c ({signal_3689, signal_2231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2217 ( .a ({signal_6380, signal_6374}), .b ({signal_3631, signal_2173}), .clk ( clk ), .r ( Fresh[755] ), .c ({signal_3690, signal_2232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2218 ( .a ({signal_6388, signal_6384}), .b ({signal_3633, signal_2175}), .clk ( clk ), .r ( Fresh[756] ), .c ({signal_3691, signal_2233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2219 ( .a ({signal_6404, signal_6396}), .b ({signal_3634, signal_2176}), .clk ( clk ), .r ( Fresh[757] ), .c ({signal_3692, signal_2234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2220 ( .a ({signal_6416, signal_6410}), .b ({signal_3636, signal_2178}), .clk ( clk ), .r ( Fresh[758] ), .c ({signal_3693, signal_2235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2222 ( .a ({signal_3609, signal_2151}), .b ({signal_3585, signal_2127}), .clk ( clk ), .r ( Fresh[759] ), .c ({signal_3695, signal_2237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2223 ( .a ({signal_3611, signal_2153}), .b ({signal_3640, signal_2182}), .clk ( clk ), .r ( Fresh[760] ), .c ({signal_3696, signal_2238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2224 ( .a ({signal_6428, signal_6422}), .b ({signal_3642, signal_2184}), .clk ( clk ), .r ( Fresh[761] ), .c ({signal_3697, signal_2239}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2239 ( .a ({signal_3681, signal_2223}), .b ({signal_3712, signal_2254}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2241 ( .a ({signal_3690, signal_2232}), .b ({signal_3714, signal_2256}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2243 ( .a ({signal_3697, signal_2239}), .b ({signal_3716, signal_2258}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2249 ( .a ({signal_3620, signal_2162}), .b ({signal_6432, signal_6430}), .clk ( clk ), .r ( Fresh[762] ), .c ({signal_3722, signal_2264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2250 ( .a ({signal_3602, signal_2144}), .b ({signal_3661, signal_2203}), .clk ( clk ), .r ( Fresh[763] ), .c ({signal_3723, signal_2265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2251 ( .a ({signal_6436, signal_6434}), .b ({signal_3662, signal_2204}), .clk ( clk ), .r ( Fresh[764] ), .c ({signal_3724, signal_2266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2252 ( .a ({signal_6448, signal_6442}), .b ({signal_3664, signal_2206}), .clk ( clk ), .r ( Fresh[765] ), .c ({signal_3725, signal_2267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2253 ( .a ({signal_6452, signal_6450}), .b ({signal_3665, signal_2207}), .clk ( clk ), .r ( Fresh[766] ), .c ({signal_3726, signal_2268}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2254 ( .a ({signal_6456, signal_6454}), .b ({signal_3667, signal_2209}), .clk ( clk ), .r ( Fresh[767] ), .c ({signal_3727, signal_2269}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2271 ( .a ({signal_3724, signal_2266}), .b ({signal_3744, signal_2286}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2272 ( .a ({signal_3725, signal_2267}), .b ({signal_3745, signal_2287}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2273 ( .a ({signal_3726, signal_2268}), .b ({signal_3746, signal_2288}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2274 ( .a ({signal_3727, signal_2269}), .b ({signal_3747, signal_2289}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2282 ( .a ({signal_3708, signal_2250}), .b ({signal_6468, signal_6462}), .clk ( clk ), .r ( Fresh[768] ), .c ({signal_3755, signal_2297}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2283 ( .a ({signal_6452, signal_6450}), .b ({signal_3706, signal_2248}), .clk ( clk ), .r ( Fresh[769] ), .c ({signal_3756, signal_2298}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2285 ( .a ({signal_6480, signal_6474}), .b ({signal_3721, signal_2263}), .clk ( clk ), .r ( Fresh[770] ), .c ({signal_3758, signal_2300}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2286 ( .a ({signal_6488, signal_6484}), .b ({signal_3709, signal_2251}), .clk ( clk ), .r ( Fresh[771] ), .c ({signal_3759, signal_2301}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2297 ( .a ({signal_3756, signal_2298}), .b ({signal_3770, signal_2312}) ) ;
    buf_clk cell_4138 ( .C ( clk ), .D ( signal_6497 ), .Q ( signal_6498 ) ) ;
    buf_clk cell_4148 ( .C ( clk ), .D ( signal_6507 ), .Q ( signal_6508 ) ) ;
    buf_clk cell_4154 ( .C ( clk ), .D ( signal_6513 ), .Q ( signal_6514 ) ) ;
    buf_clk cell_4160 ( .C ( clk ), .D ( signal_6519 ), .Q ( signal_6520 ) ) ;
    buf_clk cell_4168 ( .C ( clk ), .D ( signal_6527 ), .Q ( signal_6528 ) ) ;
    buf_clk cell_4176 ( .C ( clk ), .D ( signal_6535 ), .Q ( signal_6536 ) ) ;
    buf_clk cell_4184 ( .C ( clk ), .D ( signal_6543 ), .Q ( signal_6544 ) ) ;
    buf_clk cell_4192 ( .C ( clk ), .D ( signal_6551 ), .Q ( signal_6552 ) ) ;
    buf_clk cell_4196 ( .C ( clk ), .D ( signal_6555 ), .Q ( signal_6556 ) ) ;
    buf_clk cell_4200 ( .C ( clk ), .D ( signal_6559 ), .Q ( signal_6560 ) ) ;
    buf_clk cell_4204 ( .C ( clk ), .D ( signal_6563 ), .Q ( signal_6564 ) ) ;
    buf_clk cell_4208 ( .C ( clk ), .D ( signal_6567 ), .Q ( signal_6568 ) ) ;
    buf_clk cell_4210 ( .C ( clk ), .D ( signal_6569 ), .Q ( signal_6570 ) ) ;
    buf_clk cell_4212 ( .C ( clk ), .D ( signal_6571 ), .Q ( signal_6572 ) ) ;
    buf_clk cell_4214 ( .C ( clk ), .D ( signal_6573 ), .Q ( signal_6574 ) ) ;
    buf_clk cell_4216 ( .C ( clk ), .D ( signal_6575 ), .Q ( signal_6576 ) ) ;
    buf_clk cell_4220 ( .C ( clk ), .D ( signal_6579 ), .Q ( signal_6580 ) ) ;
    buf_clk cell_4224 ( .C ( clk ), .D ( signal_6583 ), .Q ( signal_6584 ) ) ;
    buf_clk cell_4234 ( .C ( clk ), .D ( signal_6593 ), .Q ( signal_6594 ) ) ;
    buf_clk cell_4244 ( .C ( clk ), .D ( signal_6603 ), .Q ( signal_6604 ) ) ;
    buf_clk cell_4250 ( .C ( clk ), .D ( signal_6609 ), .Q ( signal_6610 ) ) ;
    buf_clk cell_4256 ( .C ( clk ), .D ( signal_6615 ), .Q ( signal_6616 ) ) ;
    buf_clk cell_4258 ( .C ( clk ), .D ( signal_6617 ), .Q ( signal_6618 ) ) ;
    buf_clk cell_4260 ( .C ( clk ), .D ( signal_6619 ), .Q ( signal_6620 ) ) ;
    buf_clk cell_4268 ( .C ( clk ), .D ( signal_6627 ), .Q ( signal_6628 ) ) ;
    buf_clk cell_4276 ( .C ( clk ), .D ( signal_6635 ), .Q ( signal_6636 ) ) ;
    buf_clk cell_4282 ( .C ( clk ), .D ( signal_6641 ), .Q ( signal_6642 ) ) ;
    buf_clk cell_4288 ( .C ( clk ), .D ( signal_6647 ), .Q ( signal_6648 ) ) ;
    buf_clk cell_4296 ( .C ( clk ), .D ( signal_6655 ), .Q ( signal_6656 ) ) ;
    buf_clk cell_4304 ( .C ( clk ), .D ( signal_6663 ), .Q ( signal_6664 ) ) ;
    buf_clk cell_4312 ( .C ( clk ), .D ( signal_6671 ), .Q ( signal_6672 ) ) ;
    buf_clk cell_4320 ( .C ( clk ), .D ( signal_6679 ), .Q ( signal_6680 ) ) ;
    buf_clk cell_4328 ( .C ( clk ), .D ( signal_6687 ), .Q ( signal_6688 ) ) ;
    buf_clk cell_4336 ( .C ( clk ), .D ( signal_6695 ), .Q ( signal_6696 ) ) ;
    buf_clk cell_4346 ( .C ( clk ), .D ( signal_6705 ), .Q ( signal_6706 ) ) ;
    buf_clk cell_4356 ( .C ( clk ), .D ( signal_6715 ), .Q ( signal_6716 ) ) ;
    buf_clk cell_4364 ( .C ( clk ), .D ( signal_6723 ), .Q ( signal_6724 ) ) ;
    buf_clk cell_4372 ( .C ( clk ), .D ( signal_6731 ), .Q ( signal_6732 ) ) ;
    buf_clk cell_4380 ( .C ( clk ), .D ( signal_6739 ), .Q ( signal_6740 ) ) ;
    buf_clk cell_4388 ( .C ( clk ), .D ( signal_6747 ), .Q ( signal_6748 ) ) ;
    buf_clk cell_4390 ( .C ( clk ), .D ( signal_6749 ), .Q ( signal_6750 ) ) ;
    buf_clk cell_4392 ( .C ( clk ), .D ( signal_6751 ), .Q ( signal_6752 ) ) ;
    buf_clk cell_4400 ( .C ( clk ), .D ( signal_6759 ), .Q ( signal_6760 ) ) ;
    buf_clk cell_4408 ( .C ( clk ), .D ( signal_6767 ), .Q ( signal_6768 ) ) ;
    buf_clk cell_4416 ( .C ( clk ), .D ( signal_6775 ), .Q ( signal_6776 ) ) ;
    buf_clk cell_4424 ( .C ( clk ), .D ( signal_6783 ), .Q ( signal_6784 ) ) ;
    buf_clk cell_4432 ( .C ( clk ), .D ( signal_6791 ), .Q ( signal_6792 ) ) ;
    buf_clk cell_4440 ( .C ( clk ), .D ( signal_6799 ), .Q ( signal_6800 ) ) ;
    buf_clk cell_4444 ( .C ( clk ), .D ( signal_6803 ), .Q ( signal_6804 ) ) ;
    buf_clk cell_4450 ( .C ( clk ), .D ( signal_6809 ), .Q ( signal_6810 ) ) ;
    buf_clk cell_4458 ( .C ( clk ), .D ( signal_6817 ), .Q ( signal_6818 ) ) ;
    buf_clk cell_4466 ( .C ( clk ), .D ( signal_6825 ), .Q ( signal_6826 ) ) ;
    buf_clk cell_4472 ( .C ( clk ), .D ( signal_6831 ), .Q ( signal_6832 ) ) ;
    buf_clk cell_4478 ( .C ( clk ), .D ( signal_6837 ), .Q ( signal_6838 ) ) ;
    buf_clk cell_4484 ( .C ( clk ), .D ( signal_6843 ), .Q ( signal_6844 ) ) ;
    buf_clk cell_4490 ( .C ( clk ), .D ( signal_6849 ), .Q ( signal_6850 ) ) ;
    buf_clk cell_4498 ( .C ( clk ), .D ( signal_6857 ), .Q ( signal_6858 ) ) ;
    buf_clk cell_4506 ( .C ( clk ), .D ( signal_6865 ), .Q ( signal_6866 ) ) ;
    buf_clk cell_4516 ( .C ( clk ), .D ( signal_6875 ), .Q ( signal_6876 ) ) ;
    buf_clk cell_4526 ( .C ( clk ), .D ( signal_6885 ), .Q ( signal_6886 ) ) ;
    buf_clk cell_4536 ( .C ( clk ), .D ( signal_6895 ), .Q ( signal_6896 ) ) ;
    buf_clk cell_4542 ( .C ( clk ), .D ( signal_6901 ), .Q ( signal_6902 ) ) ;
    buf_clk cell_4550 ( .C ( clk ), .D ( signal_6909 ), .Q ( signal_6910 ) ) ;
    buf_clk cell_4558 ( .C ( clk ), .D ( signal_6917 ), .Q ( signal_6918 ) ) ;
    buf_clk cell_4568 ( .C ( clk ), .D ( signal_6927 ), .Q ( signal_6928 ) ) ;
    buf_clk cell_4578 ( .C ( clk ), .D ( signal_6937 ), .Q ( signal_6938 ) ) ;
    buf_clk cell_4586 ( .C ( clk ), .D ( signal_6945 ), .Q ( signal_6946 ) ) ;
    buf_clk cell_4594 ( .C ( clk ), .D ( signal_6953 ), .Q ( signal_6954 ) ) ;
    buf_clk cell_4600 ( .C ( clk ), .D ( signal_6959 ), .Q ( signal_6960 ) ) ;
    buf_clk cell_4606 ( .C ( clk ), .D ( signal_6965 ), .Q ( signal_6966 ) ) ;
    buf_clk cell_4612 ( .C ( clk ), .D ( signal_6971 ), .Q ( signal_6972 ) ) ;
    buf_clk cell_4618 ( .C ( clk ), .D ( signal_6977 ), .Q ( signal_6978 ) ) ;
    buf_clk cell_4626 ( .C ( clk ), .D ( signal_6985 ), .Q ( signal_6986 ) ) ;
    buf_clk cell_4630 ( .C ( clk ), .D ( signal_6989 ), .Q ( signal_6990 ) ) ;
    buf_clk cell_4634 ( .C ( clk ), .D ( signal_6993 ), .Q ( signal_6994 ) ) ;
    buf_clk cell_4638 ( .C ( clk ), .D ( signal_6997 ), .Q ( signal_6998 ) ) ;
    buf_clk cell_4644 ( .C ( clk ), .D ( signal_7003 ), .Q ( signal_7004 ) ) ;
    buf_clk cell_4650 ( .C ( clk ), .D ( signal_7009 ), .Q ( signal_7010 ) ) ;
    buf_clk cell_4660 ( .C ( clk ), .D ( signal_7019 ), .Q ( signal_7020 ) ) ;
    buf_clk cell_4666 ( .C ( clk ), .D ( signal_7025 ), .Q ( signal_7026 ) ) ;
    buf_clk cell_4670 ( .C ( clk ), .D ( signal_7029 ), .Q ( signal_7030 ) ) ;
    buf_clk cell_4674 ( .C ( clk ), .D ( signal_7033 ), .Q ( signal_7034 ) ) ;
    buf_clk cell_4680 ( .C ( clk ), .D ( signal_7039 ), .Q ( signal_7040 ) ) ;
    buf_clk cell_4686 ( .C ( clk ), .D ( signal_7045 ), .Q ( signal_7046 ) ) ;
    buf_clk cell_4694 ( .C ( clk ), .D ( signal_7053 ), .Q ( signal_7054 ) ) ;
    buf_clk cell_4698 ( .C ( clk ), .D ( signal_7057 ), .Q ( signal_7058 ) ) ;
    buf_clk cell_4702 ( .C ( clk ), .D ( signal_7061 ), .Q ( signal_7062 ) ) ;
    buf_clk cell_4708 ( .C ( clk ), .D ( signal_7067 ), .Q ( signal_7068 ) ) ;
    buf_clk cell_4716 ( .C ( clk ), .D ( signal_7075 ), .Q ( signal_7076 ) ) ;
    buf_clk cell_4724 ( .C ( clk ), .D ( signal_7083 ), .Q ( signal_7084 ) ) ;
    buf_clk cell_4730 ( .C ( clk ), .D ( signal_7089 ), .Q ( signal_7090 ) ) ;
    buf_clk cell_4736 ( .C ( clk ), .D ( signal_7095 ), .Q ( signal_7096 ) ) ;
    buf_clk cell_4746 ( .C ( clk ), .D ( signal_7105 ), .Q ( signal_7106 ) ) ;
    buf_clk cell_4756 ( .C ( clk ), .D ( signal_7115 ), .Q ( signal_7116 ) ) ;
    buf_clk cell_4762 ( .C ( clk ), .D ( signal_7121 ), .Q ( signal_7122 ) ) ;
    buf_clk cell_4768 ( .C ( clk ), .D ( signal_7127 ), .Q ( signal_7128 ) ) ;
    buf_clk cell_4784 ( .C ( clk ), .D ( signal_7143 ), .Q ( signal_7144 ) ) ;
    buf_clk cell_4792 ( .C ( clk ), .D ( signal_7151 ), .Q ( signal_7152 ) ) ;
    buf_clk cell_4798 ( .C ( clk ), .D ( signal_7157 ), .Q ( signal_7158 ) ) ;
    buf_clk cell_4804 ( .C ( clk ), .D ( signal_7163 ), .Q ( signal_7164 ) ) ;
    buf_clk cell_4812 ( .C ( clk ), .D ( signal_7171 ), .Q ( signal_7172 ) ) ;
    buf_clk cell_4820 ( .C ( clk ), .D ( signal_7179 ), .Q ( signal_7180 ) ) ;
    buf_clk cell_4826 ( .C ( clk ), .D ( signal_7185 ), .Q ( signal_7186 ) ) ;
    buf_clk cell_4832 ( .C ( clk ), .D ( signal_7191 ), .Q ( signal_7192 ) ) ;
    buf_clk cell_4840 ( .C ( clk ), .D ( signal_7199 ), .Q ( signal_7200 ) ) ;
    buf_clk cell_4848 ( .C ( clk ), .D ( signal_7207 ), .Q ( signal_7208 ) ) ;
    buf_clk cell_4862 ( .C ( clk ), .D ( signal_7221 ), .Q ( signal_7222 ) ) ;
    buf_clk cell_4868 ( .C ( clk ), .D ( signal_7227 ), .Q ( signal_7228 ) ) ;
    buf_clk cell_4874 ( .C ( clk ), .D ( signal_7233 ), .Q ( signal_7234 ) ) ;
    buf_clk cell_4880 ( .C ( clk ), .D ( signal_7239 ), .Q ( signal_7240 ) ) ;
    buf_clk cell_4902 ( .C ( clk ), .D ( signal_7261 ), .Q ( signal_7262 ) ) ;
    buf_clk cell_4910 ( .C ( clk ), .D ( signal_7269 ), .Q ( signal_7270 ) ) ;
    buf_clk cell_4922 ( .C ( clk ), .D ( signal_7281 ), .Q ( signal_7282 ) ) ;
    buf_clk cell_4934 ( .C ( clk ), .D ( signal_7293 ), .Q ( signal_7294 ) ) ;
    buf_clk cell_4972 ( .C ( clk ), .D ( signal_7331 ), .Q ( signal_7332 ) ) ;
    buf_clk cell_4986 ( .C ( clk ), .D ( signal_7345 ), .Q ( signal_7346 ) ) ;
    buf_clk cell_4994 ( .C ( clk ), .D ( signal_7353 ), .Q ( signal_7354 ) ) ;
    buf_clk cell_5002 ( .C ( clk ), .D ( signal_7361 ), .Q ( signal_7362 ) ) ;
    buf_clk cell_5016 ( .C ( clk ), .D ( signal_7375 ), .Q ( signal_7376 ) ) ;
    buf_clk cell_5030 ( .C ( clk ), .D ( signal_7389 ), .Q ( signal_7390 ) ) ;
    buf_clk cell_5038 ( .C ( clk ), .D ( signal_7397 ), .Q ( signal_7398 ) ) ;
    buf_clk cell_5046 ( .C ( clk ), .D ( signal_7405 ), .Q ( signal_7406 ) ) ;
    buf_clk cell_5062 ( .C ( clk ), .D ( signal_7421 ), .Q ( signal_7422 ) ) ;
    buf_clk cell_5072 ( .C ( clk ), .D ( signal_7431 ), .Q ( signal_7432 ) ) ;
    buf_clk cell_5096 ( .C ( clk ), .D ( signal_7455 ), .Q ( signal_7456 ) ) ;
    buf_clk cell_5112 ( .C ( clk ), .D ( signal_7471 ), .Q ( signal_7472 ) ) ;
    buf_clk cell_5136 ( .C ( clk ), .D ( signal_7495 ), .Q ( signal_7496 ) ) ;
    buf_clk cell_5152 ( .C ( clk ), .D ( signal_7511 ), .Q ( signal_7512 ) ) ;
    buf_clk cell_5162 ( .C ( clk ), .D ( signal_7521 ), .Q ( signal_7522 ) ) ;
    buf_clk cell_5172 ( .C ( clk ), .D ( signal_7531 ), .Q ( signal_7532 ) ) ;
    buf_clk cell_5258 ( .C ( clk ), .D ( signal_7617 ), .Q ( signal_7618 ) ) ;
    buf_clk cell_5274 ( .C ( clk ), .D ( signal_7633 ), .Q ( signal_7634 ) ) ;
    buf_clk cell_5292 ( .C ( clk ), .D ( signal_7651 ), .Q ( signal_7652 ) ) ;
    buf_clk cell_5310 ( .C ( clk ), .D ( signal_7669 ), .Q ( signal_7670 ) ) ;
    buf_clk cell_5392 ( .C ( clk ), .D ( signal_7751 ), .Q ( signal_7752 ) ) ;
    buf_clk cell_5412 ( .C ( clk ), .D ( signal_7771 ), .Q ( signal_7772 ) ) ;

    /* cells in depth 15 */
    buf_clk cell_4445 ( .C ( clk ), .D ( signal_6804 ), .Q ( signal_6805 ) ) ;
    buf_clk cell_4451 ( .C ( clk ), .D ( signal_6810 ), .Q ( signal_6811 ) ) ;
    buf_clk cell_4459 ( .C ( clk ), .D ( signal_6818 ), .Q ( signal_6819 ) ) ;
    buf_clk cell_4467 ( .C ( clk ), .D ( signal_6826 ), .Q ( signal_6827 ) ) ;
    buf_clk cell_4473 ( .C ( clk ), .D ( signal_6832 ), .Q ( signal_6833 ) ) ;
    buf_clk cell_4479 ( .C ( clk ), .D ( signal_6838 ), .Q ( signal_6839 ) ) ;
    buf_clk cell_4485 ( .C ( clk ), .D ( signal_6844 ), .Q ( signal_6845 ) ) ;
    buf_clk cell_4491 ( .C ( clk ), .D ( signal_6850 ), .Q ( signal_6851 ) ) ;
    buf_clk cell_4499 ( .C ( clk ), .D ( signal_6858 ), .Q ( signal_6859 ) ) ;
    buf_clk cell_4507 ( .C ( clk ), .D ( signal_6866 ), .Q ( signal_6867 ) ) ;
    buf_clk cell_4517 ( .C ( clk ), .D ( signal_6876 ), .Q ( signal_6877 ) ) ;
    buf_clk cell_4527 ( .C ( clk ), .D ( signal_6886 ), .Q ( signal_6887 ) ) ;
    buf_clk cell_4529 ( .C ( clk ), .D ( signal_2258 ), .Q ( signal_6889 ) ) ;
    buf_clk cell_4531 ( .C ( clk ), .D ( signal_3716 ), .Q ( signal_6891 ) ) ;
    buf_clk cell_4537 ( .C ( clk ), .D ( signal_6896 ), .Q ( signal_6897 ) ) ;
    buf_clk cell_4543 ( .C ( clk ), .D ( signal_6902 ), .Q ( signal_6903 ) ) ;
    buf_clk cell_4551 ( .C ( clk ), .D ( signal_6910 ), .Q ( signal_6911 ) ) ;
    buf_clk cell_4559 ( .C ( clk ), .D ( signal_6918 ), .Q ( signal_6919 ) ) ;
    buf_clk cell_4569 ( .C ( clk ), .D ( signal_6928 ), .Q ( signal_6929 ) ) ;
    buf_clk cell_4579 ( .C ( clk ), .D ( signal_6938 ), .Q ( signal_6939 ) ) ;
    buf_clk cell_4587 ( .C ( clk ), .D ( signal_6946 ), .Q ( signal_6947 ) ) ;
    buf_clk cell_4595 ( .C ( clk ), .D ( signal_6954 ), .Q ( signal_6955 ) ) ;
    buf_clk cell_4601 ( .C ( clk ), .D ( signal_6960 ), .Q ( signal_6961 ) ) ;
    buf_clk cell_4607 ( .C ( clk ), .D ( signal_6966 ), .Q ( signal_6967 ) ) ;
    buf_clk cell_4613 ( .C ( clk ), .D ( signal_6972 ), .Q ( signal_6973 ) ) ;
    buf_clk cell_4619 ( .C ( clk ), .D ( signal_6978 ), .Q ( signal_6979 ) ) ;
    buf_clk cell_4621 ( .C ( clk ), .D ( signal_6570 ), .Q ( signal_6981 ) ) ;
    buf_clk cell_4623 ( .C ( clk ), .D ( signal_6572 ), .Q ( signal_6983 ) ) ;
    buf_clk cell_4627 ( .C ( clk ), .D ( signal_6986 ), .Q ( signal_6987 ) ) ;
    buf_clk cell_4631 ( .C ( clk ), .D ( signal_6990 ), .Q ( signal_6991 ) ) ;
    buf_clk cell_4635 ( .C ( clk ), .D ( signal_6994 ), .Q ( signal_6995 ) ) ;
    buf_clk cell_4639 ( .C ( clk ), .D ( signal_6998 ), .Q ( signal_6999 ) ) ;
    buf_clk cell_4645 ( .C ( clk ), .D ( signal_7004 ), .Q ( signal_7005 ) ) ;
    buf_clk cell_4651 ( .C ( clk ), .D ( signal_7010 ), .Q ( signal_7011 ) ) ;
    buf_clk cell_4653 ( .C ( clk ), .D ( signal_2287 ), .Q ( signal_7013 ) ) ;
    buf_clk cell_4655 ( .C ( clk ), .D ( signal_3745 ), .Q ( signal_7015 ) ) ;
    buf_clk cell_4661 ( .C ( clk ), .D ( signal_7020 ), .Q ( signal_7021 ) ) ;
    buf_clk cell_4667 ( .C ( clk ), .D ( signal_7026 ), .Q ( signal_7027 ) ) ;
    buf_clk cell_4671 ( .C ( clk ), .D ( signal_7030 ), .Q ( signal_7031 ) ) ;
    buf_clk cell_4675 ( .C ( clk ), .D ( signal_7034 ), .Q ( signal_7035 ) ) ;
    buf_clk cell_4681 ( .C ( clk ), .D ( signal_7040 ), .Q ( signal_7041 ) ) ;
    buf_clk cell_4687 ( .C ( clk ), .D ( signal_7046 ), .Q ( signal_7047 ) ) ;
    buf_clk cell_4689 ( .C ( clk ), .D ( signal_2312 ), .Q ( signal_7049 ) ) ;
    buf_clk cell_4691 ( .C ( clk ), .D ( signal_3770 ), .Q ( signal_7051 ) ) ;
    buf_clk cell_4695 ( .C ( clk ), .D ( signal_7054 ), .Q ( signal_7055 ) ) ;
    buf_clk cell_4699 ( .C ( clk ), .D ( signal_7058 ), .Q ( signal_7059 ) ) ;
    buf_clk cell_4703 ( .C ( clk ), .D ( signal_7062 ), .Q ( signal_7063 ) ) ;
    buf_clk cell_4709 ( .C ( clk ), .D ( signal_7068 ), .Q ( signal_7069 ) ) ;
    buf_clk cell_4717 ( .C ( clk ), .D ( signal_7076 ), .Q ( signal_7077 ) ) ;
    buf_clk cell_4725 ( .C ( clk ), .D ( signal_7084 ), .Q ( signal_7085 ) ) ;
    buf_clk cell_4731 ( .C ( clk ), .D ( signal_7090 ), .Q ( signal_7091 ) ) ;
    buf_clk cell_4737 ( .C ( clk ), .D ( signal_7096 ), .Q ( signal_7097 ) ) ;
    buf_clk cell_4747 ( .C ( clk ), .D ( signal_7106 ), .Q ( signal_7107 ) ) ;
    buf_clk cell_4757 ( .C ( clk ), .D ( signal_7116 ), .Q ( signal_7117 ) ) ;
    buf_clk cell_4763 ( .C ( clk ), .D ( signal_7122 ), .Q ( signal_7123 ) ) ;
    buf_clk cell_4769 ( .C ( clk ), .D ( signal_7128 ), .Q ( signal_7129 ) ) ;
    buf_clk cell_4773 ( .C ( clk ), .D ( signal_2288 ), .Q ( signal_7133 ) ) ;
    buf_clk cell_4777 ( .C ( clk ), .D ( signal_3746 ), .Q ( signal_7137 ) ) ;
    buf_clk cell_4785 ( .C ( clk ), .D ( signal_7144 ), .Q ( signal_7145 ) ) ;
    buf_clk cell_4793 ( .C ( clk ), .D ( signal_7152 ), .Q ( signal_7153 ) ) ;
    buf_clk cell_4799 ( .C ( clk ), .D ( signal_7158 ), .Q ( signal_7159 ) ) ;
    buf_clk cell_4805 ( .C ( clk ), .D ( signal_7164 ), .Q ( signal_7165 ) ) ;
    buf_clk cell_4813 ( .C ( clk ), .D ( signal_7172 ), .Q ( signal_7173 ) ) ;
    buf_clk cell_4821 ( .C ( clk ), .D ( signal_7180 ), .Q ( signal_7181 ) ) ;
    buf_clk cell_4827 ( .C ( clk ), .D ( signal_7186 ), .Q ( signal_7187 ) ) ;
    buf_clk cell_4833 ( .C ( clk ), .D ( signal_7192 ), .Q ( signal_7193 ) ) ;
    buf_clk cell_4841 ( .C ( clk ), .D ( signal_7200 ), .Q ( signal_7201 ) ) ;
    buf_clk cell_4849 ( .C ( clk ), .D ( signal_7208 ), .Q ( signal_7209 ) ) ;
    buf_clk cell_4853 ( .C ( clk ), .D ( signal_2213 ), .Q ( signal_7213 ) ) ;
    buf_clk cell_4857 ( .C ( clk ), .D ( signal_3671 ), .Q ( signal_7217 ) ) ;
    buf_clk cell_4863 ( .C ( clk ), .D ( signal_7222 ), .Q ( signal_7223 ) ) ;
    buf_clk cell_4869 ( .C ( clk ), .D ( signal_7228 ), .Q ( signal_7229 ) ) ;
    buf_clk cell_4875 ( .C ( clk ), .D ( signal_7234 ), .Q ( signal_7235 ) ) ;
    buf_clk cell_4881 ( .C ( clk ), .D ( signal_7240 ), .Q ( signal_7241 ) ) ;
    buf_clk cell_4885 ( .C ( clk ), .D ( signal_2189 ), .Q ( signal_7245 ) ) ;
    buf_clk cell_4889 ( .C ( clk ), .D ( signal_3647 ), .Q ( signal_7249 ) ) ;
    buf_clk cell_4893 ( .C ( clk ), .D ( signal_2138 ), .Q ( signal_7253 ) ) ;
    buf_clk cell_4897 ( .C ( clk ), .D ( signal_3596 ), .Q ( signal_7257 ) ) ;
    buf_clk cell_4903 ( .C ( clk ), .D ( signal_7262 ), .Q ( signal_7263 ) ) ;
    buf_clk cell_4911 ( .C ( clk ), .D ( signal_7270 ), .Q ( signal_7271 ) ) ;
    buf_clk cell_4923 ( .C ( clk ), .D ( signal_7282 ), .Q ( signal_7283 ) ) ;
    buf_clk cell_4935 ( .C ( clk ), .D ( signal_7294 ), .Q ( signal_7295 ) ) ;
    buf_clk cell_4941 ( .C ( clk ), .D ( signal_2238 ), .Q ( signal_7301 ) ) ;
    buf_clk cell_4947 ( .C ( clk ), .D ( signal_3696 ), .Q ( signal_7307 ) ) ;
    buf_clk cell_4953 ( .C ( clk ), .D ( signal_2210 ), .Q ( signal_7313 ) ) ;
    buf_clk cell_4959 ( .C ( clk ), .D ( signal_3668 ), .Q ( signal_7319 ) ) ;
    buf_clk cell_4973 ( .C ( clk ), .D ( signal_7332 ), .Q ( signal_7333 ) ) ;
    buf_clk cell_4987 ( .C ( clk ), .D ( signal_7346 ), .Q ( signal_7347 ) ) ;
    buf_clk cell_4995 ( .C ( clk ), .D ( signal_7354 ), .Q ( signal_7355 ) ) ;
    buf_clk cell_5003 ( .C ( clk ), .D ( signal_7362 ), .Q ( signal_7363 ) ) ;
    buf_clk cell_5017 ( .C ( clk ), .D ( signal_7376 ), .Q ( signal_7377 ) ) ;
    buf_clk cell_5031 ( .C ( clk ), .D ( signal_7390 ), .Q ( signal_7391 ) ) ;
    buf_clk cell_5039 ( .C ( clk ), .D ( signal_7398 ), .Q ( signal_7399 ) ) ;
    buf_clk cell_5047 ( .C ( clk ), .D ( signal_7406 ), .Q ( signal_7407 ) ) ;
    buf_clk cell_5063 ( .C ( clk ), .D ( signal_7422 ), .Q ( signal_7423 ) ) ;
    buf_clk cell_5073 ( .C ( clk ), .D ( signal_7432 ), .Q ( signal_7433 ) ) ;
    buf_clk cell_5097 ( .C ( clk ), .D ( signal_7456 ), .Q ( signal_7457 ) ) ;
    buf_clk cell_5113 ( .C ( clk ), .D ( signal_7472 ), .Q ( signal_7473 ) ) ;
    buf_clk cell_5137 ( .C ( clk ), .D ( signal_7496 ), .Q ( signal_7497 ) ) ;
    buf_clk cell_5153 ( .C ( clk ), .D ( signal_7512 ), .Q ( signal_7513 ) ) ;
    buf_clk cell_5163 ( .C ( clk ), .D ( signal_7522 ), .Q ( signal_7523 ) ) ;
    buf_clk cell_5173 ( .C ( clk ), .D ( signal_7532 ), .Q ( signal_7533 ) ) ;
    buf_clk cell_5201 ( .C ( clk ), .D ( signal_2289 ), .Q ( signal_7561 ) ) ;
    buf_clk cell_5211 ( .C ( clk ), .D ( signal_3747 ), .Q ( signal_7571 ) ) ;
    buf_clk cell_5233 ( .C ( clk ), .D ( signal_2265 ), .Q ( signal_7593 ) ) ;
    buf_clk cell_5243 ( .C ( clk ), .D ( signal_3723 ), .Q ( signal_7603 ) ) ;
    buf_clk cell_5259 ( .C ( clk ), .D ( signal_7618 ), .Q ( signal_7619 ) ) ;
    buf_clk cell_5275 ( .C ( clk ), .D ( signal_7634 ), .Q ( signal_7635 ) ) ;
    buf_clk cell_5293 ( .C ( clk ), .D ( signal_7652 ), .Q ( signal_7653 ) ) ;
    buf_clk cell_5311 ( .C ( clk ), .D ( signal_7670 ), .Q ( signal_7671 ) ) ;
    buf_clk cell_5393 ( .C ( clk ), .D ( signal_7752 ), .Q ( signal_7753 ) ) ;
    buf_clk cell_5413 ( .C ( clk ), .D ( signal_7772 ), .Q ( signal_7773 ) ) ;

    /* cells in depth 16 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2180 ( .a ({signal_6508, signal_6498}), .b ({signal_3589, signal_2131}), .clk ( clk ), .r ( Fresh[772] ), .c ({signal_3653, signal_2195}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2181 ( .a ({signal_6520, signal_6514}), .b ({signal_3591, signal_2133}), .clk ( clk ), .r ( Fresh[773] ), .c ({signal_3654, signal_2196}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2182 ( .a ({signal_6536, signal_6528}), .b ({signal_3594, signal_2136}), .clk ( clk ), .r ( Fresh[774] ), .c ({signal_3655, signal_2197}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2183 ( .a ({signal_6552, signal_6544}), .b ({signal_3595, signal_2137}), .clk ( clk ), .r ( Fresh[775] ), .c ({signal_3656, signal_2198}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2199 ( .a ({signal_3653, signal_2195}), .b ({signal_3672, signal_2214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2225 ( .a ({signal_6560, signal_6556}), .b ({signal_3643, signal_2185}), .clk ( clk ), .r ( Fresh[776] ), .c ({signal_3698, signal_2240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2226 ( .a ({signal_6568, signal_6564}), .b ({signal_3645, signal_2187}), .clk ( clk ), .r ( Fresh[777] ), .c ({signal_3699, signal_2241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2227 ( .a ({signal_6572, signal_6570}), .b ({signal_3613, signal_2155}), .clk ( clk ), .r ( Fresh[778] ), .c ({signal_3700, signal_2242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2228 ( .a ({signal_3650, signal_2192}), .b ({signal_6576, signal_6574}), .clk ( clk ), .r ( Fresh[779] ), .c ({signal_3701, signal_2243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2229 ( .a ({signal_6584, signal_6580}), .b ({signal_3652, signal_2194}), .clk ( clk ), .r ( Fresh[780] ), .c ({signal_3702, signal_2244}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2244 ( .a ({signal_3698, signal_2240}), .b ({signal_3717, signal_2259}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2245 ( .a ({signal_3700, signal_2242}), .b ({signal_3718, signal_2260}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2246 ( .a ({signal_3702, signal_2244}), .b ({signal_3719, signal_2261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2247 ( .a ({signal_6604, signal_6594}), .b ({signal_3673, signal_2215}), .clk ( clk ), .r ( Fresh[781] ), .c ({signal_3720, signal_2262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2255 ( .a ({signal_6616, signal_6610}), .b ({signal_3682, signal_2224}), .clk ( clk ), .r ( Fresh[782] ), .c ({signal_3728, signal_2270}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2256 ( .a ({signal_6620, signal_6618}), .b ({signal_3683, signal_2225}), .clk ( clk ), .r ( Fresh[783] ), .c ({signal_3729, signal_2271}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2257 ( .a ({signal_6636, signal_6628}), .b ({signal_3684, signal_2226}), .clk ( clk ), .r ( Fresh[784] ), .c ({signal_3730, signal_2272}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2258 ( .a ({signal_6648, signal_6642}), .b ({signal_3685, signal_2227}), .clk ( clk ), .r ( Fresh[785] ), .c ({signal_3731, signal_2273}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2259 ( .a ({signal_6664, signal_6656}), .b ({signal_3687, signal_2229}), .clk ( clk ), .r ( Fresh[786] ), .c ({signal_3732, signal_2274}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2260 ( .a ({signal_6680, signal_6672}), .b ({signal_3688, signal_2230}), .clk ( clk ), .r ( Fresh[787] ), .c ({signal_3733, signal_2275}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2261 ( .a ({signal_6696, signal_6688}), .b ({signal_3689, signal_2231}), .clk ( clk ), .r ( Fresh[788] ), .c ({signal_3734, signal_2276}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2262 ( .a ({signal_6560, signal_6556}), .b ({signal_3669, signal_2211}), .clk ( clk ), .r ( Fresh[789] ), .c ({signal_3735, signal_2277}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2263 ( .a ({signal_6716, signal_6706}), .b ({signal_3692, signal_2234}), .clk ( clk ), .r ( Fresh[790] ), .c ({signal_3736, signal_2278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2264 ( .a ({signal_3663, signal_2205}), .b ({signal_3693, signal_2235}), .clk ( clk ), .r ( Fresh[791] ), .c ({signal_3737, signal_2279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2265 ( .a ({signal_6732, signal_6724}), .b ({signal_3670, signal_2212}), .clk ( clk ), .r ( Fresh[792] ), .c ({signal_3738, signal_2280}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2266 ( .a ({signal_6748, signal_6740}), .b ({signal_3695, signal_2237}), .clk ( clk ), .r ( Fresh[793] ), .c ({signal_3739, signal_2281}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2275 ( .a ({signal_3729, signal_2271}), .b ({signal_3748, signal_2290}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2276 ( .a ({signal_3730, signal_2272}), .b ({signal_3749, signal_2291}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2277 ( .a ({signal_3732, signal_2274}), .b ({signal_3750, signal_2292}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2278 ( .a ({signal_3734, signal_2276}), .b ({signal_3751, signal_2293}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2279 ( .a ({signal_3735, signal_2277}), .b ({signal_3752, signal_2294}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2280 ( .a ({signal_3738, signal_2280}), .b ({signal_3753, signal_2295}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2287 ( .a ({signal_3722, signal_2264}), .b ({signal_3680, signal_2222}), .clk ( clk ), .r ( Fresh[794] ), .c ({signal_3760, signal_2302}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2288 ( .a ({signal_6752, signal_6750}), .b ({signal_3712, signal_2254}), .clk ( clk ), .r ( Fresh[795] ), .c ({signal_3761, signal_2303}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2290 ( .a ({signal_6752, signal_6750}), .b ({signal_3714, signal_2256}), .clk ( clk ), .r ( Fresh[796] ), .c ({signal_3763, signal_2305}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2299 ( .a ({signal_3761, signal_2303}), .b ({signal_3772, signal_2314}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2301 ( .a ({signal_3763, signal_2305}), .b ({signal_3774, signal_2316}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2304 ( .a ({signal_6768, signal_6760}), .b ({signal_3755, signal_2297}), .clk ( clk ), .r ( Fresh[797] ), .c ({signal_3777, signal_2319}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2305 ( .a ({signal_6784, signal_6776}), .b ({signal_3758, signal_2300}), .clk ( clk ), .r ( Fresh[798] ), .c ({signal_3778, signal_2320}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2306 ( .a ({signal_6800, signal_6792}), .b ({signal_3759, signal_2301}), .clk ( clk ), .r ( Fresh[799] ), .c ({signal_3779, signal_2321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2307 ( .a ({signal_3744, signal_2286}), .b ({signal_3691, signal_2233}), .clk ( clk ), .r ( Fresh[800] ), .c ({signal_3780, signal_2322}) ) ;
    buf_clk cell_4446 ( .C ( clk ), .D ( signal_6805 ), .Q ( signal_6806 ) ) ;
    buf_clk cell_4452 ( .C ( clk ), .D ( signal_6811 ), .Q ( signal_6812 ) ) ;
    buf_clk cell_4460 ( .C ( clk ), .D ( signal_6819 ), .Q ( signal_6820 ) ) ;
    buf_clk cell_4468 ( .C ( clk ), .D ( signal_6827 ), .Q ( signal_6828 ) ) ;
    buf_clk cell_4474 ( .C ( clk ), .D ( signal_6833 ), .Q ( signal_6834 ) ) ;
    buf_clk cell_4480 ( .C ( clk ), .D ( signal_6839 ), .Q ( signal_6840 ) ) ;
    buf_clk cell_4486 ( .C ( clk ), .D ( signal_6845 ), .Q ( signal_6846 ) ) ;
    buf_clk cell_4492 ( .C ( clk ), .D ( signal_6851 ), .Q ( signal_6852 ) ) ;
    buf_clk cell_4500 ( .C ( clk ), .D ( signal_6859 ), .Q ( signal_6860 ) ) ;
    buf_clk cell_4508 ( .C ( clk ), .D ( signal_6867 ), .Q ( signal_6868 ) ) ;
    buf_clk cell_4518 ( .C ( clk ), .D ( signal_6877 ), .Q ( signal_6878 ) ) ;
    buf_clk cell_4528 ( .C ( clk ), .D ( signal_6887 ), .Q ( signal_6888 ) ) ;
    buf_clk cell_4530 ( .C ( clk ), .D ( signal_6889 ), .Q ( signal_6890 ) ) ;
    buf_clk cell_4532 ( .C ( clk ), .D ( signal_6891 ), .Q ( signal_6892 ) ) ;
    buf_clk cell_4538 ( .C ( clk ), .D ( signal_6897 ), .Q ( signal_6898 ) ) ;
    buf_clk cell_4544 ( .C ( clk ), .D ( signal_6903 ), .Q ( signal_6904 ) ) ;
    buf_clk cell_4552 ( .C ( clk ), .D ( signal_6911 ), .Q ( signal_6912 ) ) ;
    buf_clk cell_4560 ( .C ( clk ), .D ( signal_6919 ), .Q ( signal_6920 ) ) ;
    buf_clk cell_4570 ( .C ( clk ), .D ( signal_6929 ), .Q ( signal_6930 ) ) ;
    buf_clk cell_4580 ( .C ( clk ), .D ( signal_6939 ), .Q ( signal_6940 ) ) ;
    buf_clk cell_4588 ( .C ( clk ), .D ( signal_6947 ), .Q ( signal_6948 ) ) ;
    buf_clk cell_4596 ( .C ( clk ), .D ( signal_6955 ), .Q ( signal_6956 ) ) ;
    buf_clk cell_4602 ( .C ( clk ), .D ( signal_6961 ), .Q ( signal_6962 ) ) ;
    buf_clk cell_4608 ( .C ( clk ), .D ( signal_6967 ), .Q ( signal_6968 ) ) ;
    buf_clk cell_4614 ( .C ( clk ), .D ( signal_6973 ), .Q ( signal_6974 ) ) ;
    buf_clk cell_4620 ( .C ( clk ), .D ( signal_6979 ), .Q ( signal_6980 ) ) ;
    buf_clk cell_4622 ( .C ( clk ), .D ( signal_6981 ), .Q ( signal_6982 ) ) ;
    buf_clk cell_4624 ( .C ( clk ), .D ( signal_6983 ), .Q ( signal_6984 ) ) ;
    buf_clk cell_4628 ( .C ( clk ), .D ( signal_6987 ), .Q ( signal_6988 ) ) ;
    buf_clk cell_4632 ( .C ( clk ), .D ( signal_6991 ), .Q ( signal_6992 ) ) ;
    buf_clk cell_4636 ( .C ( clk ), .D ( signal_6995 ), .Q ( signal_6996 ) ) ;
    buf_clk cell_4640 ( .C ( clk ), .D ( signal_6999 ), .Q ( signal_7000 ) ) ;
    buf_clk cell_4646 ( .C ( clk ), .D ( signal_7005 ), .Q ( signal_7006 ) ) ;
    buf_clk cell_4652 ( .C ( clk ), .D ( signal_7011 ), .Q ( signal_7012 ) ) ;
    buf_clk cell_4654 ( .C ( clk ), .D ( signal_7013 ), .Q ( signal_7014 ) ) ;
    buf_clk cell_4656 ( .C ( clk ), .D ( signal_7015 ), .Q ( signal_7016 ) ) ;
    buf_clk cell_4662 ( .C ( clk ), .D ( signal_7021 ), .Q ( signal_7022 ) ) ;
    buf_clk cell_4668 ( .C ( clk ), .D ( signal_7027 ), .Q ( signal_7028 ) ) ;
    buf_clk cell_4672 ( .C ( clk ), .D ( signal_7031 ), .Q ( signal_7032 ) ) ;
    buf_clk cell_4676 ( .C ( clk ), .D ( signal_7035 ), .Q ( signal_7036 ) ) ;
    buf_clk cell_4682 ( .C ( clk ), .D ( signal_7041 ), .Q ( signal_7042 ) ) ;
    buf_clk cell_4688 ( .C ( clk ), .D ( signal_7047 ), .Q ( signal_7048 ) ) ;
    buf_clk cell_4690 ( .C ( clk ), .D ( signal_7049 ), .Q ( signal_7050 ) ) ;
    buf_clk cell_4692 ( .C ( clk ), .D ( signal_7051 ), .Q ( signal_7052 ) ) ;
    buf_clk cell_4696 ( .C ( clk ), .D ( signal_7055 ), .Q ( signal_7056 ) ) ;
    buf_clk cell_4700 ( .C ( clk ), .D ( signal_7059 ), .Q ( signal_7060 ) ) ;
    buf_clk cell_4704 ( .C ( clk ), .D ( signal_7063 ), .Q ( signal_7064 ) ) ;
    buf_clk cell_4710 ( .C ( clk ), .D ( signal_7069 ), .Q ( signal_7070 ) ) ;
    buf_clk cell_4718 ( .C ( clk ), .D ( signal_7077 ), .Q ( signal_7078 ) ) ;
    buf_clk cell_4726 ( .C ( clk ), .D ( signal_7085 ), .Q ( signal_7086 ) ) ;
    buf_clk cell_4732 ( .C ( clk ), .D ( signal_7091 ), .Q ( signal_7092 ) ) ;
    buf_clk cell_4738 ( .C ( clk ), .D ( signal_7097 ), .Q ( signal_7098 ) ) ;
    buf_clk cell_4748 ( .C ( clk ), .D ( signal_7107 ), .Q ( signal_7108 ) ) ;
    buf_clk cell_4758 ( .C ( clk ), .D ( signal_7117 ), .Q ( signal_7118 ) ) ;
    buf_clk cell_4764 ( .C ( clk ), .D ( signal_7123 ), .Q ( signal_7124 ) ) ;
    buf_clk cell_4770 ( .C ( clk ), .D ( signal_7129 ), .Q ( signal_7130 ) ) ;
    buf_clk cell_4774 ( .C ( clk ), .D ( signal_7133 ), .Q ( signal_7134 ) ) ;
    buf_clk cell_4778 ( .C ( clk ), .D ( signal_7137 ), .Q ( signal_7138 ) ) ;
    buf_clk cell_4786 ( .C ( clk ), .D ( signal_7145 ), .Q ( signal_7146 ) ) ;
    buf_clk cell_4794 ( .C ( clk ), .D ( signal_7153 ), .Q ( signal_7154 ) ) ;
    buf_clk cell_4800 ( .C ( clk ), .D ( signal_7159 ), .Q ( signal_7160 ) ) ;
    buf_clk cell_4806 ( .C ( clk ), .D ( signal_7165 ), .Q ( signal_7166 ) ) ;
    buf_clk cell_4814 ( .C ( clk ), .D ( signal_7173 ), .Q ( signal_7174 ) ) ;
    buf_clk cell_4822 ( .C ( clk ), .D ( signal_7181 ), .Q ( signal_7182 ) ) ;
    buf_clk cell_4828 ( .C ( clk ), .D ( signal_7187 ), .Q ( signal_7188 ) ) ;
    buf_clk cell_4834 ( .C ( clk ), .D ( signal_7193 ), .Q ( signal_7194 ) ) ;
    buf_clk cell_4842 ( .C ( clk ), .D ( signal_7201 ), .Q ( signal_7202 ) ) ;
    buf_clk cell_4850 ( .C ( clk ), .D ( signal_7209 ), .Q ( signal_7210 ) ) ;
    buf_clk cell_4854 ( .C ( clk ), .D ( signal_7213 ), .Q ( signal_7214 ) ) ;
    buf_clk cell_4858 ( .C ( clk ), .D ( signal_7217 ), .Q ( signal_7218 ) ) ;
    buf_clk cell_4864 ( .C ( clk ), .D ( signal_7223 ), .Q ( signal_7224 ) ) ;
    buf_clk cell_4870 ( .C ( clk ), .D ( signal_7229 ), .Q ( signal_7230 ) ) ;
    buf_clk cell_4876 ( .C ( clk ), .D ( signal_7235 ), .Q ( signal_7236 ) ) ;
    buf_clk cell_4882 ( .C ( clk ), .D ( signal_7241 ), .Q ( signal_7242 ) ) ;
    buf_clk cell_4886 ( .C ( clk ), .D ( signal_7245 ), .Q ( signal_7246 ) ) ;
    buf_clk cell_4890 ( .C ( clk ), .D ( signal_7249 ), .Q ( signal_7250 ) ) ;
    buf_clk cell_4894 ( .C ( clk ), .D ( signal_7253 ), .Q ( signal_7254 ) ) ;
    buf_clk cell_4898 ( .C ( clk ), .D ( signal_7257 ), .Q ( signal_7258 ) ) ;
    buf_clk cell_4904 ( .C ( clk ), .D ( signal_7263 ), .Q ( signal_7264 ) ) ;
    buf_clk cell_4912 ( .C ( clk ), .D ( signal_7271 ), .Q ( signal_7272 ) ) ;
    buf_clk cell_4924 ( .C ( clk ), .D ( signal_7283 ), .Q ( signal_7284 ) ) ;
    buf_clk cell_4936 ( .C ( clk ), .D ( signal_7295 ), .Q ( signal_7296 ) ) ;
    buf_clk cell_4942 ( .C ( clk ), .D ( signal_7301 ), .Q ( signal_7302 ) ) ;
    buf_clk cell_4948 ( .C ( clk ), .D ( signal_7307 ), .Q ( signal_7308 ) ) ;
    buf_clk cell_4954 ( .C ( clk ), .D ( signal_7313 ), .Q ( signal_7314 ) ) ;
    buf_clk cell_4960 ( .C ( clk ), .D ( signal_7319 ), .Q ( signal_7320 ) ) ;
    buf_clk cell_4974 ( .C ( clk ), .D ( signal_7333 ), .Q ( signal_7334 ) ) ;
    buf_clk cell_4988 ( .C ( clk ), .D ( signal_7347 ), .Q ( signal_7348 ) ) ;
    buf_clk cell_4996 ( .C ( clk ), .D ( signal_7355 ), .Q ( signal_7356 ) ) ;
    buf_clk cell_5004 ( .C ( clk ), .D ( signal_7363 ), .Q ( signal_7364 ) ) ;
    buf_clk cell_5018 ( .C ( clk ), .D ( signal_7377 ), .Q ( signal_7378 ) ) ;
    buf_clk cell_5032 ( .C ( clk ), .D ( signal_7391 ), .Q ( signal_7392 ) ) ;
    buf_clk cell_5040 ( .C ( clk ), .D ( signal_7399 ), .Q ( signal_7400 ) ) ;
    buf_clk cell_5048 ( .C ( clk ), .D ( signal_7407 ), .Q ( signal_7408 ) ) ;
    buf_clk cell_5064 ( .C ( clk ), .D ( signal_7423 ), .Q ( signal_7424 ) ) ;
    buf_clk cell_5074 ( .C ( clk ), .D ( signal_7433 ), .Q ( signal_7434 ) ) ;
    buf_clk cell_5098 ( .C ( clk ), .D ( signal_7457 ), .Q ( signal_7458 ) ) ;
    buf_clk cell_5114 ( .C ( clk ), .D ( signal_7473 ), .Q ( signal_7474 ) ) ;
    buf_clk cell_5138 ( .C ( clk ), .D ( signal_7497 ), .Q ( signal_7498 ) ) ;
    buf_clk cell_5154 ( .C ( clk ), .D ( signal_7513 ), .Q ( signal_7514 ) ) ;
    buf_clk cell_5164 ( .C ( clk ), .D ( signal_7523 ), .Q ( signal_7524 ) ) ;
    buf_clk cell_5174 ( .C ( clk ), .D ( signal_7533 ), .Q ( signal_7534 ) ) ;
    buf_clk cell_5202 ( .C ( clk ), .D ( signal_7561 ), .Q ( signal_7562 ) ) ;
    buf_clk cell_5212 ( .C ( clk ), .D ( signal_7571 ), .Q ( signal_7572 ) ) ;
    buf_clk cell_5234 ( .C ( clk ), .D ( signal_7593 ), .Q ( signal_7594 ) ) ;
    buf_clk cell_5244 ( .C ( clk ), .D ( signal_7603 ), .Q ( signal_7604 ) ) ;
    buf_clk cell_5260 ( .C ( clk ), .D ( signal_7619 ), .Q ( signal_7620 ) ) ;
    buf_clk cell_5276 ( .C ( clk ), .D ( signal_7635 ), .Q ( signal_7636 ) ) ;
    buf_clk cell_5294 ( .C ( clk ), .D ( signal_7653 ), .Q ( signal_7654 ) ) ;
    buf_clk cell_5312 ( .C ( clk ), .D ( signal_7671 ), .Q ( signal_7672 ) ) ;
    buf_clk cell_5394 ( .C ( clk ), .D ( signal_7753 ), .Q ( signal_7754 ) ) ;
    buf_clk cell_5414 ( .C ( clk ), .D ( signal_7773 ), .Q ( signal_7774 ) ) ;

    /* cells in depth 17 */
    buf_clk cell_4705 ( .C ( clk ), .D ( signal_7064 ), .Q ( signal_7065 ) ) ;
    buf_clk cell_4711 ( .C ( clk ), .D ( signal_7070 ), .Q ( signal_7071 ) ) ;
    buf_clk cell_4719 ( .C ( clk ), .D ( signal_7078 ), .Q ( signal_7079 ) ) ;
    buf_clk cell_4727 ( .C ( clk ), .D ( signal_7086 ), .Q ( signal_7087 ) ) ;
    buf_clk cell_4733 ( .C ( clk ), .D ( signal_7092 ), .Q ( signal_7093 ) ) ;
    buf_clk cell_4739 ( .C ( clk ), .D ( signal_7098 ), .Q ( signal_7099 ) ) ;
    buf_clk cell_4749 ( .C ( clk ), .D ( signal_7108 ), .Q ( signal_7109 ) ) ;
    buf_clk cell_4759 ( .C ( clk ), .D ( signal_7118 ), .Q ( signal_7119 ) ) ;
    buf_clk cell_4765 ( .C ( clk ), .D ( signal_7124 ), .Q ( signal_7125 ) ) ;
    buf_clk cell_4771 ( .C ( clk ), .D ( signal_7130 ), .Q ( signal_7131 ) ) ;
    buf_clk cell_4775 ( .C ( clk ), .D ( signal_7134 ), .Q ( signal_7135 ) ) ;
    buf_clk cell_4779 ( .C ( clk ), .D ( signal_7138 ), .Q ( signal_7139 ) ) ;
    buf_clk cell_4787 ( .C ( clk ), .D ( signal_7146 ), .Q ( signal_7147 ) ) ;
    buf_clk cell_4795 ( .C ( clk ), .D ( signal_7154 ), .Q ( signal_7155 ) ) ;
    buf_clk cell_4801 ( .C ( clk ), .D ( signal_7160 ), .Q ( signal_7161 ) ) ;
    buf_clk cell_4807 ( .C ( clk ), .D ( signal_7166 ), .Q ( signal_7167 ) ) ;
    buf_clk cell_4815 ( .C ( clk ), .D ( signal_7174 ), .Q ( signal_7175 ) ) ;
    buf_clk cell_4823 ( .C ( clk ), .D ( signal_7182 ), .Q ( signal_7183 ) ) ;
    buf_clk cell_4829 ( .C ( clk ), .D ( signal_7188 ), .Q ( signal_7189 ) ) ;
    buf_clk cell_4835 ( .C ( clk ), .D ( signal_7194 ), .Q ( signal_7195 ) ) ;
    buf_clk cell_4843 ( .C ( clk ), .D ( signal_7202 ), .Q ( signal_7203 ) ) ;
    buf_clk cell_4851 ( .C ( clk ), .D ( signal_7210 ), .Q ( signal_7211 ) ) ;
    buf_clk cell_4855 ( .C ( clk ), .D ( signal_7214 ), .Q ( signal_7215 ) ) ;
    buf_clk cell_4859 ( .C ( clk ), .D ( signal_7218 ), .Q ( signal_7219 ) ) ;
    buf_clk cell_4865 ( .C ( clk ), .D ( signal_7224 ), .Q ( signal_7225 ) ) ;
    buf_clk cell_4871 ( .C ( clk ), .D ( signal_7230 ), .Q ( signal_7231 ) ) ;
    buf_clk cell_4877 ( .C ( clk ), .D ( signal_7236 ), .Q ( signal_7237 ) ) ;
    buf_clk cell_4883 ( .C ( clk ), .D ( signal_7242 ), .Q ( signal_7243 ) ) ;
    buf_clk cell_4887 ( .C ( clk ), .D ( signal_7246 ), .Q ( signal_7247 ) ) ;
    buf_clk cell_4891 ( .C ( clk ), .D ( signal_7250 ), .Q ( signal_7251 ) ) ;
    buf_clk cell_4895 ( .C ( clk ), .D ( signal_7254 ), .Q ( signal_7255 ) ) ;
    buf_clk cell_4899 ( .C ( clk ), .D ( signal_7258 ), .Q ( signal_7259 ) ) ;
    buf_clk cell_4905 ( .C ( clk ), .D ( signal_7264 ), .Q ( signal_7265 ) ) ;
    buf_clk cell_4913 ( .C ( clk ), .D ( signal_7272 ), .Q ( signal_7273 ) ) ;
    buf_clk cell_4925 ( .C ( clk ), .D ( signal_7284 ), .Q ( signal_7285 ) ) ;
    buf_clk cell_4937 ( .C ( clk ), .D ( signal_7296 ), .Q ( signal_7297 ) ) ;
    buf_clk cell_4943 ( .C ( clk ), .D ( signal_7302 ), .Q ( signal_7303 ) ) ;
    buf_clk cell_4949 ( .C ( clk ), .D ( signal_7308 ), .Q ( signal_7309 ) ) ;
    buf_clk cell_4955 ( .C ( clk ), .D ( signal_7314 ), .Q ( signal_7315 ) ) ;
    buf_clk cell_4961 ( .C ( clk ), .D ( signal_7320 ), .Q ( signal_7321 ) ) ;
    buf_clk cell_4975 ( .C ( clk ), .D ( signal_7334 ), .Q ( signal_7335 ) ) ;
    buf_clk cell_4989 ( .C ( clk ), .D ( signal_7348 ), .Q ( signal_7349 ) ) ;
    buf_clk cell_4997 ( .C ( clk ), .D ( signal_7356 ), .Q ( signal_7357 ) ) ;
    buf_clk cell_5005 ( .C ( clk ), .D ( signal_7364 ), .Q ( signal_7365 ) ) ;
    buf_clk cell_5019 ( .C ( clk ), .D ( signal_7378 ), .Q ( signal_7379 ) ) ;
    buf_clk cell_5033 ( .C ( clk ), .D ( signal_7392 ), .Q ( signal_7393 ) ) ;
    buf_clk cell_5041 ( .C ( clk ), .D ( signal_7400 ), .Q ( signal_7401 ) ) ;
    buf_clk cell_5049 ( .C ( clk ), .D ( signal_7408 ), .Q ( signal_7409 ) ) ;
    buf_clk cell_5065 ( .C ( clk ), .D ( signal_7424 ), .Q ( signal_7425 ) ) ;
    buf_clk cell_5075 ( .C ( clk ), .D ( signal_7434 ), .Q ( signal_7435 ) ) ;
    buf_clk cell_5099 ( .C ( clk ), .D ( signal_7458 ), .Q ( signal_7459 ) ) ;
    buf_clk cell_5115 ( .C ( clk ), .D ( signal_7474 ), .Q ( signal_7475 ) ) ;
    buf_clk cell_5139 ( .C ( clk ), .D ( signal_7498 ), .Q ( signal_7499 ) ) ;
    buf_clk cell_5155 ( .C ( clk ), .D ( signal_7514 ), .Q ( signal_7515 ) ) ;
    buf_clk cell_5165 ( .C ( clk ), .D ( signal_7524 ), .Q ( signal_7525 ) ) ;
    buf_clk cell_5175 ( .C ( clk ), .D ( signal_7534 ), .Q ( signal_7535 ) ) ;
    buf_clk cell_5203 ( .C ( clk ), .D ( signal_7562 ), .Q ( signal_7563 ) ) ;
    buf_clk cell_5213 ( .C ( clk ), .D ( signal_7572 ), .Q ( signal_7573 ) ) ;
    buf_clk cell_5235 ( .C ( clk ), .D ( signal_7594 ), .Q ( signal_7595 ) ) ;
    buf_clk cell_5245 ( .C ( clk ), .D ( signal_7604 ), .Q ( signal_7605 ) ) ;
    buf_clk cell_5261 ( .C ( clk ), .D ( signal_7620 ), .Q ( signal_7621 ) ) ;
    buf_clk cell_5277 ( .C ( clk ), .D ( signal_7636 ), .Q ( signal_7637 ) ) ;
    buf_clk cell_5295 ( .C ( clk ), .D ( signal_7654 ), .Q ( signal_7655 ) ) ;
    buf_clk cell_5313 ( .C ( clk ), .D ( signal_7672 ), .Q ( signal_7673 ) ) ;
    buf_clk cell_5329 ( .C ( clk ), .D ( signal_2281 ), .Q ( signal_7689 ) ) ;
    buf_clk cell_5337 ( .C ( clk ), .D ( signal_3739 ), .Q ( signal_7697 ) ) ;
    buf_clk cell_5395 ( .C ( clk ), .D ( signal_7754 ), .Q ( signal_7755 ) ) ;
    buf_clk cell_5415 ( .C ( clk ), .D ( signal_7774 ), .Q ( signal_7775 ) ) ;
    buf_clk cell_5441 ( .C ( clk ), .D ( signal_2260 ), .Q ( signal_7801 ) ) ;
    buf_clk cell_5453 ( .C ( clk ), .D ( signal_3718 ), .Q ( signal_7813 ) ) ;
    buf_clk cell_5465 ( .C ( clk ), .D ( signal_2322 ), .Q ( signal_7825 ) ) ;
    buf_clk cell_5479 ( .C ( clk ), .D ( signal_3780 ), .Q ( signal_7839 ) ) ;

    /* cells in depth 18 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2230 ( .a ({signal_6812, signal_6806}), .b ({signal_3654, signal_2196}), .clk ( clk ), .r ( Fresh[801] ), .c ({signal_3703, signal_2245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2231 ( .a ({signal_6828, signal_6820}), .b ({signal_3655, signal_2197}), .clk ( clk ), .r ( Fresh[802] ), .c ({signal_3704, signal_2246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2232 ( .a ({signal_6840, signal_6834}), .b ({signal_3656, signal_2198}), .clk ( clk ), .r ( Fresh[803] ), .c ({signal_3705, signal_2247}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2267 ( .a ({signal_6852, signal_6846}), .b ({signal_3699, signal_2241}), .clk ( clk ), .r ( Fresh[804] ), .c ({signal_3740, signal_2282}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2268 ( .a ({signal_6868, signal_6860}), .b ({signal_3672, signal_2214}), .clk ( clk ), .r ( Fresh[805] ), .c ({signal_3741, signal_2283}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2281 ( .a ({signal_3741, signal_2283}), .b ({signal_3754, signal_2296}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2284 ( .a ({signal_6888, signal_6878}), .b ({signal_3720, signal_2262}), .clk ( clk ), .r ( Fresh[806] ), .c ({signal_3757, signal_2299}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2289 ( .a ({signal_6892, signal_6890}), .b ({signal_3717, signal_2259}), .clk ( clk ), .r ( Fresh[807] ), .c ({signal_3762, signal_2304}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2291 ( .a ({signal_6904, signal_6898}), .b ({signal_3728, signal_2270}), .clk ( clk ), .r ( Fresh[808] ), .c ({signal_3764, signal_2306}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2292 ( .a ({signal_6920, signal_6912}), .b ({signal_3731, signal_2273}), .clk ( clk ), .r ( Fresh[809] ), .c ({signal_3765, signal_2307}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2293 ( .a ({signal_6940, signal_6930}), .b ({signal_3733, signal_2275}), .clk ( clk ), .r ( Fresh[810] ), .c ({signal_3766, signal_2308}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2294 ( .a ({signal_6956, signal_6948}), .b ({signal_3736, signal_2278}), .clk ( clk ), .r ( Fresh[811] ), .c ({signal_3767, signal_2309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2295 ( .a ({signal_6968, signal_6962}), .b ({signal_3719, signal_2261}), .clk ( clk ), .r ( Fresh[812] ), .c ({signal_3768, signal_2310}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2298 ( .a ({signal_3757, signal_2299}), .b ({signal_3771, signal_2313}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2300 ( .a ({signal_3762, signal_2304}), .b ({signal_3773, signal_2315}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2302 ( .a ({signal_3767, signal_2309}), .b ({signal_3775, signal_2317}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2303 ( .a ({signal_3768, signal_2310}), .b ({signal_3776, signal_2318}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2308 ( .a ({signal_6980, signal_6974}), .b ({signal_3748, signal_2290}), .clk ( clk ), .r ( Fresh[813] ), .c ({signal_3781, signal_2323}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2309 ( .a ({signal_6984, signal_6982}), .b ({signal_3749, signal_2291}), .clk ( clk ), .r ( Fresh[814] ), .c ({signal_3782, signal_2324}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2310 ( .a ({signal_6984, signal_6982}), .b ({signal_3750, signal_2292}), .clk ( clk ), .r ( Fresh[815] ), .c ({signal_3783, signal_2325}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2311 ( .a ({signal_6992, signal_6988}), .b ({signal_3751, signal_2293}), .clk ( clk ), .r ( Fresh[816] ), .c ({signal_3784, signal_2326}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2312 ( .a ({signal_7000, signal_6996}), .b ({signal_3752, signal_2294}), .clk ( clk ), .r ( Fresh[817] ), .c ({signal_3785, signal_2327}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2313 ( .a ({signal_3760, signal_2302}), .b ({signal_3737, signal_2279}), .clk ( clk ), .r ( Fresh[818] ), .c ({signal_3786, signal_2328}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2314 ( .a ({signal_7012, signal_7006}), .b ({signal_3753, signal_2295}), .clk ( clk ), .r ( Fresh[819] ), .c ({signal_3787, signal_2329}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2315 ( .a ({signal_7016, signal_7014}), .b ({signal_3701, signal_2243}), .clk ( clk ), .r ( Fresh[820] ), .c ({signal_3788, signal_2330}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2320 ( .a ({signal_3781, signal_2323}), .b ({signal_3793, signal_2335}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2321 ( .a ({signal_3782, signal_2324}), .b ({signal_3794, signal_2336}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2322 ( .a ({signal_3783, signal_2325}), .b ({signal_3795, signal_2337}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2323 ( .a ({signal_3784, signal_2326}), .b ({signal_3796, signal_2338}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2324 ( .a ({signal_7028, signal_7022}), .b ({signal_3777, signal_2319}), .clk ( clk ), .r ( Fresh[821] ), .c ({signal_3797, signal_2339}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2326 ( .a ({signal_7036, signal_7032}), .b ({signal_3772, signal_2314}), .clk ( clk ), .r ( Fresh[822] ), .c ({signal_3799, signal_2341}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2328 ( .a ({signal_7048, signal_7042}), .b ({signal_3778, signal_2320}), .clk ( clk ), .r ( Fresh[823] ), .c ({signal_3801, signal_2343}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2329 ( .a ({signal_7052, signal_7050}), .b ({signal_3779, signal_2321}), .clk ( clk ), .r ( Fresh[824] ), .c ({signal_3802, signal_2344}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2330 ( .a ({signal_7060, signal_7056}), .b ({signal_3774, signal_2316}), .clk ( clk ), .r ( Fresh[825] ), .c ({signal_3803, signal_2345}) ) ;
    buf_clk cell_4706 ( .C ( clk ), .D ( signal_7065 ), .Q ( signal_7066 ) ) ;
    buf_clk cell_4712 ( .C ( clk ), .D ( signal_7071 ), .Q ( signal_7072 ) ) ;
    buf_clk cell_4720 ( .C ( clk ), .D ( signal_7079 ), .Q ( signal_7080 ) ) ;
    buf_clk cell_4728 ( .C ( clk ), .D ( signal_7087 ), .Q ( signal_7088 ) ) ;
    buf_clk cell_4734 ( .C ( clk ), .D ( signal_7093 ), .Q ( signal_7094 ) ) ;
    buf_clk cell_4740 ( .C ( clk ), .D ( signal_7099 ), .Q ( signal_7100 ) ) ;
    buf_clk cell_4750 ( .C ( clk ), .D ( signal_7109 ), .Q ( signal_7110 ) ) ;
    buf_clk cell_4760 ( .C ( clk ), .D ( signal_7119 ), .Q ( signal_7120 ) ) ;
    buf_clk cell_4766 ( .C ( clk ), .D ( signal_7125 ), .Q ( signal_7126 ) ) ;
    buf_clk cell_4772 ( .C ( clk ), .D ( signal_7131 ), .Q ( signal_7132 ) ) ;
    buf_clk cell_4776 ( .C ( clk ), .D ( signal_7135 ), .Q ( signal_7136 ) ) ;
    buf_clk cell_4780 ( .C ( clk ), .D ( signal_7139 ), .Q ( signal_7140 ) ) ;
    buf_clk cell_4788 ( .C ( clk ), .D ( signal_7147 ), .Q ( signal_7148 ) ) ;
    buf_clk cell_4796 ( .C ( clk ), .D ( signal_7155 ), .Q ( signal_7156 ) ) ;
    buf_clk cell_4802 ( .C ( clk ), .D ( signal_7161 ), .Q ( signal_7162 ) ) ;
    buf_clk cell_4808 ( .C ( clk ), .D ( signal_7167 ), .Q ( signal_7168 ) ) ;
    buf_clk cell_4816 ( .C ( clk ), .D ( signal_7175 ), .Q ( signal_7176 ) ) ;
    buf_clk cell_4824 ( .C ( clk ), .D ( signal_7183 ), .Q ( signal_7184 ) ) ;
    buf_clk cell_4830 ( .C ( clk ), .D ( signal_7189 ), .Q ( signal_7190 ) ) ;
    buf_clk cell_4836 ( .C ( clk ), .D ( signal_7195 ), .Q ( signal_7196 ) ) ;
    buf_clk cell_4844 ( .C ( clk ), .D ( signal_7203 ), .Q ( signal_7204 ) ) ;
    buf_clk cell_4852 ( .C ( clk ), .D ( signal_7211 ), .Q ( signal_7212 ) ) ;
    buf_clk cell_4856 ( .C ( clk ), .D ( signal_7215 ), .Q ( signal_7216 ) ) ;
    buf_clk cell_4860 ( .C ( clk ), .D ( signal_7219 ), .Q ( signal_7220 ) ) ;
    buf_clk cell_4866 ( .C ( clk ), .D ( signal_7225 ), .Q ( signal_7226 ) ) ;
    buf_clk cell_4872 ( .C ( clk ), .D ( signal_7231 ), .Q ( signal_7232 ) ) ;
    buf_clk cell_4878 ( .C ( clk ), .D ( signal_7237 ), .Q ( signal_7238 ) ) ;
    buf_clk cell_4884 ( .C ( clk ), .D ( signal_7243 ), .Q ( signal_7244 ) ) ;
    buf_clk cell_4888 ( .C ( clk ), .D ( signal_7247 ), .Q ( signal_7248 ) ) ;
    buf_clk cell_4892 ( .C ( clk ), .D ( signal_7251 ), .Q ( signal_7252 ) ) ;
    buf_clk cell_4896 ( .C ( clk ), .D ( signal_7255 ), .Q ( signal_7256 ) ) ;
    buf_clk cell_4900 ( .C ( clk ), .D ( signal_7259 ), .Q ( signal_7260 ) ) ;
    buf_clk cell_4906 ( .C ( clk ), .D ( signal_7265 ), .Q ( signal_7266 ) ) ;
    buf_clk cell_4914 ( .C ( clk ), .D ( signal_7273 ), .Q ( signal_7274 ) ) ;
    buf_clk cell_4926 ( .C ( clk ), .D ( signal_7285 ), .Q ( signal_7286 ) ) ;
    buf_clk cell_4938 ( .C ( clk ), .D ( signal_7297 ), .Q ( signal_7298 ) ) ;
    buf_clk cell_4944 ( .C ( clk ), .D ( signal_7303 ), .Q ( signal_7304 ) ) ;
    buf_clk cell_4950 ( .C ( clk ), .D ( signal_7309 ), .Q ( signal_7310 ) ) ;
    buf_clk cell_4956 ( .C ( clk ), .D ( signal_7315 ), .Q ( signal_7316 ) ) ;
    buf_clk cell_4962 ( .C ( clk ), .D ( signal_7321 ), .Q ( signal_7322 ) ) ;
    buf_clk cell_4976 ( .C ( clk ), .D ( signal_7335 ), .Q ( signal_7336 ) ) ;
    buf_clk cell_4990 ( .C ( clk ), .D ( signal_7349 ), .Q ( signal_7350 ) ) ;
    buf_clk cell_4998 ( .C ( clk ), .D ( signal_7357 ), .Q ( signal_7358 ) ) ;
    buf_clk cell_5006 ( .C ( clk ), .D ( signal_7365 ), .Q ( signal_7366 ) ) ;
    buf_clk cell_5020 ( .C ( clk ), .D ( signal_7379 ), .Q ( signal_7380 ) ) ;
    buf_clk cell_5034 ( .C ( clk ), .D ( signal_7393 ), .Q ( signal_7394 ) ) ;
    buf_clk cell_5042 ( .C ( clk ), .D ( signal_7401 ), .Q ( signal_7402 ) ) ;
    buf_clk cell_5050 ( .C ( clk ), .D ( signal_7409 ), .Q ( signal_7410 ) ) ;
    buf_clk cell_5066 ( .C ( clk ), .D ( signal_7425 ), .Q ( signal_7426 ) ) ;
    buf_clk cell_5076 ( .C ( clk ), .D ( signal_7435 ), .Q ( signal_7436 ) ) ;
    buf_clk cell_5100 ( .C ( clk ), .D ( signal_7459 ), .Q ( signal_7460 ) ) ;
    buf_clk cell_5116 ( .C ( clk ), .D ( signal_7475 ), .Q ( signal_7476 ) ) ;
    buf_clk cell_5140 ( .C ( clk ), .D ( signal_7499 ), .Q ( signal_7500 ) ) ;
    buf_clk cell_5156 ( .C ( clk ), .D ( signal_7515 ), .Q ( signal_7516 ) ) ;
    buf_clk cell_5166 ( .C ( clk ), .D ( signal_7525 ), .Q ( signal_7526 ) ) ;
    buf_clk cell_5176 ( .C ( clk ), .D ( signal_7535 ), .Q ( signal_7536 ) ) ;
    buf_clk cell_5204 ( .C ( clk ), .D ( signal_7563 ), .Q ( signal_7564 ) ) ;
    buf_clk cell_5214 ( .C ( clk ), .D ( signal_7573 ), .Q ( signal_7574 ) ) ;
    buf_clk cell_5236 ( .C ( clk ), .D ( signal_7595 ), .Q ( signal_7596 ) ) ;
    buf_clk cell_5246 ( .C ( clk ), .D ( signal_7605 ), .Q ( signal_7606 ) ) ;
    buf_clk cell_5262 ( .C ( clk ), .D ( signal_7621 ), .Q ( signal_7622 ) ) ;
    buf_clk cell_5278 ( .C ( clk ), .D ( signal_7637 ), .Q ( signal_7638 ) ) ;
    buf_clk cell_5296 ( .C ( clk ), .D ( signal_7655 ), .Q ( signal_7656 ) ) ;
    buf_clk cell_5314 ( .C ( clk ), .D ( signal_7673 ), .Q ( signal_7674 ) ) ;
    buf_clk cell_5330 ( .C ( clk ), .D ( signal_7689 ), .Q ( signal_7690 ) ) ;
    buf_clk cell_5338 ( .C ( clk ), .D ( signal_7697 ), .Q ( signal_7698 ) ) ;
    buf_clk cell_5396 ( .C ( clk ), .D ( signal_7755 ), .Q ( signal_7756 ) ) ;
    buf_clk cell_5416 ( .C ( clk ), .D ( signal_7775 ), .Q ( signal_7776 ) ) ;
    buf_clk cell_5442 ( .C ( clk ), .D ( signal_7801 ), .Q ( signal_7802 ) ) ;
    buf_clk cell_5454 ( .C ( clk ), .D ( signal_7813 ), .Q ( signal_7814 ) ) ;
    buf_clk cell_5466 ( .C ( clk ), .D ( signal_7825 ), .Q ( signal_7826 ) ) ;
    buf_clk cell_5480 ( .C ( clk ), .D ( signal_7839 ), .Q ( signal_7840 ) ) ;

    /* cells in depth 19 */
    buf_clk cell_4907 ( .C ( clk ), .D ( signal_7266 ), .Q ( signal_7267 ) ) ;
    buf_clk cell_4915 ( .C ( clk ), .D ( signal_7274 ), .Q ( signal_7275 ) ) ;
    buf_clk cell_4927 ( .C ( clk ), .D ( signal_7286 ), .Q ( signal_7287 ) ) ;
    buf_clk cell_4939 ( .C ( clk ), .D ( signal_7298 ), .Q ( signal_7299 ) ) ;
    buf_clk cell_4945 ( .C ( clk ), .D ( signal_7304 ), .Q ( signal_7305 ) ) ;
    buf_clk cell_4951 ( .C ( clk ), .D ( signal_7310 ), .Q ( signal_7311 ) ) ;
    buf_clk cell_4957 ( .C ( clk ), .D ( signal_7316 ), .Q ( signal_7317 ) ) ;
    buf_clk cell_4963 ( .C ( clk ), .D ( signal_7322 ), .Q ( signal_7323 ) ) ;
    buf_clk cell_4977 ( .C ( clk ), .D ( signal_7336 ), .Q ( signal_7337 ) ) ;
    buf_clk cell_4991 ( .C ( clk ), .D ( signal_7350 ), .Q ( signal_7351 ) ) ;
    buf_clk cell_4999 ( .C ( clk ), .D ( signal_7358 ), .Q ( signal_7359 ) ) ;
    buf_clk cell_5007 ( .C ( clk ), .D ( signal_7366 ), .Q ( signal_7367 ) ) ;
    buf_clk cell_5021 ( .C ( clk ), .D ( signal_7380 ), .Q ( signal_7381 ) ) ;
    buf_clk cell_5035 ( .C ( clk ), .D ( signal_7394 ), .Q ( signal_7395 ) ) ;
    buf_clk cell_5043 ( .C ( clk ), .D ( signal_7402 ), .Q ( signal_7403 ) ) ;
    buf_clk cell_5051 ( .C ( clk ), .D ( signal_7410 ), .Q ( signal_7411 ) ) ;
    buf_clk cell_5053 ( .C ( clk ), .D ( signal_2335 ), .Q ( signal_7413 ) ) ;
    buf_clk cell_5057 ( .C ( clk ), .D ( signal_3793 ), .Q ( signal_7417 ) ) ;
    buf_clk cell_5067 ( .C ( clk ), .D ( signal_7426 ), .Q ( signal_7427 ) ) ;
    buf_clk cell_5077 ( .C ( clk ), .D ( signal_7436 ), .Q ( signal_7437 ) ) ;
    buf_clk cell_5101 ( .C ( clk ), .D ( signal_7460 ), .Q ( signal_7461 ) ) ;
    buf_clk cell_5117 ( .C ( clk ), .D ( signal_7476 ), .Q ( signal_7477 ) ) ;
    buf_clk cell_5121 ( .C ( clk ), .D ( signal_2308 ), .Q ( signal_7481 ) ) ;
    buf_clk cell_5125 ( .C ( clk ), .D ( signal_3766 ), .Q ( signal_7485 ) ) ;
    buf_clk cell_5141 ( .C ( clk ), .D ( signal_7500 ), .Q ( signal_7501 ) ) ;
    buf_clk cell_5157 ( .C ( clk ), .D ( signal_7516 ), .Q ( signal_7517 ) ) ;
    buf_clk cell_5167 ( .C ( clk ), .D ( signal_7526 ), .Q ( signal_7527 ) ) ;
    buf_clk cell_5177 ( .C ( clk ), .D ( signal_7536 ), .Q ( signal_7537 ) ) ;
    buf_clk cell_5181 ( .C ( clk ), .D ( signal_2318 ), .Q ( signal_7541 ) ) ;
    buf_clk cell_5185 ( .C ( clk ), .D ( signal_3776 ), .Q ( signal_7545 ) ) ;
    buf_clk cell_5189 ( .C ( clk ), .D ( signal_2336 ), .Q ( signal_7549 ) ) ;
    buf_clk cell_5195 ( .C ( clk ), .D ( signal_3794 ), .Q ( signal_7555 ) ) ;
    buf_clk cell_5205 ( .C ( clk ), .D ( signal_7564 ), .Q ( signal_7565 ) ) ;
    buf_clk cell_5215 ( .C ( clk ), .D ( signal_7574 ), .Q ( signal_7575 ) ) ;
    buf_clk cell_5221 ( .C ( clk ), .D ( signal_2343 ), .Q ( signal_7581 ) ) ;
    buf_clk cell_5227 ( .C ( clk ), .D ( signal_3801 ), .Q ( signal_7587 ) ) ;
    buf_clk cell_5237 ( .C ( clk ), .D ( signal_7596 ), .Q ( signal_7597 ) ) ;
    buf_clk cell_5247 ( .C ( clk ), .D ( signal_7606 ), .Q ( signal_7607 ) ) ;
    buf_clk cell_5263 ( .C ( clk ), .D ( signal_7622 ), .Q ( signal_7623 ) ) ;
    buf_clk cell_5279 ( .C ( clk ), .D ( signal_7638 ), .Q ( signal_7639 ) ) ;
    buf_clk cell_5297 ( .C ( clk ), .D ( signal_7656 ), .Q ( signal_7657 ) ) ;
    buf_clk cell_5315 ( .C ( clk ), .D ( signal_7674 ), .Q ( signal_7675 ) ) ;
    buf_clk cell_5331 ( .C ( clk ), .D ( signal_7690 ), .Q ( signal_7691 ) ) ;
    buf_clk cell_5339 ( .C ( clk ), .D ( signal_7698 ), .Q ( signal_7699 ) ) ;
    buf_clk cell_5345 ( .C ( clk ), .D ( signal_2306 ), .Q ( signal_7705 ) ) ;
    buf_clk cell_5353 ( .C ( clk ), .D ( signal_3764 ), .Q ( signal_7713 ) ) ;
    buf_clk cell_5397 ( .C ( clk ), .D ( signal_7756 ), .Q ( signal_7757 ) ) ;
    buf_clk cell_5417 ( .C ( clk ), .D ( signal_7776 ), .Q ( signal_7777 ) ) ;
    buf_clk cell_5443 ( .C ( clk ), .D ( signal_7802 ), .Q ( signal_7803 ) ) ;
    buf_clk cell_5455 ( .C ( clk ), .D ( signal_7814 ), .Q ( signal_7815 ) ) ;
    buf_clk cell_5467 ( .C ( clk ), .D ( signal_7826 ), .Q ( signal_7827 ) ) ;
    buf_clk cell_5481 ( .C ( clk ), .D ( signal_7840 ), .Q ( signal_7841 ) ) ;
    buf_clk cell_5493 ( .C ( clk ), .D ( signal_2328 ), .Q ( signal_7853 ) ) ;
    buf_clk cell_5507 ( .C ( clk ), .D ( signal_3786 ), .Q ( signal_7867 ) ) ;

    /* cells in depth 20 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2269 ( .a ({signal_7072, signal_7066}), .b ({signal_3703, signal_2245}), .clk ( clk ), .r ( Fresh[826] ), .c ({signal_3742, signal_2284}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2270 ( .a ({signal_7088, signal_7080}), .b ({signal_3705, signal_2247}), .clk ( clk ), .r ( Fresh[827] ), .c ({signal_3743, signal_2285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2296 ( .a ({signal_7100, signal_7094}), .b ({signal_3740, signal_2282}), .clk ( clk ), .r ( Fresh[828] ), .c ({signal_3769, signal_2311}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2316 ( .a ({signal_7120, signal_7110}), .b ({signal_3765, signal_2307}), .clk ( clk ), .r ( Fresh[829] ), .c ({signal_3789, signal_2331}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2317 ( .a ({signal_7132, signal_7126}), .b ({signal_3754, signal_2296}), .clk ( clk ), .r ( Fresh[830] ), .c ({signal_3790, signal_2332}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2318 ( .a ({signal_7140, signal_7136}), .b ({signal_3704, signal_2246}), .clk ( clk ), .r ( Fresh[831] ), .c ({signal_3791, signal_2333}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2325 ( .a ({signal_7156, signal_7148}), .b ({signal_3771, signal_2313}), .clk ( clk ), .r ( Fresh[832] ), .c ({signal_3798, signal_2340}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2327 ( .a ({signal_7168, signal_7162}), .b ({signal_3773, signal_2315}), .clk ( clk ), .r ( Fresh[833] ), .c ({signal_3800, signal_2342}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2331 ( .a ({signal_7184, signal_7176}), .b ({signal_3785, signal_2327}), .clk ( clk ), .r ( Fresh[834] ), .c ({signal_3804, signal_2346}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2332 ( .a ({signal_7196, signal_7190}), .b ({signal_3775, signal_2317}), .clk ( clk ), .r ( Fresh[835] ), .c ({signal_3805, signal_2347}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2333 ( .a ({signal_7212, signal_7204}), .b ({signal_3787, signal_2329}), .clk ( clk ), .r ( Fresh[836] ), .c ({signal_3806, signal_2348}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2335 ( .a ({signal_3798, signal_2340}), .b ({signal_3808, signal_2350}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2336 ( .a ({signal_3805, signal_2347}), .b ({signal_3809, signal_2351}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2337 ( .a ({signal_7220, signal_7216}), .b ({signal_3799, signal_2341}), .clk ( clk ), .r ( Fresh[837] ), .c ({signal_3810, signal_2352}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2339 ( .a ({signal_7232, signal_7226}), .b ({signal_3802, signal_2344}), .clk ( clk ), .r ( Fresh[838] ), .c ({signal_3812, signal_2354}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2340 ( .a ({signal_7244, signal_7238}), .b ({signal_3795, signal_2337}), .clk ( clk ), .r ( Fresh[839] ), .c ({signal_3813, signal_2355}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2341 ( .a ({signal_7252, signal_7248}), .b ({signal_3796, signal_2338}), .clk ( clk ), .r ( Fresh[840] ), .c ({signal_3814, signal_2356}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2342 ( .a ({signal_7260, signal_7256}), .b ({signal_3803, signal_2345}), .clk ( clk ), .r ( Fresh[841] ), .c ({signal_3815, signal_2357}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2343 ( .a ({signal_3797, signal_2339}), .b ({signal_3788, signal_2330}), .clk ( clk ), .r ( Fresh[842] ), .c ({signal_3816, signal_2358}) ) ;
    buf_clk cell_4908 ( .C ( clk ), .D ( signal_7267 ), .Q ( signal_7268 ) ) ;
    buf_clk cell_4916 ( .C ( clk ), .D ( signal_7275 ), .Q ( signal_7276 ) ) ;
    buf_clk cell_4928 ( .C ( clk ), .D ( signal_7287 ), .Q ( signal_7288 ) ) ;
    buf_clk cell_4940 ( .C ( clk ), .D ( signal_7299 ), .Q ( signal_7300 ) ) ;
    buf_clk cell_4946 ( .C ( clk ), .D ( signal_7305 ), .Q ( signal_7306 ) ) ;
    buf_clk cell_4952 ( .C ( clk ), .D ( signal_7311 ), .Q ( signal_7312 ) ) ;
    buf_clk cell_4958 ( .C ( clk ), .D ( signal_7317 ), .Q ( signal_7318 ) ) ;
    buf_clk cell_4964 ( .C ( clk ), .D ( signal_7323 ), .Q ( signal_7324 ) ) ;
    buf_clk cell_4978 ( .C ( clk ), .D ( signal_7337 ), .Q ( signal_7338 ) ) ;
    buf_clk cell_4992 ( .C ( clk ), .D ( signal_7351 ), .Q ( signal_7352 ) ) ;
    buf_clk cell_5000 ( .C ( clk ), .D ( signal_7359 ), .Q ( signal_7360 ) ) ;
    buf_clk cell_5008 ( .C ( clk ), .D ( signal_7367 ), .Q ( signal_7368 ) ) ;
    buf_clk cell_5022 ( .C ( clk ), .D ( signal_7381 ), .Q ( signal_7382 ) ) ;
    buf_clk cell_5036 ( .C ( clk ), .D ( signal_7395 ), .Q ( signal_7396 ) ) ;
    buf_clk cell_5044 ( .C ( clk ), .D ( signal_7403 ), .Q ( signal_7404 ) ) ;
    buf_clk cell_5052 ( .C ( clk ), .D ( signal_7411 ), .Q ( signal_7412 ) ) ;
    buf_clk cell_5054 ( .C ( clk ), .D ( signal_7413 ), .Q ( signal_7414 ) ) ;
    buf_clk cell_5058 ( .C ( clk ), .D ( signal_7417 ), .Q ( signal_7418 ) ) ;
    buf_clk cell_5068 ( .C ( clk ), .D ( signal_7427 ), .Q ( signal_7428 ) ) ;
    buf_clk cell_5078 ( .C ( clk ), .D ( signal_7437 ), .Q ( signal_7438 ) ) ;
    buf_clk cell_5102 ( .C ( clk ), .D ( signal_7461 ), .Q ( signal_7462 ) ) ;
    buf_clk cell_5118 ( .C ( clk ), .D ( signal_7477 ), .Q ( signal_7478 ) ) ;
    buf_clk cell_5122 ( .C ( clk ), .D ( signal_7481 ), .Q ( signal_7482 ) ) ;
    buf_clk cell_5126 ( .C ( clk ), .D ( signal_7485 ), .Q ( signal_7486 ) ) ;
    buf_clk cell_5142 ( .C ( clk ), .D ( signal_7501 ), .Q ( signal_7502 ) ) ;
    buf_clk cell_5158 ( .C ( clk ), .D ( signal_7517 ), .Q ( signal_7518 ) ) ;
    buf_clk cell_5168 ( .C ( clk ), .D ( signal_7527 ), .Q ( signal_7528 ) ) ;
    buf_clk cell_5178 ( .C ( clk ), .D ( signal_7537 ), .Q ( signal_7538 ) ) ;
    buf_clk cell_5182 ( .C ( clk ), .D ( signal_7541 ), .Q ( signal_7542 ) ) ;
    buf_clk cell_5186 ( .C ( clk ), .D ( signal_7545 ), .Q ( signal_7546 ) ) ;
    buf_clk cell_5190 ( .C ( clk ), .D ( signal_7549 ), .Q ( signal_7550 ) ) ;
    buf_clk cell_5196 ( .C ( clk ), .D ( signal_7555 ), .Q ( signal_7556 ) ) ;
    buf_clk cell_5206 ( .C ( clk ), .D ( signal_7565 ), .Q ( signal_7566 ) ) ;
    buf_clk cell_5216 ( .C ( clk ), .D ( signal_7575 ), .Q ( signal_7576 ) ) ;
    buf_clk cell_5222 ( .C ( clk ), .D ( signal_7581 ), .Q ( signal_7582 ) ) ;
    buf_clk cell_5228 ( .C ( clk ), .D ( signal_7587 ), .Q ( signal_7588 ) ) ;
    buf_clk cell_5238 ( .C ( clk ), .D ( signal_7597 ), .Q ( signal_7598 ) ) ;
    buf_clk cell_5248 ( .C ( clk ), .D ( signal_7607 ), .Q ( signal_7608 ) ) ;
    buf_clk cell_5264 ( .C ( clk ), .D ( signal_7623 ), .Q ( signal_7624 ) ) ;
    buf_clk cell_5280 ( .C ( clk ), .D ( signal_7639 ), .Q ( signal_7640 ) ) ;
    buf_clk cell_5298 ( .C ( clk ), .D ( signal_7657 ), .Q ( signal_7658 ) ) ;
    buf_clk cell_5316 ( .C ( clk ), .D ( signal_7675 ), .Q ( signal_7676 ) ) ;
    buf_clk cell_5332 ( .C ( clk ), .D ( signal_7691 ), .Q ( signal_7692 ) ) ;
    buf_clk cell_5340 ( .C ( clk ), .D ( signal_7699 ), .Q ( signal_7700 ) ) ;
    buf_clk cell_5346 ( .C ( clk ), .D ( signal_7705 ), .Q ( signal_7706 ) ) ;
    buf_clk cell_5354 ( .C ( clk ), .D ( signal_7713 ), .Q ( signal_7714 ) ) ;
    buf_clk cell_5398 ( .C ( clk ), .D ( signal_7757 ), .Q ( signal_7758 ) ) ;
    buf_clk cell_5418 ( .C ( clk ), .D ( signal_7777 ), .Q ( signal_7778 ) ) ;
    buf_clk cell_5444 ( .C ( clk ), .D ( signal_7803 ), .Q ( signal_7804 ) ) ;
    buf_clk cell_5456 ( .C ( clk ), .D ( signal_7815 ), .Q ( signal_7816 ) ) ;
    buf_clk cell_5468 ( .C ( clk ), .D ( signal_7827 ), .Q ( signal_7828 ) ) ;
    buf_clk cell_5482 ( .C ( clk ), .D ( signal_7841 ), .Q ( signal_7842 ) ) ;
    buf_clk cell_5494 ( .C ( clk ), .D ( signal_7853 ), .Q ( signal_7854 ) ) ;
    buf_clk cell_5508 ( .C ( clk ), .D ( signal_7867 ), .Q ( signal_7868 ) ) ;

    /* cells in depth 21 */
    buf_clk cell_5055 ( .C ( clk ), .D ( signal_7414 ), .Q ( signal_7415 ) ) ;
    buf_clk cell_5059 ( .C ( clk ), .D ( signal_7418 ), .Q ( signal_7419 ) ) ;
    buf_clk cell_5069 ( .C ( clk ), .D ( signal_7428 ), .Q ( signal_7429 ) ) ;
    buf_clk cell_5079 ( .C ( clk ), .D ( signal_7438 ), .Q ( signal_7439 ) ) ;
    buf_clk cell_5081 ( .C ( clk ), .D ( signal_2354 ), .Q ( signal_7441 ) ) ;
    buf_clk cell_5083 ( .C ( clk ), .D ( signal_3812 ), .Q ( signal_7443 ) ) ;
    buf_clk cell_5085 ( .C ( clk ), .D ( signal_2357 ), .Q ( signal_7445 ) ) ;
    buf_clk cell_5087 ( .C ( clk ), .D ( signal_3815 ), .Q ( signal_7447 ) ) ;
    buf_clk cell_5103 ( .C ( clk ), .D ( signal_7462 ), .Q ( signal_7463 ) ) ;
    buf_clk cell_5119 ( .C ( clk ), .D ( signal_7478 ), .Q ( signal_7479 ) ) ;
    buf_clk cell_5123 ( .C ( clk ), .D ( signal_7482 ), .Q ( signal_7483 ) ) ;
    buf_clk cell_5127 ( .C ( clk ), .D ( signal_7486 ), .Q ( signal_7487 ) ) ;
    buf_clk cell_5143 ( .C ( clk ), .D ( signal_7502 ), .Q ( signal_7503 ) ) ;
    buf_clk cell_5159 ( .C ( clk ), .D ( signal_7518 ), .Q ( signal_7519 ) ) ;
    buf_clk cell_5169 ( .C ( clk ), .D ( signal_7528 ), .Q ( signal_7529 ) ) ;
    buf_clk cell_5179 ( .C ( clk ), .D ( signal_7538 ), .Q ( signal_7539 ) ) ;
    buf_clk cell_5183 ( .C ( clk ), .D ( signal_7542 ), .Q ( signal_7543 ) ) ;
    buf_clk cell_5187 ( .C ( clk ), .D ( signal_7546 ), .Q ( signal_7547 ) ) ;
    buf_clk cell_5191 ( .C ( clk ), .D ( signal_7550 ), .Q ( signal_7551 ) ) ;
    buf_clk cell_5197 ( .C ( clk ), .D ( signal_7556 ), .Q ( signal_7557 ) ) ;
    buf_clk cell_5207 ( .C ( clk ), .D ( signal_7566 ), .Q ( signal_7567 ) ) ;
    buf_clk cell_5217 ( .C ( clk ), .D ( signal_7576 ), .Q ( signal_7577 ) ) ;
    buf_clk cell_5223 ( .C ( clk ), .D ( signal_7582 ), .Q ( signal_7583 ) ) ;
    buf_clk cell_5229 ( .C ( clk ), .D ( signal_7588 ), .Q ( signal_7589 ) ) ;
    buf_clk cell_5239 ( .C ( clk ), .D ( signal_7598 ), .Q ( signal_7599 ) ) ;
    buf_clk cell_5249 ( .C ( clk ), .D ( signal_7608 ), .Q ( signal_7609 ) ) ;
    buf_clk cell_5265 ( .C ( clk ), .D ( signal_7624 ), .Q ( signal_7625 ) ) ;
    buf_clk cell_5281 ( .C ( clk ), .D ( signal_7640 ), .Q ( signal_7641 ) ) ;
    buf_clk cell_5299 ( .C ( clk ), .D ( signal_7658 ), .Q ( signal_7659 ) ) ;
    buf_clk cell_5317 ( .C ( clk ), .D ( signal_7676 ), .Q ( signal_7677 ) ) ;
    buf_clk cell_5321 ( .C ( clk ), .D ( signal_2348 ), .Q ( signal_7681 ) ) ;
    buf_clk cell_5325 ( .C ( clk ), .D ( signal_3806 ), .Q ( signal_7685 ) ) ;
    buf_clk cell_5333 ( .C ( clk ), .D ( signal_7692 ), .Q ( signal_7693 ) ) ;
    buf_clk cell_5341 ( .C ( clk ), .D ( signal_7700 ), .Q ( signal_7701 ) ) ;
    buf_clk cell_5347 ( .C ( clk ), .D ( signal_7706 ), .Q ( signal_7707 ) ) ;
    buf_clk cell_5355 ( .C ( clk ), .D ( signal_7714 ), .Q ( signal_7715 ) ) ;
    buf_clk cell_5361 ( .C ( clk ), .D ( signal_2285 ), .Q ( signal_7721 ) ) ;
    buf_clk cell_5367 ( .C ( clk ), .D ( signal_3743 ), .Q ( signal_7727 ) ) ;
    buf_clk cell_5399 ( .C ( clk ), .D ( signal_7758 ), .Q ( signal_7759 ) ) ;
    buf_clk cell_5419 ( .C ( clk ), .D ( signal_7778 ), .Q ( signal_7779 ) ) ;
    buf_clk cell_5425 ( .C ( clk ), .D ( signal_2332 ), .Q ( signal_7785 ) ) ;
    buf_clk cell_5433 ( .C ( clk ), .D ( signal_3790 ), .Q ( signal_7793 ) ) ;
    buf_clk cell_5445 ( .C ( clk ), .D ( signal_7804 ), .Q ( signal_7805 ) ) ;
    buf_clk cell_5457 ( .C ( clk ), .D ( signal_7816 ), .Q ( signal_7817 ) ) ;
    buf_clk cell_5469 ( .C ( clk ), .D ( signal_7828 ), .Q ( signal_7829 ) ) ;
    buf_clk cell_5483 ( .C ( clk ), .D ( signal_7842 ), .Q ( signal_7843 ) ) ;
    buf_clk cell_5495 ( .C ( clk ), .D ( signal_7854 ), .Q ( signal_7855 ) ) ;
    buf_clk cell_5509 ( .C ( clk ), .D ( signal_7868 ), .Q ( signal_7869 ) ) ;

    /* cells in depth 22 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2319 ( .a ({signal_7276, signal_7268}), .b ({signal_3769, signal_2311}), .clk ( clk ), .r ( Fresh[843] ), .c ({signal_3792, signal_2334}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2334 ( .a ({signal_7300, signal_7288}), .b ({signal_3789, signal_2331}), .clk ( clk ), .r ( Fresh[844] ), .c ({signal_3807, signal_2349}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2338 ( .a ({signal_7312, signal_7306}), .b ({signal_3800, signal_2342}), .clk ( clk ), .r ( Fresh[845] ), .c ({signal_3811, signal_2353}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2344 ( .a ({signal_3804, signal_2346}), .b ({signal_3742, signal_2284}), .clk ( clk ), .r ( Fresh[846] ), .c ({signal_3817, signal_2359}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2346 ( .a ({signal_7324, signal_7318}), .b ({signal_3808, signal_2350}), .clk ( clk ), .r ( Fresh[847] ), .c ({signal_3819, signal_2361}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2348 ( .a ({signal_7352, signal_7338}), .b ({signal_3813, signal_2355}), .clk ( clk ), .r ( Fresh[848] ), .c ({signal_3821, signal_2363}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2349 ( .a ({signal_7368, signal_7360}), .b ({signal_3814, signal_2356}), .clk ( clk ), .r ( Fresh[849] ), .c ({signal_3822, signal_2364}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2350 ( .a ({signal_7396, signal_7382}), .b ({signal_3809, signal_2351}), .clk ( clk ), .r ( Fresh[850] ), .c ({signal_3823, signal_2365}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2351 ( .a ({signal_7412, signal_7404}), .b ({signal_3816, signal_2358}), .clk ( clk ), .r ( Fresh[851] ), .c ({signal_3824, signal_2366}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2352 ( .a ({signal_3810, signal_2352}), .b ({signal_3791, signal_2333}), .clk ( clk ), .r ( Fresh[852] ), .c ({signal_3825, signal_2367}) ) ;
    buf_clk cell_5056 ( .C ( clk ), .D ( signal_7415 ), .Q ( signal_7416 ) ) ;
    buf_clk cell_5060 ( .C ( clk ), .D ( signal_7419 ), .Q ( signal_7420 ) ) ;
    buf_clk cell_5070 ( .C ( clk ), .D ( signal_7429 ), .Q ( signal_7430 ) ) ;
    buf_clk cell_5080 ( .C ( clk ), .D ( signal_7439 ), .Q ( signal_7440 ) ) ;
    buf_clk cell_5082 ( .C ( clk ), .D ( signal_7441 ), .Q ( signal_7442 ) ) ;
    buf_clk cell_5084 ( .C ( clk ), .D ( signal_7443 ), .Q ( signal_7444 ) ) ;
    buf_clk cell_5086 ( .C ( clk ), .D ( signal_7445 ), .Q ( signal_7446 ) ) ;
    buf_clk cell_5088 ( .C ( clk ), .D ( signal_7447 ), .Q ( signal_7448 ) ) ;
    buf_clk cell_5104 ( .C ( clk ), .D ( signal_7463 ), .Q ( signal_7464 ) ) ;
    buf_clk cell_5120 ( .C ( clk ), .D ( signal_7479 ), .Q ( signal_7480 ) ) ;
    buf_clk cell_5124 ( .C ( clk ), .D ( signal_7483 ), .Q ( signal_7484 ) ) ;
    buf_clk cell_5128 ( .C ( clk ), .D ( signal_7487 ), .Q ( signal_7488 ) ) ;
    buf_clk cell_5144 ( .C ( clk ), .D ( signal_7503 ), .Q ( signal_7504 ) ) ;
    buf_clk cell_5160 ( .C ( clk ), .D ( signal_7519 ), .Q ( signal_7520 ) ) ;
    buf_clk cell_5170 ( .C ( clk ), .D ( signal_7529 ), .Q ( signal_7530 ) ) ;
    buf_clk cell_5180 ( .C ( clk ), .D ( signal_7539 ), .Q ( signal_7540 ) ) ;
    buf_clk cell_5184 ( .C ( clk ), .D ( signal_7543 ), .Q ( signal_7544 ) ) ;
    buf_clk cell_5188 ( .C ( clk ), .D ( signal_7547 ), .Q ( signal_7548 ) ) ;
    buf_clk cell_5192 ( .C ( clk ), .D ( signal_7551 ), .Q ( signal_7552 ) ) ;
    buf_clk cell_5198 ( .C ( clk ), .D ( signal_7557 ), .Q ( signal_7558 ) ) ;
    buf_clk cell_5208 ( .C ( clk ), .D ( signal_7567 ), .Q ( signal_7568 ) ) ;
    buf_clk cell_5218 ( .C ( clk ), .D ( signal_7577 ), .Q ( signal_7578 ) ) ;
    buf_clk cell_5224 ( .C ( clk ), .D ( signal_7583 ), .Q ( signal_7584 ) ) ;
    buf_clk cell_5230 ( .C ( clk ), .D ( signal_7589 ), .Q ( signal_7590 ) ) ;
    buf_clk cell_5240 ( .C ( clk ), .D ( signal_7599 ), .Q ( signal_7600 ) ) ;
    buf_clk cell_5250 ( .C ( clk ), .D ( signal_7609 ), .Q ( signal_7610 ) ) ;
    buf_clk cell_5266 ( .C ( clk ), .D ( signal_7625 ), .Q ( signal_7626 ) ) ;
    buf_clk cell_5282 ( .C ( clk ), .D ( signal_7641 ), .Q ( signal_7642 ) ) ;
    buf_clk cell_5300 ( .C ( clk ), .D ( signal_7659 ), .Q ( signal_7660 ) ) ;
    buf_clk cell_5318 ( .C ( clk ), .D ( signal_7677 ), .Q ( signal_7678 ) ) ;
    buf_clk cell_5322 ( .C ( clk ), .D ( signal_7681 ), .Q ( signal_7682 ) ) ;
    buf_clk cell_5326 ( .C ( clk ), .D ( signal_7685 ), .Q ( signal_7686 ) ) ;
    buf_clk cell_5334 ( .C ( clk ), .D ( signal_7693 ), .Q ( signal_7694 ) ) ;
    buf_clk cell_5342 ( .C ( clk ), .D ( signal_7701 ), .Q ( signal_7702 ) ) ;
    buf_clk cell_5348 ( .C ( clk ), .D ( signal_7707 ), .Q ( signal_7708 ) ) ;
    buf_clk cell_5356 ( .C ( clk ), .D ( signal_7715 ), .Q ( signal_7716 ) ) ;
    buf_clk cell_5362 ( .C ( clk ), .D ( signal_7721 ), .Q ( signal_7722 ) ) ;
    buf_clk cell_5368 ( .C ( clk ), .D ( signal_7727 ), .Q ( signal_7728 ) ) ;
    buf_clk cell_5400 ( .C ( clk ), .D ( signal_7759 ), .Q ( signal_7760 ) ) ;
    buf_clk cell_5420 ( .C ( clk ), .D ( signal_7779 ), .Q ( signal_7780 ) ) ;
    buf_clk cell_5426 ( .C ( clk ), .D ( signal_7785 ), .Q ( signal_7786 ) ) ;
    buf_clk cell_5434 ( .C ( clk ), .D ( signal_7793 ), .Q ( signal_7794 ) ) ;
    buf_clk cell_5446 ( .C ( clk ), .D ( signal_7805 ), .Q ( signal_7806 ) ) ;
    buf_clk cell_5458 ( .C ( clk ), .D ( signal_7817 ), .Q ( signal_7818 ) ) ;
    buf_clk cell_5470 ( .C ( clk ), .D ( signal_7829 ), .Q ( signal_7830 ) ) ;
    buf_clk cell_5484 ( .C ( clk ), .D ( signal_7843 ), .Q ( signal_7844 ) ) ;
    buf_clk cell_5496 ( .C ( clk ), .D ( signal_7855 ), .Q ( signal_7856 ) ) ;
    buf_clk cell_5510 ( .C ( clk ), .D ( signal_7869 ), .Q ( signal_7870 ) ) ;

    /* cells in depth 23 */
    buf_clk cell_5193 ( .C ( clk ), .D ( signal_7552 ), .Q ( signal_7553 ) ) ;
    buf_clk cell_5199 ( .C ( clk ), .D ( signal_7558 ), .Q ( signal_7559 ) ) ;
    buf_clk cell_5209 ( .C ( clk ), .D ( signal_7568 ), .Q ( signal_7569 ) ) ;
    buf_clk cell_5219 ( .C ( clk ), .D ( signal_7578 ), .Q ( signal_7579 ) ) ;
    buf_clk cell_5225 ( .C ( clk ), .D ( signal_7584 ), .Q ( signal_7585 ) ) ;
    buf_clk cell_5231 ( .C ( clk ), .D ( signal_7590 ), .Q ( signal_7591 ) ) ;
    buf_clk cell_5241 ( .C ( clk ), .D ( signal_7600 ), .Q ( signal_7601 ) ) ;
    buf_clk cell_5251 ( .C ( clk ), .D ( signal_7610 ), .Q ( signal_7611 ) ) ;
    buf_clk cell_5267 ( .C ( clk ), .D ( signal_7626 ), .Q ( signal_7627 ) ) ;
    buf_clk cell_5283 ( .C ( clk ), .D ( signal_7642 ), .Q ( signal_7643 ) ) ;
    buf_clk cell_5301 ( .C ( clk ), .D ( signal_7660 ), .Q ( signal_7661 ) ) ;
    buf_clk cell_5319 ( .C ( clk ), .D ( signal_7678 ), .Q ( signal_7679 ) ) ;
    buf_clk cell_5323 ( .C ( clk ), .D ( signal_7682 ), .Q ( signal_7683 ) ) ;
    buf_clk cell_5327 ( .C ( clk ), .D ( signal_7686 ), .Q ( signal_7687 ) ) ;
    buf_clk cell_5335 ( .C ( clk ), .D ( signal_7694 ), .Q ( signal_7695 ) ) ;
    buf_clk cell_5343 ( .C ( clk ), .D ( signal_7702 ), .Q ( signal_7703 ) ) ;
    buf_clk cell_5349 ( .C ( clk ), .D ( signal_7708 ), .Q ( signal_7709 ) ) ;
    buf_clk cell_5357 ( .C ( clk ), .D ( signal_7716 ), .Q ( signal_7717 ) ) ;
    buf_clk cell_5363 ( .C ( clk ), .D ( signal_7722 ), .Q ( signal_7723 ) ) ;
    buf_clk cell_5369 ( .C ( clk ), .D ( signal_7728 ), .Q ( signal_7729 ) ) ;
    buf_clk cell_5373 ( .C ( clk ), .D ( signal_2361 ), .Q ( signal_7733 ) ) ;
    buf_clk cell_5377 ( .C ( clk ), .D ( signal_3819 ), .Q ( signal_7737 ) ) ;
    buf_clk cell_5401 ( .C ( clk ), .D ( signal_7760 ), .Q ( signal_7761 ) ) ;
    buf_clk cell_5421 ( .C ( clk ), .D ( signal_7780 ), .Q ( signal_7781 ) ) ;
    buf_clk cell_5427 ( .C ( clk ), .D ( signal_7786 ), .Q ( signal_7787 ) ) ;
    buf_clk cell_5435 ( .C ( clk ), .D ( signal_7794 ), .Q ( signal_7795 ) ) ;
    buf_clk cell_5447 ( .C ( clk ), .D ( signal_7806 ), .Q ( signal_7807 ) ) ;
    buf_clk cell_5459 ( .C ( clk ), .D ( signal_7818 ), .Q ( signal_7819 ) ) ;
    buf_clk cell_5471 ( .C ( clk ), .D ( signal_7830 ), .Q ( signal_7831 ) ) ;
    buf_clk cell_5485 ( .C ( clk ), .D ( signal_7844 ), .Q ( signal_7845 ) ) ;
    buf_clk cell_5497 ( .C ( clk ), .D ( signal_7856 ), .Q ( signal_7857 ) ) ;
    buf_clk cell_5511 ( .C ( clk ), .D ( signal_7870 ), .Q ( signal_7871 ) ) ;

    /* cells in depth 24 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2345 ( .a ({signal_7420, signal_7416}), .b ({signal_3792, signal_2334}), .clk ( clk ), .r ( Fresh[853] ), .c ({signal_3818, signal_2360}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2347 ( .a ({signal_7440, signal_7430}), .b ({signal_3811, signal_2353}), .clk ( clk ), .r ( Fresh[854] ), .c ({signal_3820, signal_2362}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2353 ( .a ({signal_7444, signal_7442}), .b ({signal_3807, signal_2349}), .clk ( clk ), .r ( Fresh[855] ), .c ({signal_3826, signal_2368}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2354 ( .a ({signal_7448, signal_7446}), .b ({signal_3817, signal_2359}), .clk ( clk ), .r ( Fresh[856] ), .c ({signal_3827, signal_2369}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2357 ( .a ({signal_7480, signal_7464}), .b ({signal_3821, signal_2363}), .clk ( clk ), .r ( Fresh[857] ), .c ({signal_3830, signal_2372}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2358 ( .a ({signal_7488, signal_7484}), .b ({signal_3822, signal_2364}), .clk ( clk ), .r ( Fresh[858] ), .c ({signal_3831, signal_2373}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2359 ( .a ({signal_7520, signal_7504}), .b ({signal_3823, signal_2365}), .clk ( clk ), .r ( Fresh[859] ), .c ({signal_3832, signal_2374}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2360 ( .a ({signal_7540, signal_7530}), .b ({signal_3824, signal_2366}), .clk ( clk ), .r ( Fresh[860] ), .c ({signal_3833, signal_2375}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2361 ( .a ({signal_7548, signal_7544}), .b ({signal_3825, signal_2367}), .clk ( clk ), .r ( Fresh[861] ), .c ({signal_3834, signal_2376}) ) ;
    buf_clk cell_5194 ( .C ( clk ), .D ( signal_7553 ), .Q ( signal_7554 ) ) ;
    buf_clk cell_5200 ( .C ( clk ), .D ( signal_7559 ), .Q ( signal_7560 ) ) ;
    buf_clk cell_5210 ( .C ( clk ), .D ( signal_7569 ), .Q ( signal_7570 ) ) ;
    buf_clk cell_5220 ( .C ( clk ), .D ( signal_7579 ), .Q ( signal_7580 ) ) ;
    buf_clk cell_5226 ( .C ( clk ), .D ( signal_7585 ), .Q ( signal_7586 ) ) ;
    buf_clk cell_5232 ( .C ( clk ), .D ( signal_7591 ), .Q ( signal_7592 ) ) ;
    buf_clk cell_5242 ( .C ( clk ), .D ( signal_7601 ), .Q ( signal_7602 ) ) ;
    buf_clk cell_5252 ( .C ( clk ), .D ( signal_7611 ), .Q ( signal_7612 ) ) ;
    buf_clk cell_5268 ( .C ( clk ), .D ( signal_7627 ), .Q ( signal_7628 ) ) ;
    buf_clk cell_5284 ( .C ( clk ), .D ( signal_7643 ), .Q ( signal_7644 ) ) ;
    buf_clk cell_5302 ( .C ( clk ), .D ( signal_7661 ), .Q ( signal_7662 ) ) ;
    buf_clk cell_5320 ( .C ( clk ), .D ( signal_7679 ), .Q ( signal_7680 ) ) ;
    buf_clk cell_5324 ( .C ( clk ), .D ( signal_7683 ), .Q ( signal_7684 ) ) ;
    buf_clk cell_5328 ( .C ( clk ), .D ( signal_7687 ), .Q ( signal_7688 ) ) ;
    buf_clk cell_5336 ( .C ( clk ), .D ( signal_7695 ), .Q ( signal_7696 ) ) ;
    buf_clk cell_5344 ( .C ( clk ), .D ( signal_7703 ), .Q ( signal_7704 ) ) ;
    buf_clk cell_5350 ( .C ( clk ), .D ( signal_7709 ), .Q ( signal_7710 ) ) ;
    buf_clk cell_5358 ( .C ( clk ), .D ( signal_7717 ), .Q ( signal_7718 ) ) ;
    buf_clk cell_5364 ( .C ( clk ), .D ( signal_7723 ), .Q ( signal_7724 ) ) ;
    buf_clk cell_5370 ( .C ( clk ), .D ( signal_7729 ), .Q ( signal_7730 ) ) ;
    buf_clk cell_5374 ( .C ( clk ), .D ( signal_7733 ), .Q ( signal_7734 ) ) ;
    buf_clk cell_5378 ( .C ( clk ), .D ( signal_7737 ), .Q ( signal_7738 ) ) ;
    buf_clk cell_5402 ( .C ( clk ), .D ( signal_7761 ), .Q ( signal_7762 ) ) ;
    buf_clk cell_5422 ( .C ( clk ), .D ( signal_7781 ), .Q ( signal_7782 ) ) ;
    buf_clk cell_5428 ( .C ( clk ), .D ( signal_7787 ), .Q ( signal_7788 ) ) ;
    buf_clk cell_5436 ( .C ( clk ), .D ( signal_7795 ), .Q ( signal_7796 ) ) ;
    buf_clk cell_5448 ( .C ( clk ), .D ( signal_7807 ), .Q ( signal_7808 ) ) ;
    buf_clk cell_5460 ( .C ( clk ), .D ( signal_7819 ), .Q ( signal_7820 ) ) ;
    buf_clk cell_5472 ( .C ( clk ), .D ( signal_7831 ), .Q ( signal_7832 ) ) ;
    buf_clk cell_5486 ( .C ( clk ), .D ( signal_7845 ), .Q ( signal_7846 ) ) ;
    buf_clk cell_5498 ( .C ( clk ), .D ( signal_7857 ), .Q ( signal_7858 ) ) ;
    buf_clk cell_5512 ( .C ( clk ), .D ( signal_7871 ), .Q ( signal_7872 ) ) ;

    /* cells in depth 25 */
    buf_clk cell_5351 ( .C ( clk ), .D ( signal_7710 ), .Q ( signal_7711 ) ) ;
    buf_clk cell_5359 ( .C ( clk ), .D ( signal_7718 ), .Q ( signal_7719 ) ) ;
    buf_clk cell_5365 ( .C ( clk ), .D ( signal_7724 ), .Q ( signal_7725 ) ) ;
    buf_clk cell_5371 ( .C ( clk ), .D ( signal_7730 ), .Q ( signal_7731 ) ) ;
    buf_clk cell_5375 ( .C ( clk ), .D ( signal_7734 ), .Q ( signal_7735 ) ) ;
    buf_clk cell_5379 ( .C ( clk ), .D ( signal_7738 ), .Q ( signal_7739 ) ) ;
    buf_clk cell_5381 ( .C ( clk ), .D ( signal_2373 ), .Q ( signal_7741 ) ) ;
    buf_clk cell_5383 ( .C ( clk ), .D ( signal_3831 ), .Q ( signal_7743 ) ) ;
    buf_clk cell_5403 ( .C ( clk ), .D ( signal_7762 ), .Q ( signal_7763 ) ) ;
    buf_clk cell_5423 ( .C ( clk ), .D ( signal_7782 ), .Q ( signal_7783 ) ) ;
    buf_clk cell_5429 ( .C ( clk ), .D ( signal_7788 ), .Q ( signal_7789 ) ) ;
    buf_clk cell_5437 ( .C ( clk ), .D ( signal_7796 ), .Q ( signal_7797 ) ) ;
    buf_clk cell_5449 ( .C ( clk ), .D ( signal_7808 ), .Q ( signal_7809 ) ) ;
    buf_clk cell_5461 ( .C ( clk ), .D ( signal_7820 ), .Q ( signal_7821 ) ) ;
    buf_clk cell_5473 ( .C ( clk ), .D ( signal_7832 ), .Q ( signal_7833 ) ) ;
    buf_clk cell_5487 ( .C ( clk ), .D ( signal_7846 ), .Q ( signal_7847 ) ) ;
    buf_clk cell_5499 ( .C ( clk ), .D ( signal_7858 ), .Q ( signal_7859 ) ) ;
    buf_clk cell_5513 ( .C ( clk ), .D ( signal_7872 ), .Q ( signal_7873 ) ) ;

    /* cells in depth 26 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2355 ( .a ({signal_7560, signal_7554}), .b ({signal_3818, signal_2360}), .clk ( clk ), .r ( Fresh[862] ), .c ({signal_3828, signal_2370}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2356 ( .a ({signal_7580, signal_7570}), .b ({signal_3820, signal_2362}), .clk ( clk ), .r ( Fresh[863] ), .c ({signal_3829, signal_2371}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2362 ( .a ({signal_7592, signal_7586}), .b ({signal_3826, signal_2368}), .clk ( clk ), .r ( Fresh[864] ), .c ({signal_3835, signal_2377}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2363 ( .a ({signal_7612, signal_7602}), .b ({signal_3827, signal_2369}), .clk ( clk ), .r ( Fresh[865] ), .c ({signal_3836, signal_2378}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2365 ( .a ({signal_3836, signal_2378}), .b ({signal_3838, signal_26}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2368 ( .a ({signal_7644, signal_7628}), .b ({signal_3830, signal_2372}), .clk ( clk ), .r ( Fresh[866] ), .c ({signal_3841, signal_2381}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2369 ( .a ({signal_7680, signal_7662}), .b ({signal_3832, signal_2374}), .clk ( clk ), .r ( Fresh[867] ), .c ({signal_3842, signal_2382}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2370 ( .a ({signal_7688, signal_7684}), .b ({signal_3833, signal_2375}), .clk ( clk ), .r ( Fresh[868] ), .c ({signal_3843, signal_2383}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2371 ( .a ({signal_7704, signal_7696}), .b ({signal_3834, signal_2376}), .clk ( clk ), .r ( Fresh[869] ), .c ({signal_3844, signal_2384}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2374 ( .a ({signal_3843, signal_2383}), .b ({signal_3847, signal_28}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2375 ( .a ({signal_3844, signal_2384}), .b ({signal_3848, signal_29}) ) ;
    buf_clk cell_5352 ( .C ( clk ), .D ( signal_7711 ), .Q ( signal_7712 ) ) ;
    buf_clk cell_5360 ( .C ( clk ), .D ( signal_7719 ), .Q ( signal_7720 ) ) ;
    buf_clk cell_5366 ( .C ( clk ), .D ( signal_7725 ), .Q ( signal_7726 ) ) ;
    buf_clk cell_5372 ( .C ( clk ), .D ( signal_7731 ), .Q ( signal_7732 ) ) ;
    buf_clk cell_5376 ( .C ( clk ), .D ( signal_7735 ), .Q ( signal_7736 ) ) ;
    buf_clk cell_5380 ( .C ( clk ), .D ( signal_7739 ), .Q ( signal_7740 ) ) ;
    buf_clk cell_5382 ( .C ( clk ), .D ( signal_7741 ), .Q ( signal_7742 ) ) ;
    buf_clk cell_5384 ( .C ( clk ), .D ( signal_7743 ), .Q ( signal_7744 ) ) ;
    buf_clk cell_5404 ( .C ( clk ), .D ( signal_7763 ), .Q ( signal_7764 ) ) ;
    buf_clk cell_5424 ( .C ( clk ), .D ( signal_7783 ), .Q ( signal_7784 ) ) ;
    buf_clk cell_5430 ( .C ( clk ), .D ( signal_7789 ), .Q ( signal_7790 ) ) ;
    buf_clk cell_5438 ( .C ( clk ), .D ( signal_7797 ), .Q ( signal_7798 ) ) ;
    buf_clk cell_5450 ( .C ( clk ), .D ( signal_7809 ), .Q ( signal_7810 ) ) ;
    buf_clk cell_5462 ( .C ( clk ), .D ( signal_7821 ), .Q ( signal_7822 ) ) ;
    buf_clk cell_5474 ( .C ( clk ), .D ( signal_7833 ), .Q ( signal_7834 ) ) ;
    buf_clk cell_5488 ( .C ( clk ), .D ( signal_7847 ), .Q ( signal_7848 ) ) ;
    buf_clk cell_5500 ( .C ( clk ), .D ( signal_7859 ), .Q ( signal_7860 ) ) ;
    buf_clk cell_5514 ( .C ( clk ), .D ( signal_7873 ), .Q ( signal_7874 ) ) ;

    /* cells in depth 27 */
    buf_clk cell_5431 ( .C ( clk ), .D ( signal_7790 ), .Q ( signal_7791 ) ) ;
    buf_clk cell_5439 ( .C ( clk ), .D ( signal_7798 ), .Q ( signal_7799 ) ) ;
    buf_clk cell_5451 ( .C ( clk ), .D ( signal_7810 ), .Q ( signal_7811 ) ) ;
    buf_clk cell_5463 ( .C ( clk ), .D ( signal_7822 ), .Q ( signal_7823 ) ) ;
    buf_clk cell_5475 ( .C ( clk ), .D ( signal_7834 ), .Q ( signal_7835 ) ) ;
    buf_clk cell_5489 ( .C ( clk ), .D ( signal_7848 ), .Q ( signal_7849 ) ) ;
    buf_clk cell_5501 ( .C ( clk ), .D ( signal_7860 ), .Q ( signal_7861 ) ) ;
    buf_clk cell_5515 ( .C ( clk ), .D ( signal_7874 ), .Q ( signal_7875 ) ) ;
    buf_clk cell_5553 ( .C ( clk ), .D ( signal_26 ), .Q ( signal_7913 ) ) ;
    buf_clk cell_5561 ( .C ( clk ), .D ( signal_3838 ), .Q ( signal_7921 ) ) ;
    buf_clk cell_5569 ( .C ( clk ), .D ( signal_28 ), .Q ( signal_7929 ) ) ;
    buf_clk cell_5577 ( .C ( clk ), .D ( signal_3847 ), .Q ( signal_7937 ) ) ;
    buf_clk cell_5585 ( .C ( clk ), .D ( signal_29 ), .Q ( signal_7945 ) ) ;
    buf_clk cell_5593 ( .C ( clk ), .D ( signal_3848 ), .Q ( signal_7953 ) ) ;

    /* cells in depth 28 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2364 ( .a ({signal_7720, signal_7712}), .b ({signal_3828, signal_2370}), .clk ( clk ), .r ( Fresh[870] ), .c ({signal_3837, signal_2379}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2366 ( .a ({signal_3837, signal_2379}), .b ({signal_3839, signal_23}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2367 ( .a ({signal_7732, signal_7726}), .b ({signal_3829, signal_2371}), .clk ( clk ), .r ( Fresh[871] ), .c ({signal_3840, signal_2380}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2372 ( .a ({signal_7740, signal_7736}), .b ({signal_3835, signal_2377}), .clk ( clk ), .r ( Fresh[872] ), .c ({signal_3845, signal_2385}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2373 ( .a ({signal_3840, signal_2380}), .b ({signal_3846, signal_30}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2376 ( .a ({signal_3845, signal_2385}), .b ({signal_3849, signal_24}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2377 ( .a ({signal_7744, signal_7742}), .b ({signal_3841, signal_2381}), .clk ( clk ), .r ( Fresh[873] ), .c ({signal_3850, signal_2386}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2378 ( .a ({signal_7784, signal_7764}), .b ({signal_3842, signal_2382}), .clk ( clk ), .r ( Fresh[874] ), .c ({signal_3851, signal_2387}) ) ;
    buf_clk cell_5432 ( .C ( clk ), .D ( signal_7791 ), .Q ( signal_7792 ) ) ;
    buf_clk cell_5440 ( .C ( clk ), .D ( signal_7799 ), .Q ( signal_7800 ) ) ;
    buf_clk cell_5452 ( .C ( clk ), .D ( signal_7811 ), .Q ( signal_7812 ) ) ;
    buf_clk cell_5464 ( .C ( clk ), .D ( signal_7823 ), .Q ( signal_7824 ) ) ;
    buf_clk cell_5476 ( .C ( clk ), .D ( signal_7835 ), .Q ( signal_7836 ) ) ;
    buf_clk cell_5490 ( .C ( clk ), .D ( signal_7849 ), .Q ( signal_7850 ) ) ;
    buf_clk cell_5502 ( .C ( clk ), .D ( signal_7861 ), .Q ( signal_7862 ) ) ;
    buf_clk cell_5516 ( .C ( clk ), .D ( signal_7875 ), .Q ( signal_7876 ) ) ;
    buf_clk cell_5554 ( .C ( clk ), .D ( signal_7913 ), .Q ( signal_7914 ) ) ;
    buf_clk cell_5562 ( .C ( clk ), .D ( signal_7921 ), .Q ( signal_7922 ) ) ;
    buf_clk cell_5570 ( .C ( clk ), .D ( signal_7929 ), .Q ( signal_7930 ) ) ;
    buf_clk cell_5578 ( .C ( clk ), .D ( signal_7937 ), .Q ( signal_7938 ) ) ;
    buf_clk cell_5586 ( .C ( clk ), .D ( signal_7945 ), .Q ( signal_7946 ) ) ;
    buf_clk cell_5594 ( .C ( clk ), .D ( signal_7953 ), .Q ( signal_7954 ) ) ;

    /* cells in depth 29 */
    buf_clk cell_5477 ( .C ( clk ), .D ( signal_7836 ), .Q ( signal_7837 ) ) ;
    buf_clk cell_5491 ( .C ( clk ), .D ( signal_7850 ), .Q ( signal_7851 ) ) ;
    buf_clk cell_5503 ( .C ( clk ), .D ( signal_7862 ), .Q ( signal_7863 ) ) ;
    buf_clk cell_5517 ( .C ( clk ), .D ( signal_7876 ), .Q ( signal_7877 ) ) ;
    buf_clk cell_5521 ( .C ( clk ), .D ( signal_23 ), .Q ( signal_7881 ) ) ;
    buf_clk cell_5527 ( .C ( clk ), .D ( signal_3839 ), .Q ( signal_7887 ) ) ;
    buf_clk cell_5533 ( .C ( clk ), .D ( signal_24 ), .Q ( signal_7893 ) ) ;
    buf_clk cell_5539 ( .C ( clk ), .D ( signal_3849 ), .Q ( signal_7899 ) ) ;
    buf_clk cell_5555 ( .C ( clk ), .D ( signal_7914 ), .Q ( signal_7915 ) ) ;
    buf_clk cell_5563 ( .C ( clk ), .D ( signal_7922 ), .Q ( signal_7923 ) ) ;
    buf_clk cell_5571 ( .C ( clk ), .D ( signal_7930 ), .Q ( signal_7931 ) ) ;
    buf_clk cell_5579 ( .C ( clk ), .D ( signal_7938 ), .Q ( signal_7939 ) ) ;
    buf_clk cell_5587 ( .C ( clk ), .D ( signal_7946 ), .Q ( signal_7947 ) ) ;
    buf_clk cell_5595 ( .C ( clk ), .D ( signal_7954 ), .Q ( signal_7955 ) ) ;
    buf_clk cell_5601 ( .C ( clk ), .D ( signal_30 ), .Q ( signal_7961 ) ) ;
    buf_clk cell_5607 ( .C ( clk ), .D ( signal_3846 ), .Q ( signal_7967 ) ) ;

    /* cells in depth 30 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2379 ( .a ({signal_7800, signal_7792}), .b ({signal_3850, signal_2386}), .clk ( clk ), .r ( Fresh[875] ), .c ({signal_3852, signal_2388}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2380 ( .a ({signal_7824, signal_7812}), .b ({signal_3851, signal_2387}), .clk ( clk ), .r ( Fresh[876] ), .c ({signal_3853, signal_2389}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2381 ( .a ({signal_3852, signal_2388}), .b ({signal_3854, signal_25}) ) ;
    buf_clk cell_5478 ( .C ( clk ), .D ( signal_7837 ), .Q ( signal_7838 ) ) ;
    buf_clk cell_5492 ( .C ( clk ), .D ( signal_7851 ), .Q ( signal_7852 ) ) ;
    buf_clk cell_5504 ( .C ( clk ), .D ( signal_7863 ), .Q ( signal_7864 ) ) ;
    buf_clk cell_5518 ( .C ( clk ), .D ( signal_7877 ), .Q ( signal_7878 ) ) ;
    buf_clk cell_5522 ( .C ( clk ), .D ( signal_7881 ), .Q ( signal_7882 ) ) ;
    buf_clk cell_5528 ( .C ( clk ), .D ( signal_7887 ), .Q ( signal_7888 ) ) ;
    buf_clk cell_5534 ( .C ( clk ), .D ( signal_7893 ), .Q ( signal_7894 ) ) ;
    buf_clk cell_5540 ( .C ( clk ), .D ( signal_7899 ), .Q ( signal_7900 ) ) ;
    buf_clk cell_5556 ( .C ( clk ), .D ( signal_7915 ), .Q ( signal_7916 ) ) ;
    buf_clk cell_5564 ( .C ( clk ), .D ( signal_7923 ), .Q ( signal_7924 ) ) ;
    buf_clk cell_5572 ( .C ( clk ), .D ( signal_7931 ), .Q ( signal_7932 ) ) ;
    buf_clk cell_5580 ( .C ( clk ), .D ( signal_7939 ), .Q ( signal_7940 ) ) ;
    buf_clk cell_5588 ( .C ( clk ), .D ( signal_7947 ), .Q ( signal_7948 ) ) ;
    buf_clk cell_5596 ( .C ( clk ), .D ( signal_7955 ), .Q ( signal_7956 ) ) ;
    buf_clk cell_5602 ( .C ( clk ), .D ( signal_7961 ), .Q ( signal_7962 ) ) ;
    buf_clk cell_5608 ( .C ( clk ), .D ( signal_7967 ), .Q ( signal_7968 ) ) ;

    /* cells in depth 31 */
    buf_clk cell_5505 ( .C ( clk ), .D ( signal_7864 ), .Q ( signal_7865 ) ) ;
    buf_clk cell_5519 ( .C ( clk ), .D ( signal_7878 ), .Q ( signal_7879 ) ) ;
    buf_clk cell_5523 ( .C ( clk ), .D ( signal_7882 ), .Q ( signal_7883 ) ) ;
    buf_clk cell_5529 ( .C ( clk ), .D ( signal_7888 ), .Q ( signal_7889 ) ) ;
    buf_clk cell_5535 ( .C ( clk ), .D ( signal_7894 ), .Q ( signal_7895 ) ) ;
    buf_clk cell_5541 ( .C ( clk ), .D ( signal_7900 ), .Q ( signal_7901 ) ) ;
    buf_clk cell_5545 ( .C ( clk ), .D ( signal_25 ), .Q ( signal_7905 ) ) ;
    buf_clk cell_5549 ( .C ( clk ), .D ( signal_3854 ), .Q ( signal_7909 ) ) ;
    buf_clk cell_5557 ( .C ( clk ), .D ( signal_7916 ), .Q ( signal_7917 ) ) ;
    buf_clk cell_5565 ( .C ( clk ), .D ( signal_7924 ), .Q ( signal_7925 ) ) ;
    buf_clk cell_5573 ( .C ( clk ), .D ( signal_7932 ), .Q ( signal_7933 ) ) ;
    buf_clk cell_5581 ( .C ( clk ), .D ( signal_7940 ), .Q ( signal_7941 ) ) ;
    buf_clk cell_5589 ( .C ( clk ), .D ( signal_7948 ), .Q ( signal_7949 ) ) ;
    buf_clk cell_5597 ( .C ( clk ), .D ( signal_7956 ), .Q ( signal_7957 ) ) ;
    buf_clk cell_5603 ( .C ( clk ), .D ( signal_7962 ), .Q ( signal_7963 ) ) ;
    buf_clk cell_5609 ( .C ( clk ), .D ( signal_7968 ), .Q ( signal_7969 ) ) ;

    /* cells in depth 32 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2382 ( .a ({signal_7852, signal_7838}), .b ({signal_3853, signal_2389}), .clk ( clk ), .r ( Fresh[877] ), .c ({signal_3855, signal_2390}) ) ;
    buf_clk cell_5506 ( .C ( clk ), .D ( signal_7865 ), .Q ( signal_7866 ) ) ;
    buf_clk cell_5520 ( .C ( clk ), .D ( signal_7879 ), .Q ( signal_7880 ) ) ;
    buf_clk cell_5524 ( .C ( clk ), .D ( signal_7883 ), .Q ( signal_7884 ) ) ;
    buf_clk cell_5530 ( .C ( clk ), .D ( signal_7889 ), .Q ( signal_7890 ) ) ;
    buf_clk cell_5536 ( .C ( clk ), .D ( signal_7895 ), .Q ( signal_7896 ) ) ;
    buf_clk cell_5542 ( .C ( clk ), .D ( signal_7901 ), .Q ( signal_7902 ) ) ;
    buf_clk cell_5546 ( .C ( clk ), .D ( signal_7905 ), .Q ( signal_7906 ) ) ;
    buf_clk cell_5550 ( .C ( clk ), .D ( signal_7909 ), .Q ( signal_7910 ) ) ;
    buf_clk cell_5558 ( .C ( clk ), .D ( signal_7917 ), .Q ( signal_7918 ) ) ;
    buf_clk cell_5566 ( .C ( clk ), .D ( signal_7925 ), .Q ( signal_7926 ) ) ;
    buf_clk cell_5574 ( .C ( clk ), .D ( signal_7933 ), .Q ( signal_7934 ) ) ;
    buf_clk cell_5582 ( .C ( clk ), .D ( signal_7941 ), .Q ( signal_7942 ) ) ;
    buf_clk cell_5590 ( .C ( clk ), .D ( signal_7949 ), .Q ( signal_7950 ) ) ;
    buf_clk cell_5598 ( .C ( clk ), .D ( signal_7957 ), .Q ( signal_7958 ) ) ;
    buf_clk cell_5604 ( .C ( clk ), .D ( signal_7963 ), .Q ( signal_7964 ) ) ;
    buf_clk cell_5610 ( .C ( clk ), .D ( signal_7969 ), .Q ( signal_7970 ) ) ;

    /* cells in depth 33 */
    buf_clk cell_5525 ( .C ( clk ), .D ( signal_7884 ), .Q ( signal_7885 ) ) ;
    buf_clk cell_5531 ( .C ( clk ), .D ( signal_7890 ), .Q ( signal_7891 ) ) ;
    buf_clk cell_5537 ( .C ( clk ), .D ( signal_7896 ), .Q ( signal_7897 ) ) ;
    buf_clk cell_5543 ( .C ( clk ), .D ( signal_7902 ), .Q ( signal_7903 ) ) ;
    buf_clk cell_5547 ( .C ( clk ), .D ( signal_7906 ), .Q ( signal_7907 ) ) ;
    buf_clk cell_5551 ( .C ( clk ), .D ( signal_7910 ), .Q ( signal_7911 ) ) ;
    buf_clk cell_5559 ( .C ( clk ), .D ( signal_7918 ), .Q ( signal_7919 ) ) ;
    buf_clk cell_5567 ( .C ( clk ), .D ( signal_7926 ), .Q ( signal_7927 ) ) ;
    buf_clk cell_5575 ( .C ( clk ), .D ( signal_7934 ), .Q ( signal_7935 ) ) ;
    buf_clk cell_5583 ( .C ( clk ), .D ( signal_7942 ), .Q ( signal_7943 ) ) ;
    buf_clk cell_5591 ( .C ( clk ), .D ( signal_7950 ), .Q ( signal_7951 ) ) ;
    buf_clk cell_5599 ( .C ( clk ), .D ( signal_7958 ), .Q ( signal_7959 ) ) ;
    buf_clk cell_5605 ( .C ( clk ), .D ( signal_7964 ), .Q ( signal_7965 ) ) ;
    buf_clk cell_5611 ( .C ( clk ), .D ( signal_7970 ), .Q ( signal_7971 ) ) ;

    /* cells in depth 34 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_2383 ( .a ({signal_7880, signal_7866}), .b ({signal_3855, signal_2390}), .clk ( clk ), .r ( Fresh[878] ), .c ({signal_3856, signal_2391}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_2384 ( .a ({signal_3856, signal_2391}), .b ({signal_3857, signal_27}) ) ;
    buf_clk cell_5526 ( .C ( clk ), .D ( signal_7885 ), .Q ( signal_7886 ) ) ;
    buf_clk cell_5532 ( .C ( clk ), .D ( signal_7891 ), .Q ( signal_7892 ) ) ;
    buf_clk cell_5538 ( .C ( clk ), .D ( signal_7897 ), .Q ( signal_7898 ) ) ;
    buf_clk cell_5544 ( .C ( clk ), .D ( signal_7903 ), .Q ( signal_7904 ) ) ;
    buf_clk cell_5548 ( .C ( clk ), .D ( signal_7907 ), .Q ( signal_7908 ) ) ;
    buf_clk cell_5552 ( .C ( clk ), .D ( signal_7911 ), .Q ( signal_7912 ) ) ;
    buf_clk cell_5560 ( .C ( clk ), .D ( signal_7919 ), .Q ( signal_7920 ) ) ;
    buf_clk cell_5568 ( .C ( clk ), .D ( signal_7927 ), .Q ( signal_7928 ) ) ;
    buf_clk cell_5576 ( .C ( clk ), .D ( signal_7935 ), .Q ( signal_7936 ) ) ;
    buf_clk cell_5584 ( .C ( clk ), .D ( signal_7943 ), .Q ( signal_7944 ) ) ;
    buf_clk cell_5592 ( .C ( clk ), .D ( signal_7951 ), .Q ( signal_7952 ) ) ;
    buf_clk cell_5600 ( .C ( clk ), .D ( signal_7959 ), .Q ( signal_7960 ) ) ;
    buf_clk cell_5606 ( .C ( clk ), .D ( signal_7965 ), .Q ( signal_7966 ) ) ;
    buf_clk cell_5612 ( .C ( clk ), .D ( signal_7971 ), .Q ( signal_7972 ) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_7892, signal_7886}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_7904, signal_7898}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_7912, signal_7908}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_7928, signal_7920}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_4 ( .clk ( clk ), .D ({signal_3857, signal_27}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_5 ( .clk ( clk ), .D ({signal_7944, signal_7936}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_6 ( .clk ( clk ), .D ({signal_7960, signal_7952}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_7 ( .clk ( clk ), .D ({signal_7972, signal_7966}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
