/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 12 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 13 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d1 (SI_s0, clk, SI_s1, Fresh, SO_s0, SO_s1);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [16:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    wire signal_15 ;
    wire signal_16 ;
    wire signal_17 ;
    wire signal_18 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_57 ;
    wire signal_58 ;
    wire signal_59 ;
    wire signal_60 ;
    wire signal_61 ;
    wire signal_62 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_66 ;
    wire signal_68 ;
    wire signal_70 ;
    wire signal_72 ;
    wire signal_73 ;
    wire signal_74 ;
    wire signal_75 ;
    wire signal_76 ;
    wire signal_77 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_83 ;
    wire signal_84 ;
    wire signal_85 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_141 ;
    wire signal_142 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(1)) cell_23 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_66, signal_34}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_24 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_68, signal_35}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_25 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_70, signal_36}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_26 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_72, signal_37}) ) ;

    /* cells in depth 1 */
    buf_clk cell_58 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( signal_125 ) ) ;
    buf_clk cell_60 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( signal_127 ) ) ;
    buf_clk cell_62 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( signal_129 ) ) ;
    buf_clk cell_64 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( signal_131 ) ) ;
    buf_clk cell_66 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( signal_133 ) ) ;
    buf_clk cell_68 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( signal_135 ) ) ;
    buf_clk cell_70 ( .C ( clk ), .D ( signal_34 ), .Q ( signal_137 ) ) ;
    buf_clk cell_72 ( .C ( clk ), .D ( signal_66 ), .Q ( signal_139 ) ) ;
    buf_clk cell_74 ( .C ( clk ), .D ( signal_36 ), .Q ( signal_141 ) ) ;
    buf_clk cell_76 ( .C ( clk ), .D ( signal_70 ), .Q ( signal_143 ) ) ;
    buf_clk cell_90 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( signal_157 ) ) ;
    buf_clk cell_96 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( signal_163 ) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_27 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_73, signal_38}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_28 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_74, signal_39}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_29 ( .a ({signal_73, signal_38}), .b ({signal_75, signal_40}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_30 ( .a ({signal_74, signal_39}), .b ({signal_76, signal_41}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_31 ( .a ({signal_68, signal_35}), .b ({signal_70, signal_36}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_77, signal_42}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_32 ( .a ({signal_66, signal_34}), .b ({signal_72, signal_37}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_78, signal_43}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_33 ( .a ({signal_68, signal_35}), .b ({signal_72, signal_37}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_79, signal_44}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_34 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_68, signal_35}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_80, signal_45}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_35 ( .a ({signal_66, signal_34}), .b ({signal_68, signal_35}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_81, signal_46}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_36 ( .a ({signal_79, signal_44}), .b ({signal_82, signal_47}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_39 ( .a ({signal_128, signal_126}), .b ({signal_77, signal_42}), .c ({signal_85, signal_16}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_40 ( .a ({signal_132, signal_130}), .b ({signal_80, signal_45}), .c ({signal_86, signal_50}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_41 ( .a ({signal_132, signal_130}), .b ({signal_81, signal_46}), .c ({signal_87, signal_15}) ) ;
    buf_clk cell_59 ( .C ( clk ), .D ( signal_125 ), .Q ( signal_126 ) ) ;
    buf_clk cell_61 ( .C ( clk ), .D ( signal_127 ), .Q ( signal_128 ) ) ;
    buf_clk cell_63 ( .C ( clk ), .D ( signal_129 ), .Q ( signal_130 ) ) ;
    buf_clk cell_65 ( .C ( clk ), .D ( signal_131 ), .Q ( signal_132 ) ) ;
    buf_clk cell_67 ( .C ( clk ), .D ( signal_133 ), .Q ( signal_134 ) ) ;
    buf_clk cell_69 ( .C ( clk ), .D ( signal_135 ), .Q ( signal_136 ) ) ;
    buf_clk cell_71 ( .C ( clk ), .D ( signal_137 ), .Q ( signal_138 ) ) ;
    buf_clk cell_73 ( .C ( clk ), .D ( signal_139 ), .Q ( signal_140 ) ) ;
    buf_clk cell_75 ( .C ( clk ), .D ( signal_141 ), .Q ( signal_142 ) ) ;
    buf_clk cell_77 ( .C ( clk ), .D ( signal_143 ), .Q ( signal_144 ) ) ;
    buf_clk cell_91 ( .C ( clk ), .D ( signal_157 ), .Q ( signal_158 ) ) ;
    buf_clk cell_97 ( .C ( clk ), .D ( signal_163 ), .Q ( signal_164 ) ) ;

    /* cells in depth 3 */
    buf_clk cell_78 ( .C ( clk ), .D ( signal_40 ), .Q ( signal_145 ) ) ;
    buf_clk cell_80 ( .C ( clk ), .D ( signal_75 ), .Q ( signal_147 ) ) ;
    buf_clk cell_82 ( .C ( clk ), .D ( signal_142 ), .Q ( signal_149 ) ) ;
    buf_clk cell_84 ( .C ( clk ), .D ( signal_144 ), .Q ( signal_151 ) ) ;
    buf_clk cell_86 ( .C ( clk ), .D ( signal_41 ), .Q ( signal_153 ) ) ;
    buf_clk cell_88 ( .C ( clk ), .D ( signal_76 ), .Q ( signal_155 ) ) ;
    buf_clk cell_92 ( .C ( clk ), .D ( signal_158 ), .Q ( signal_159 ) ) ;
    buf_clk cell_98 ( .C ( clk ), .D ( signal_164 ), .Q ( signal_165 ) ) ;
    buf_clk cell_118 ( .C ( clk ), .D ( signal_15 ), .Q ( signal_185 ) ) ;
    buf_clk cell_128 ( .C ( clk ), .D ( signal_87 ), .Q ( signal_195 ) ) ;
    buf_clk cell_138 ( .C ( clk ), .D ( signal_16 ), .Q ( signal_205 ) ) ;
    buf_clk cell_148 ( .C ( clk ), .D ( signal_85 ), .Q ( signal_215 ) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_37 ( .a ({signal_136, signal_134}), .b ({signal_78, signal_43}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_83, signal_48}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_38 ( .a ({signal_128, signal_126}), .b ({signal_79, signal_44}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_84, signal_49}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_42 ( .a ({signal_83, signal_48}), .b ({signal_88, signal_51}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_43 ( .a ({signal_84, signal_49}), .b ({signal_89, signal_52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_44 ( .a ({signal_140, signal_138}), .b ({signal_82, signal_47}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_90, signal_53}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_45 ( .a ({signal_144, signal_142}), .b ({signal_86, signal_50}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_91, signal_54}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_46 ( .a ({signal_91, signal_54}), .b ({signal_92, signal_55}) ) ;
    buf_clk cell_79 ( .C ( clk ), .D ( signal_145 ), .Q ( signal_146 ) ) ;
    buf_clk cell_81 ( .C ( clk ), .D ( signal_147 ), .Q ( signal_148 ) ) ;
    buf_clk cell_83 ( .C ( clk ), .D ( signal_149 ), .Q ( signal_150 ) ) ;
    buf_clk cell_85 ( .C ( clk ), .D ( signal_151 ), .Q ( signal_152 ) ) ;
    buf_clk cell_87 ( .C ( clk ), .D ( signal_153 ), .Q ( signal_154 ) ) ;
    buf_clk cell_89 ( .C ( clk ), .D ( signal_155 ), .Q ( signal_156 ) ) ;
    buf_clk cell_93 ( .C ( clk ), .D ( signal_159 ), .Q ( signal_160 ) ) ;
    buf_clk cell_99 ( .C ( clk ), .D ( signal_165 ), .Q ( signal_166 ) ) ;
    buf_clk cell_119 ( .C ( clk ), .D ( signal_185 ), .Q ( signal_186 ) ) ;
    buf_clk cell_129 ( .C ( clk ), .D ( signal_195 ), .Q ( signal_196 ) ) ;
    buf_clk cell_139 ( .C ( clk ), .D ( signal_205 ), .Q ( signal_206 ) ) ;
    buf_clk cell_149 ( .C ( clk ), .D ( signal_215 ), .Q ( signal_216 ) ) ;

    /* cells in depth 5 */
    buf_clk cell_94 ( .C ( clk ), .D ( signal_160 ), .Q ( signal_161 ) ) ;
    buf_clk cell_100 ( .C ( clk ), .D ( signal_166 ), .Q ( signal_167 ) ) ;
    buf_clk cell_106 ( .C ( clk ), .D ( signal_52 ), .Q ( signal_173 ) ) ;
    buf_clk cell_112 ( .C ( clk ), .D ( signal_89 ), .Q ( signal_179 ) ) ;
    buf_clk cell_120 ( .C ( clk ), .D ( signal_186 ), .Q ( signal_187 ) ) ;
    buf_clk cell_130 ( .C ( clk ), .D ( signal_196 ), .Q ( signal_197 ) ) ;
    buf_clk cell_140 ( .C ( clk ), .D ( signal_206 ), .Q ( signal_207 ) ) ;
    buf_clk cell_150 ( .C ( clk ), .D ( signal_216 ), .Q ( signal_217 ) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_47 ( .a ({signal_148, signal_146}), .b ({signal_90, signal_53}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_93, signal_56}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_48 ( .a ({signal_152, signal_150}), .b ({signal_88, signal_51}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_94, signal_57}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_49 ( .a ({signal_94, signal_57}), .b ({signal_95, signal_58}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_50 ( .a ({signal_92, signal_55}), .b ({signal_156, signal_154}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_96, signal_59}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_52 ( .a ({signal_96, signal_59}), .b ({signal_98, signal_17}) ) ;
    buf_clk cell_95 ( .C ( clk ), .D ( signal_161 ), .Q ( signal_162 ) ) ;
    buf_clk cell_101 ( .C ( clk ), .D ( signal_167 ), .Q ( signal_168 ) ) ;
    buf_clk cell_107 ( .C ( clk ), .D ( signal_173 ), .Q ( signal_174 ) ) ;
    buf_clk cell_113 ( .C ( clk ), .D ( signal_179 ), .Q ( signal_180 ) ) ;
    buf_clk cell_121 ( .C ( clk ), .D ( signal_187 ), .Q ( signal_188 ) ) ;
    buf_clk cell_131 ( .C ( clk ), .D ( signal_197 ), .Q ( signal_198 ) ) ;
    buf_clk cell_141 ( .C ( clk ), .D ( signal_207 ), .Q ( signal_208 ) ) ;
    buf_clk cell_151 ( .C ( clk ), .D ( signal_217 ), .Q ( signal_218 ) ) ;

    /* cells in depth 7 */
    buf_clk cell_102 ( .C ( clk ), .D ( signal_58 ), .Q ( signal_169 ) ) ;
    buf_clk cell_104 ( .C ( clk ), .D ( signal_95 ), .Q ( signal_171 ) ) ;
    buf_clk cell_108 ( .C ( clk ), .D ( signal_174 ), .Q ( signal_175 ) ) ;
    buf_clk cell_114 ( .C ( clk ), .D ( signal_180 ), .Q ( signal_181 ) ) ;
    buf_clk cell_122 ( .C ( clk ), .D ( signal_188 ), .Q ( signal_189 ) ) ;
    buf_clk cell_132 ( .C ( clk ), .D ( signal_198 ), .Q ( signal_199 ) ) ;
    buf_clk cell_142 ( .C ( clk ), .D ( signal_208 ), .Q ( signal_209 ) ) ;
    buf_clk cell_152 ( .C ( clk ), .D ( signal_218 ), .Q ( signal_219 ) ) ;
    buf_clk cell_158 ( .C ( clk ), .D ( signal_17 ), .Q ( signal_225 ) ) ;
    buf_clk cell_164 ( .C ( clk ), .D ( signal_98 ), .Q ( signal_231 ) ) ;

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_51 ( .a ({signal_168, signal_162}), .b ({signal_93, signal_56}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_97, signal_60}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_53 ( .a ({signal_97, signal_60}), .b ({signal_99, signal_61}) ) ;
    buf_clk cell_103 ( .C ( clk ), .D ( signal_169 ), .Q ( signal_170 ) ) ;
    buf_clk cell_105 ( .C ( clk ), .D ( signal_171 ), .Q ( signal_172 ) ) ;
    buf_clk cell_109 ( .C ( clk ), .D ( signal_175 ), .Q ( signal_176 ) ) ;
    buf_clk cell_115 ( .C ( clk ), .D ( signal_181 ), .Q ( signal_182 ) ) ;
    buf_clk cell_123 ( .C ( clk ), .D ( signal_189 ), .Q ( signal_190 ) ) ;
    buf_clk cell_133 ( .C ( clk ), .D ( signal_199 ), .Q ( signal_200 ) ) ;
    buf_clk cell_143 ( .C ( clk ), .D ( signal_209 ), .Q ( signal_210 ) ) ;
    buf_clk cell_153 ( .C ( clk ), .D ( signal_219 ), .Q ( signal_220 ) ) ;
    buf_clk cell_159 ( .C ( clk ), .D ( signal_225 ), .Q ( signal_226 ) ) ;
    buf_clk cell_165 ( .C ( clk ), .D ( signal_231 ), .Q ( signal_232 ) ) ;

    /* cells in depth 9 */
    buf_clk cell_110 ( .C ( clk ), .D ( signal_176 ), .Q ( signal_177 ) ) ;
    buf_clk cell_116 ( .C ( clk ), .D ( signal_182 ), .Q ( signal_183 ) ) ;
    buf_clk cell_124 ( .C ( clk ), .D ( signal_190 ), .Q ( signal_191 ) ) ;
    buf_clk cell_134 ( .C ( clk ), .D ( signal_200 ), .Q ( signal_201 ) ) ;
    buf_clk cell_144 ( .C ( clk ), .D ( signal_210 ), .Q ( signal_211 ) ) ;
    buf_clk cell_154 ( .C ( clk ), .D ( signal_220 ), .Q ( signal_221 ) ) ;
    buf_clk cell_160 ( .C ( clk ), .D ( signal_226 ), .Q ( signal_227 ) ) ;
    buf_clk cell_166 ( .C ( clk ), .D ( signal_232 ), .Q ( signal_233 ) ) ;

    /* cells in depth 10 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_54 ( .a ({signal_172, signal_170}), .b ({signal_99, signal_61}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_100, signal_62}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_55 ( .a ({signal_100, signal_62}), .b ({signal_101, signal_63}) ) ;
    buf_clk cell_111 ( .C ( clk ), .D ( signal_177 ), .Q ( signal_178 ) ) ;
    buf_clk cell_117 ( .C ( clk ), .D ( signal_183 ), .Q ( signal_184 ) ) ;
    buf_clk cell_125 ( .C ( clk ), .D ( signal_191 ), .Q ( signal_192 ) ) ;
    buf_clk cell_135 ( .C ( clk ), .D ( signal_201 ), .Q ( signal_202 ) ) ;
    buf_clk cell_145 ( .C ( clk ), .D ( signal_211 ), .Q ( signal_212 ) ) ;
    buf_clk cell_155 ( .C ( clk ), .D ( signal_221 ), .Q ( signal_222 ) ) ;
    buf_clk cell_161 ( .C ( clk ), .D ( signal_227 ), .Q ( signal_228 ) ) ;
    buf_clk cell_167 ( .C ( clk ), .D ( signal_233 ), .Q ( signal_234 ) ) ;

    /* cells in depth 11 */
    buf_clk cell_126 ( .C ( clk ), .D ( signal_192 ), .Q ( signal_193 ) ) ;
    buf_clk cell_136 ( .C ( clk ), .D ( signal_202 ), .Q ( signal_203 ) ) ;
    buf_clk cell_146 ( .C ( clk ), .D ( signal_212 ), .Q ( signal_213 ) ) ;
    buf_clk cell_156 ( .C ( clk ), .D ( signal_222 ), .Q ( signal_223 ) ) ;
    buf_clk cell_162 ( .C ( clk ), .D ( signal_228 ), .Q ( signal_229 ) ) ;
    buf_clk cell_168 ( .C ( clk ), .D ( signal_234 ), .Q ( signal_235 ) ) ;

    /* cells in depth 12 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_56 ( .a ({signal_184, signal_178}), .b ({signal_101, signal_63}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_102, signal_64}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_57 ( .a ({signal_102, signal_64}), .b ({signal_103, signal_18}) ) ;
    buf_clk cell_127 ( .C ( clk ), .D ( signal_193 ), .Q ( signal_194 ) ) ;
    buf_clk cell_137 ( .C ( clk ), .D ( signal_203 ), .Q ( signal_204 ) ) ;
    buf_clk cell_147 ( .C ( clk ), .D ( signal_213 ), .Q ( signal_214 ) ) ;
    buf_clk cell_157 ( .C ( clk ), .D ( signal_223 ), .Q ( signal_224 ) ) ;
    buf_clk cell_163 ( .C ( clk ), .D ( signal_229 ), .Q ( signal_230 ) ) ;
    buf_clk cell_169 ( .C ( clk ), .D ( signal_235 ), .Q ( signal_236 ) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk ( clk ), .D ({signal_204, signal_194}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk ( clk ), .D ({signal_224, signal_214}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk ( clk ), .D ({signal_236, signal_230}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk ( clk ), .D ({signal_103, signal_18}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
