/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* 34 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 35 register stage(s) in total */

module sbox_HPC2_Pipeline_d3 (SI_s0, clk, SI_s1, SI_s2, SI_s3, Fresh, SO_s0, SO_s1, SO_s2, SO_s3);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input [7:0] SI_s2 ;
    input [7:0] SI_s3 ;
    input [5207:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output [7:0] SO_s2 ;
    output [7:0] SO_s3 ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_946 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_952 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13393 ;
    wire new_AGEMA_signal_13394 ;
    wire new_AGEMA_signal_13395 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13399 ;
    wire new_AGEMA_signal_13400 ;
    wire new_AGEMA_signal_13401 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13405 ;
    wire new_AGEMA_signal_13406 ;
    wire new_AGEMA_signal_13407 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13891 ;
    wire new_AGEMA_signal_13892 ;
    wire new_AGEMA_signal_13893 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13897 ;
    wire new_AGEMA_signal_13898 ;
    wire new_AGEMA_signal_13899 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13903 ;
    wire new_AGEMA_signal_13904 ;
    wire new_AGEMA_signal_13905 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13909 ;
    wire new_AGEMA_signal_13910 ;
    wire new_AGEMA_signal_13911 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13915 ;
    wire new_AGEMA_signal_13916 ;
    wire new_AGEMA_signal_13917 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13921 ;
    wire new_AGEMA_signal_13922 ;
    wire new_AGEMA_signal_13923 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13927 ;
    wire new_AGEMA_signal_13928 ;
    wire new_AGEMA_signal_13929 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13933 ;
    wire new_AGEMA_signal_13934 ;
    wire new_AGEMA_signal_13935 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13939 ;
    wire new_AGEMA_signal_13940 ;
    wire new_AGEMA_signal_13941 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13945 ;
    wire new_AGEMA_signal_13946 ;
    wire new_AGEMA_signal_13947 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13951 ;
    wire new_AGEMA_signal_13952 ;
    wire new_AGEMA_signal_13953 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13957 ;
    wire new_AGEMA_signal_13958 ;
    wire new_AGEMA_signal_13959 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13963 ;
    wire new_AGEMA_signal_13964 ;
    wire new_AGEMA_signal_13965 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13969 ;
    wire new_AGEMA_signal_13970 ;
    wire new_AGEMA_signal_13971 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13975 ;
    wire new_AGEMA_signal_13976 ;
    wire new_AGEMA_signal_13977 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13981 ;
    wire new_AGEMA_signal_13982 ;
    wire new_AGEMA_signal_13983 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13987 ;
    wire new_AGEMA_signal_13988 ;
    wire new_AGEMA_signal_13989 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13993 ;
    wire new_AGEMA_signal_13994 ;
    wire new_AGEMA_signal_13995 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_13999 ;
    wire new_AGEMA_signal_14000 ;
    wire new_AGEMA_signal_14001 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14005 ;
    wire new_AGEMA_signal_14006 ;
    wire new_AGEMA_signal_14007 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14011 ;
    wire new_AGEMA_signal_14012 ;
    wire new_AGEMA_signal_14013 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14017 ;
    wire new_AGEMA_signal_14018 ;
    wire new_AGEMA_signal_14019 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14023 ;
    wire new_AGEMA_signal_14024 ;
    wire new_AGEMA_signal_14025 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14029 ;
    wire new_AGEMA_signal_14030 ;
    wire new_AGEMA_signal_14031 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14035 ;
    wire new_AGEMA_signal_14036 ;
    wire new_AGEMA_signal_14037 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14521 ;
    wire new_AGEMA_signal_14522 ;
    wire new_AGEMA_signal_14523 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14527 ;
    wire new_AGEMA_signal_14528 ;
    wire new_AGEMA_signal_14529 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14533 ;
    wire new_AGEMA_signal_14534 ;
    wire new_AGEMA_signal_14535 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14539 ;
    wire new_AGEMA_signal_14540 ;
    wire new_AGEMA_signal_14541 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14545 ;
    wire new_AGEMA_signal_14546 ;
    wire new_AGEMA_signal_14547 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14551 ;
    wire new_AGEMA_signal_14552 ;
    wire new_AGEMA_signal_14553 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14557 ;
    wire new_AGEMA_signal_14558 ;
    wire new_AGEMA_signal_14559 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14563 ;
    wire new_AGEMA_signal_14564 ;
    wire new_AGEMA_signal_14565 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14569 ;
    wire new_AGEMA_signal_14570 ;
    wire new_AGEMA_signal_14571 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14575 ;
    wire new_AGEMA_signal_14576 ;
    wire new_AGEMA_signal_14577 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14581 ;
    wire new_AGEMA_signal_14582 ;
    wire new_AGEMA_signal_14583 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14587 ;
    wire new_AGEMA_signal_14588 ;
    wire new_AGEMA_signal_14589 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14593 ;
    wire new_AGEMA_signal_14594 ;
    wire new_AGEMA_signal_14595 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14599 ;
    wire new_AGEMA_signal_14600 ;
    wire new_AGEMA_signal_14601 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14605 ;
    wire new_AGEMA_signal_14606 ;
    wire new_AGEMA_signal_14607 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14611 ;
    wire new_AGEMA_signal_14612 ;
    wire new_AGEMA_signal_14613 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14617 ;
    wire new_AGEMA_signal_14618 ;
    wire new_AGEMA_signal_14619 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14623 ;
    wire new_AGEMA_signal_14624 ;
    wire new_AGEMA_signal_14625 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14629 ;
    wire new_AGEMA_signal_14630 ;
    wire new_AGEMA_signal_14631 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14635 ;
    wire new_AGEMA_signal_14636 ;
    wire new_AGEMA_signal_14637 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14641 ;
    wire new_AGEMA_signal_14642 ;
    wire new_AGEMA_signal_14643 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14647 ;
    wire new_AGEMA_signal_14648 ;
    wire new_AGEMA_signal_14649 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14653 ;
    wire new_AGEMA_signal_14654 ;
    wire new_AGEMA_signal_14655 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14659 ;
    wire new_AGEMA_signal_14660 ;
    wire new_AGEMA_signal_14661 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14665 ;
    wire new_AGEMA_signal_14666 ;
    wire new_AGEMA_signal_14667 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14671 ;
    wire new_AGEMA_signal_14672 ;
    wire new_AGEMA_signal_14673 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14677 ;
    wire new_AGEMA_signal_14678 ;
    wire new_AGEMA_signal_14679 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14683 ;
    wire new_AGEMA_signal_14684 ;
    wire new_AGEMA_signal_14685 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14689 ;
    wire new_AGEMA_signal_14690 ;
    wire new_AGEMA_signal_14691 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14695 ;
    wire new_AGEMA_signal_14696 ;
    wire new_AGEMA_signal_14697 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14701 ;
    wire new_AGEMA_signal_14702 ;
    wire new_AGEMA_signal_14703 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14707 ;
    wire new_AGEMA_signal_14708 ;
    wire new_AGEMA_signal_14709 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15193 ;
    wire new_AGEMA_signal_15194 ;
    wire new_AGEMA_signal_15195 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15199 ;
    wire new_AGEMA_signal_15200 ;
    wire new_AGEMA_signal_15201 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15205 ;
    wire new_AGEMA_signal_15206 ;
    wire new_AGEMA_signal_15207 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15211 ;
    wire new_AGEMA_signal_15212 ;
    wire new_AGEMA_signal_15213 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15217 ;
    wire new_AGEMA_signal_15218 ;
    wire new_AGEMA_signal_15219 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15223 ;
    wire new_AGEMA_signal_15224 ;
    wire new_AGEMA_signal_15225 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15229 ;
    wire new_AGEMA_signal_15230 ;
    wire new_AGEMA_signal_15231 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15235 ;
    wire new_AGEMA_signal_15236 ;
    wire new_AGEMA_signal_15237 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15241 ;
    wire new_AGEMA_signal_15242 ;
    wire new_AGEMA_signal_15243 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15247 ;
    wire new_AGEMA_signal_15248 ;
    wire new_AGEMA_signal_15249 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15253 ;
    wire new_AGEMA_signal_15254 ;
    wire new_AGEMA_signal_15255 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15259 ;
    wire new_AGEMA_signal_15260 ;
    wire new_AGEMA_signal_15261 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15265 ;
    wire new_AGEMA_signal_15266 ;
    wire new_AGEMA_signal_15267 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15271 ;
    wire new_AGEMA_signal_15272 ;
    wire new_AGEMA_signal_15273 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15277 ;
    wire new_AGEMA_signal_15278 ;
    wire new_AGEMA_signal_15279 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15283 ;
    wire new_AGEMA_signal_15284 ;
    wire new_AGEMA_signal_15285 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15289 ;
    wire new_AGEMA_signal_15290 ;
    wire new_AGEMA_signal_15291 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15295 ;
    wire new_AGEMA_signal_15296 ;
    wire new_AGEMA_signal_15297 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15301 ;
    wire new_AGEMA_signal_15302 ;
    wire new_AGEMA_signal_15303 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15307 ;
    wire new_AGEMA_signal_15308 ;
    wire new_AGEMA_signal_15309 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15313 ;
    wire new_AGEMA_signal_15314 ;
    wire new_AGEMA_signal_15315 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15319 ;
    wire new_AGEMA_signal_15320 ;
    wire new_AGEMA_signal_15321 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15325 ;
    wire new_AGEMA_signal_15326 ;
    wire new_AGEMA_signal_15327 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15331 ;
    wire new_AGEMA_signal_15332 ;
    wire new_AGEMA_signal_15333 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15337 ;
    wire new_AGEMA_signal_15338 ;
    wire new_AGEMA_signal_15339 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15343 ;
    wire new_AGEMA_signal_15344 ;
    wire new_AGEMA_signal_15345 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15349 ;
    wire new_AGEMA_signal_15350 ;
    wire new_AGEMA_signal_15351 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15355 ;
    wire new_AGEMA_signal_15356 ;
    wire new_AGEMA_signal_15357 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15361 ;
    wire new_AGEMA_signal_15362 ;
    wire new_AGEMA_signal_15363 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15367 ;
    wire new_AGEMA_signal_15368 ;
    wire new_AGEMA_signal_15369 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15373 ;
    wire new_AGEMA_signal_15374 ;
    wire new_AGEMA_signal_15375 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15379 ;
    wire new_AGEMA_signal_15380 ;
    wire new_AGEMA_signal_15381 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(1)) U1938 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1939 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1940 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1941 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1942 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1944 ( .a ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1945 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1946 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_927 ( .C ( clk ), .D ( SI_s0[4] ), .Q ( new_AGEMA_signal_8955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C ( clk ), .D ( SI_s1[4] ), .Q ( new_AGEMA_signal_8957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C ( clk ), .D ( SI_s2[4] ), .Q ( new_AGEMA_signal_8959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C ( clk ), .D ( SI_s3[4] ), .Q ( new_AGEMA_signal_8961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C ( clk ), .D ( SI_s0[6] ), .Q ( new_AGEMA_signal_8963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C ( clk ), .D ( SI_s1[6] ), .Q ( new_AGEMA_signal_8965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C ( clk ), .D ( SI_s2[6] ), .Q ( new_AGEMA_signal_8967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C ( clk ), .D ( SI_s3[6] ), .Q ( new_AGEMA_signal_8969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C ( clk ), .D ( SI_s0[7] ), .Q ( new_AGEMA_signal_8971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C ( clk ), .D ( SI_s1[7] ), .Q ( new_AGEMA_signal_8973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C ( clk ), .D ( SI_s2[7] ), .Q ( new_AGEMA_signal_8975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C ( clk ), .D ( SI_s3[7] ), .Q ( new_AGEMA_signal_8977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C ( clk ), .D ( SI_s0[0] ), .Q ( new_AGEMA_signal_8979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C ( clk ), .D ( SI_s1[0] ), .Q ( new_AGEMA_signal_8981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C ( clk ), .D ( SI_s2[0] ), .Q ( new_AGEMA_signal_8983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C ( clk ), .D ( SI_s3[0] ), .Q ( new_AGEMA_signal_8985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_8987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_8989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_8991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( new_AGEMA_signal_8993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C ( clk ), .D ( n2630 ), .Q ( new_AGEMA_signal_8995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C ( clk ), .D ( new_AGEMA_signal_981 ), .Q ( new_AGEMA_signal_8997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C ( clk ), .D ( new_AGEMA_signal_982 ), .Q ( new_AGEMA_signal_8999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C ( clk ), .D ( new_AGEMA_signal_983 ), .Q ( new_AGEMA_signal_9001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C ( clk ), .D ( SI_s0[5] ), .Q ( new_AGEMA_signal_9003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C ( clk ), .D ( SI_s1[5] ), .Q ( new_AGEMA_signal_9005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C ( clk ), .D ( SI_s2[5] ), .Q ( new_AGEMA_signal_9007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C ( clk ), .D ( SI_s3[5] ), .Q ( new_AGEMA_signal_9009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C ( clk ), .D ( n2462 ), .Q ( new_AGEMA_signal_9011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C ( clk ), .D ( new_AGEMA_signal_957 ), .Q ( new_AGEMA_signal_9013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C ( clk ), .D ( new_AGEMA_signal_958 ), .Q ( new_AGEMA_signal_9015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C ( clk ), .D ( new_AGEMA_signal_959 ), .Q ( new_AGEMA_signal_9017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C ( clk ), .D ( n2760 ), .Q ( new_AGEMA_signal_9019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C ( clk ), .D ( new_AGEMA_signal_963 ), .Q ( new_AGEMA_signal_9021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C ( clk ), .D ( new_AGEMA_signal_964 ), .Q ( new_AGEMA_signal_9023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C ( clk ), .D ( new_AGEMA_signal_965 ), .Q ( new_AGEMA_signal_9025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C ( clk ), .D ( n2796 ), .Q ( new_AGEMA_signal_9027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C ( clk ), .D ( new_AGEMA_signal_945 ), .Q ( new_AGEMA_signal_9029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C ( clk ), .D ( new_AGEMA_signal_946 ), .Q ( new_AGEMA_signal_9031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C ( clk ), .D ( new_AGEMA_signal_947 ), .Q ( new_AGEMA_signal_9033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C ( clk ), .D ( n2765 ), .Q ( new_AGEMA_signal_9035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C ( clk ), .D ( new_AGEMA_signal_987 ), .Q ( new_AGEMA_signal_9037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C ( clk ), .D ( new_AGEMA_signal_988 ), .Q ( new_AGEMA_signal_9039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C ( clk ), .D ( new_AGEMA_signal_989 ), .Q ( new_AGEMA_signal_9041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C ( clk ), .D ( n2791 ), .Q ( new_AGEMA_signal_9043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C ( clk ), .D ( new_AGEMA_signal_969 ), .Q ( new_AGEMA_signal_9045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C ( clk ), .D ( new_AGEMA_signal_970 ), .Q ( new_AGEMA_signal_9047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C ( clk ), .D ( new_AGEMA_signal_971 ), .Q ( new_AGEMA_signal_9049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_9051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_9053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_9055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( new_AGEMA_signal_9057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C ( clk ), .D ( n2813 ), .Q ( new_AGEMA_signal_9059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C ( clk ), .D ( new_AGEMA_signal_975 ), .Q ( new_AGEMA_signal_9061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C ( clk ), .D ( new_AGEMA_signal_976 ), .Q ( new_AGEMA_signal_9063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C ( clk ), .D ( new_AGEMA_signal_977 ), .Q ( new_AGEMA_signal_9065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C ( clk ), .D ( n2810 ), .Q ( new_AGEMA_signal_9067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C ( clk ), .D ( new_AGEMA_signal_951 ), .Q ( new_AGEMA_signal_9069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C ( clk ), .D ( new_AGEMA_signal_952 ), .Q ( new_AGEMA_signal_9071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C ( clk ), .D ( new_AGEMA_signal_953 ), .Q ( new_AGEMA_signal_9073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_10099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_10105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_10111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( new_AGEMA_signal_10117 ) ) ;

    /* cells in depth 2 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1937 ( .a ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .b ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1943 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1947 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1948 ( .a ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .b ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1949 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1950 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1951 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1952 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1953 ( .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1955 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1956 ( .a ({new_AGEMA_signal_1040, new_AGEMA_signal_1039, new_AGEMA_signal_1038, n2699}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1957 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1958 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1961 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1962 ( .a ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1963 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1965 ( .a ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1966 ( .a ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1969 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1970 ( .a ({new_AGEMA_signal_1055, new_AGEMA_signal_1054, new_AGEMA_signal_1053, n2073}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1971 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1972 ( .a ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1973 ( .a ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1975 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1976 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1978 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .b ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1979 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1984 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1985 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1987 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1990 ( .a ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1991 ( .a ({new_AGEMA_signal_1073, new_AGEMA_signal_1072, new_AGEMA_signal_1071, n2538}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1995 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1996 ( .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1999 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2000 ( .a ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .b ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2004 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2008 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2009 ( .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2013 ( .a ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2014 ( .a ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2017 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2018 ( .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2020 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2021 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2025 ( .a ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2028 ( .a ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .b ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2029 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2035 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2036 ( .a ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2038 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2044 ( .a ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .b ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .clk ( clk ), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2045 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2046 ( .a ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2052 ( .a ({SI_s3[7], SI_s2[7], SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2055 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2068 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2070 ( .a ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2071 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2074 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .b ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2089 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2090 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2094 ( .a ({SI_s3[6], SI_s2[6], SI_s1[6], SI_s0[6]}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2096 ( .a ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2097 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2100 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2119 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2122 ( .a ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2131 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2133 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2134 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2138 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({new_AGEMA_signal_965, new_AGEMA_signal_964, new_AGEMA_signal_963, n2760}), .clk ( clk ), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2139 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2150 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .b ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2163 ( .a ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .b ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .clk ( clk ), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2211 ( .a ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .b ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2061}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2232 ( .a ({new_AGEMA_signal_947, new_AGEMA_signal_946, new_AGEMA_signal_945, n2796}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2276 ( .a ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .b ({new_AGEMA_signal_989, new_AGEMA_signal_988, new_AGEMA_signal_987, n2765}), .clk ( clk ), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2278 ( .a ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .b ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, new_AGEMA_signal_1356, n2118}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2307 ( .a ({SI_s3[4], SI_s2[4], SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_983, new_AGEMA_signal_982, new_AGEMA_signal_981, n2630}), .clk ( clk ), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2341 ( .a ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_971, new_AGEMA_signal_970, new_AGEMA_signal_969, n2791}), .clk ( clk ), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2383 ( .a ({SI_s3[5], SI_s2[5], SI_s1[5], SI_s0[5]}), .b ({SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2402 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_977, new_AGEMA_signal_976, new_AGEMA_signal_975, n2813}), .clk ( clk ), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2615 ( .a ({SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_959, new_AGEMA_signal_958, new_AGEMA_signal_957, n2462}), .clk ( clk ), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, n2463}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2627 ( .a ({new_AGEMA_signal_953, new_AGEMA_signal_952, new_AGEMA_signal_951, n2810}), .b ({SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2474}) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C ( clk ), .D ( new_AGEMA_signal_8955 ), .Q ( new_AGEMA_signal_8956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C ( clk ), .D ( new_AGEMA_signal_8957 ), .Q ( new_AGEMA_signal_8958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C ( clk ), .D ( new_AGEMA_signal_8959 ), .Q ( new_AGEMA_signal_8960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C ( clk ), .D ( new_AGEMA_signal_8961 ), .Q ( new_AGEMA_signal_8962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C ( clk ), .D ( new_AGEMA_signal_8963 ), .Q ( new_AGEMA_signal_8964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C ( clk ), .D ( new_AGEMA_signal_8965 ), .Q ( new_AGEMA_signal_8966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C ( clk ), .D ( new_AGEMA_signal_8967 ), .Q ( new_AGEMA_signal_8968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C ( clk ), .D ( new_AGEMA_signal_8969 ), .Q ( new_AGEMA_signal_8970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C ( clk ), .D ( new_AGEMA_signal_8971 ), .Q ( new_AGEMA_signal_8972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C ( clk ), .D ( new_AGEMA_signal_8973 ), .Q ( new_AGEMA_signal_8974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C ( clk ), .D ( new_AGEMA_signal_8975 ), .Q ( new_AGEMA_signal_8976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C ( clk ), .D ( new_AGEMA_signal_8977 ), .Q ( new_AGEMA_signal_8978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C ( clk ), .D ( new_AGEMA_signal_8979 ), .Q ( new_AGEMA_signal_8980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C ( clk ), .D ( new_AGEMA_signal_8981 ), .Q ( new_AGEMA_signal_8982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C ( clk ), .D ( new_AGEMA_signal_8983 ), .Q ( new_AGEMA_signal_8984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C ( clk ), .D ( new_AGEMA_signal_8985 ), .Q ( new_AGEMA_signal_8986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C ( clk ), .D ( new_AGEMA_signal_8987 ), .Q ( new_AGEMA_signal_8988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C ( clk ), .D ( new_AGEMA_signal_8989 ), .Q ( new_AGEMA_signal_8990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C ( clk ), .D ( new_AGEMA_signal_8991 ), .Q ( new_AGEMA_signal_8992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C ( clk ), .D ( new_AGEMA_signal_8993 ), .Q ( new_AGEMA_signal_8994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C ( clk ), .D ( new_AGEMA_signal_8995 ), .Q ( new_AGEMA_signal_8996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C ( clk ), .D ( new_AGEMA_signal_8997 ), .Q ( new_AGEMA_signal_8998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C ( clk ), .D ( new_AGEMA_signal_8999 ), .Q ( new_AGEMA_signal_9000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C ( clk ), .D ( new_AGEMA_signal_9001 ), .Q ( new_AGEMA_signal_9002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C ( clk ), .D ( new_AGEMA_signal_9003 ), .Q ( new_AGEMA_signal_9004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C ( clk ), .D ( new_AGEMA_signal_9005 ), .Q ( new_AGEMA_signal_9006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C ( clk ), .D ( new_AGEMA_signal_9007 ), .Q ( new_AGEMA_signal_9008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C ( clk ), .D ( new_AGEMA_signal_9009 ), .Q ( new_AGEMA_signal_9010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C ( clk ), .D ( new_AGEMA_signal_9011 ), .Q ( new_AGEMA_signal_9012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C ( clk ), .D ( new_AGEMA_signal_9013 ), .Q ( new_AGEMA_signal_9014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C ( clk ), .D ( new_AGEMA_signal_9015 ), .Q ( new_AGEMA_signal_9016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C ( clk ), .D ( new_AGEMA_signal_9017 ), .Q ( new_AGEMA_signal_9018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C ( clk ), .D ( new_AGEMA_signal_9019 ), .Q ( new_AGEMA_signal_9020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C ( clk ), .D ( new_AGEMA_signal_9021 ), .Q ( new_AGEMA_signal_9022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C ( clk ), .D ( new_AGEMA_signal_9023 ), .Q ( new_AGEMA_signal_9024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C ( clk ), .D ( new_AGEMA_signal_9025 ), .Q ( new_AGEMA_signal_9026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C ( clk ), .D ( new_AGEMA_signal_9027 ), .Q ( new_AGEMA_signal_9028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C ( clk ), .D ( new_AGEMA_signal_9029 ), .Q ( new_AGEMA_signal_9030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C ( clk ), .D ( new_AGEMA_signal_9031 ), .Q ( new_AGEMA_signal_9032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C ( clk ), .D ( new_AGEMA_signal_9033 ), .Q ( new_AGEMA_signal_9034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C ( clk ), .D ( new_AGEMA_signal_9035 ), .Q ( new_AGEMA_signal_9036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C ( clk ), .D ( new_AGEMA_signal_9037 ), .Q ( new_AGEMA_signal_9038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C ( clk ), .D ( new_AGEMA_signal_9039 ), .Q ( new_AGEMA_signal_9040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C ( clk ), .D ( new_AGEMA_signal_9041 ), .Q ( new_AGEMA_signal_9042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C ( clk ), .D ( new_AGEMA_signal_9043 ), .Q ( new_AGEMA_signal_9044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C ( clk ), .D ( new_AGEMA_signal_9045 ), .Q ( new_AGEMA_signal_9046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C ( clk ), .D ( new_AGEMA_signal_9047 ), .Q ( new_AGEMA_signal_9048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C ( clk ), .D ( new_AGEMA_signal_9049 ), .Q ( new_AGEMA_signal_9050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C ( clk ), .D ( new_AGEMA_signal_9051 ), .Q ( new_AGEMA_signal_9052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C ( clk ), .D ( new_AGEMA_signal_9053 ), .Q ( new_AGEMA_signal_9054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C ( clk ), .D ( new_AGEMA_signal_9055 ), .Q ( new_AGEMA_signal_9056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C ( clk ), .D ( new_AGEMA_signal_9057 ), .Q ( new_AGEMA_signal_9058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C ( clk ), .D ( new_AGEMA_signal_9059 ), .Q ( new_AGEMA_signal_9060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C ( clk ), .D ( new_AGEMA_signal_9061 ), .Q ( new_AGEMA_signal_9062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C ( clk ), .D ( new_AGEMA_signal_9063 ), .Q ( new_AGEMA_signal_9064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C ( clk ), .D ( new_AGEMA_signal_9065 ), .Q ( new_AGEMA_signal_9066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C ( clk ), .D ( new_AGEMA_signal_9067 ), .Q ( new_AGEMA_signal_9068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C ( clk ), .D ( new_AGEMA_signal_9069 ), .Q ( new_AGEMA_signal_9070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C ( clk ), .D ( new_AGEMA_signal_9071 ), .Q ( new_AGEMA_signal_9072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C ( clk ), .D ( new_AGEMA_signal_9073 ), .Q ( new_AGEMA_signal_9074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C ( clk ), .D ( new_AGEMA_signal_10099 ), .Q ( new_AGEMA_signal_10100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C ( clk ), .D ( new_AGEMA_signal_10105 ), .Q ( new_AGEMA_signal_10106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C ( clk ), .D ( new_AGEMA_signal_10111 ), .Q ( new_AGEMA_signal_10112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C ( clk ), .D ( new_AGEMA_signal_10117 ), .Q ( new_AGEMA_signal_10118 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1047 ( .C ( clk ), .D ( n2769 ), .Q ( new_AGEMA_signal_9075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C ( clk ), .D ( new_AGEMA_signal_1200 ), .Q ( new_AGEMA_signal_9077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C ( clk ), .D ( new_AGEMA_signal_1201 ), .Q ( new_AGEMA_signal_9079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C ( clk ), .D ( new_AGEMA_signal_1202 ), .Q ( new_AGEMA_signal_9081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C ( clk ), .D ( new_AGEMA_signal_9052 ), .Q ( new_AGEMA_signal_9083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C ( clk ), .D ( new_AGEMA_signal_9054 ), .Q ( new_AGEMA_signal_9085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C ( clk ), .D ( new_AGEMA_signal_9056 ), .Q ( new_AGEMA_signal_9087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C ( clk ), .D ( new_AGEMA_signal_9058 ), .Q ( new_AGEMA_signal_9089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C ( clk ), .D ( new_AGEMA_signal_8964 ), .Q ( new_AGEMA_signal_9091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C ( clk ), .D ( new_AGEMA_signal_8966 ), .Q ( new_AGEMA_signal_9093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C ( clk ), .D ( new_AGEMA_signal_8968 ), .Q ( new_AGEMA_signal_9095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C ( clk ), .D ( new_AGEMA_signal_8970 ), .Q ( new_AGEMA_signal_9097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C ( clk ), .D ( n2174 ), .Q ( new_AGEMA_signal_9099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C ( clk ), .D ( new_AGEMA_signal_1239 ), .Q ( new_AGEMA_signal_9101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C ( clk ), .D ( new_AGEMA_signal_1240 ), .Q ( new_AGEMA_signal_9103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C ( clk ), .D ( new_AGEMA_signal_1241 ), .Q ( new_AGEMA_signal_9105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C ( clk ), .D ( new_AGEMA_signal_8956 ), .Q ( new_AGEMA_signal_9107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C ( clk ), .D ( new_AGEMA_signal_8958 ), .Q ( new_AGEMA_signal_9109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C ( clk ), .D ( new_AGEMA_signal_8960 ), .Q ( new_AGEMA_signal_9111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C ( clk ), .D ( new_AGEMA_signal_8962 ), .Q ( new_AGEMA_signal_9113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C ( clk ), .D ( new_AGEMA_signal_8980 ), .Q ( new_AGEMA_signal_9115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C ( clk ), .D ( new_AGEMA_signal_8982 ), .Q ( new_AGEMA_signal_9117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C ( clk ), .D ( new_AGEMA_signal_8984 ), .Q ( new_AGEMA_signal_9119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C ( clk ), .D ( new_AGEMA_signal_8986 ), .Q ( new_AGEMA_signal_9121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C ( clk ), .D ( n2570 ), .Q ( new_AGEMA_signal_9123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C ( clk ), .D ( new_AGEMA_signal_1248 ), .Q ( new_AGEMA_signal_9125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C ( clk ), .D ( new_AGEMA_signal_1249 ), .Q ( new_AGEMA_signal_9127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C ( clk ), .D ( new_AGEMA_signal_1250 ), .Q ( new_AGEMA_signal_9129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C ( clk ), .D ( n2792 ), .Q ( new_AGEMA_signal_9131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C ( clk ), .D ( new_AGEMA_signal_1233 ), .Q ( new_AGEMA_signal_9133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C ( clk ), .D ( new_AGEMA_signal_1234 ), .Q ( new_AGEMA_signal_9135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C ( clk ), .D ( new_AGEMA_signal_1235 ), .Q ( new_AGEMA_signal_9137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C ( clk ), .D ( n2635 ), .Q ( new_AGEMA_signal_9139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C ( clk ), .D ( new_AGEMA_signal_990 ), .Q ( new_AGEMA_signal_9141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C ( clk ), .D ( new_AGEMA_signal_991 ), .Q ( new_AGEMA_signal_9143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C ( clk ), .D ( new_AGEMA_signal_992 ), .Q ( new_AGEMA_signal_9145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C ( clk ), .D ( n2587 ), .Q ( new_AGEMA_signal_9147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C ( clk ), .D ( new_AGEMA_signal_1095 ), .Q ( new_AGEMA_signal_9149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C ( clk ), .D ( new_AGEMA_signal_1096 ), .Q ( new_AGEMA_signal_9151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C ( clk ), .D ( new_AGEMA_signal_1097 ), .Q ( new_AGEMA_signal_9153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C ( clk ), .D ( n2725 ), .Q ( new_AGEMA_signal_9155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C ( clk ), .D ( new_AGEMA_signal_1062 ), .Q ( new_AGEMA_signal_9157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C ( clk ), .D ( new_AGEMA_signal_1063 ), .Q ( new_AGEMA_signal_9159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C ( clk ), .D ( new_AGEMA_signal_1064 ), .Q ( new_AGEMA_signal_9161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C ( clk ), .D ( n2708 ), .Q ( new_AGEMA_signal_9163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C ( clk ), .D ( new_AGEMA_signal_1008 ), .Q ( new_AGEMA_signal_9165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C ( clk ), .D ( new_AGEMA_signal_1009 ), .Q ( new_AGEMA_signal_9167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C ( clk ), .D ( new_AGEMA_signal_1010 ), .Q ( new_AGEMA_signal_9169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C ( clk ), .D ( n2818 ), .Q ( new_AGEMA_signal_9171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C ( clk ), .D ( new_AGEMA_signal_1290 ), .Q ( new_AGEMA_signal_9173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C ( clk ), .D ( new_AGEMA_signal_1291 ), .Q ( new_AGEMA_signal_9175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C ( clk ), .D ( new_AGEMA_signal_1292 ), .Q ( new_AGEMA_signal_9177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C ( clk ), .D ( n2790 ), .Q ( new_AGEMA_signal_9179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C ( clk ), .D ( new_AGEMA_signal_993 ), .Q ( new_AGEMA_signal_9181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C ( clk ), .D ( new_AGEMA_signal_994 ), .Q ( new_AGEMA_signal_9183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C ( clk ), .D ( new_AGEMA_signal_995 ), .Q ( new_AGEMA_signal_9185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C ( clk ), .D ( n2786 ), .Q ( new_AGEMA_signal_9187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C ( clk ), .D ( new_AGEMA_signal_1221 ), .Q ( new_AGEMA_signal_9189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C ( clk ), .D ( new_AGEMA_signal_1222 ), .Q ( new_AGEMA_signal_9191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C ( clk ), .D ( new_AGEMA_signal_1223 ), .Q ( new_AGEMA_signal_9193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C ( clk ), .D ( n2400 ), .Q ( new_AGEMA_signal_9195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C ( clk ), .D ( new_AGEMA_signal_1080 ), .Q ( new_AGEMA_signal_9197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C ( clk ), .D ( new_AGEMA_signal_1081 ), .Q ( new_AGEMA_signal_9199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C ( clk ), .D ( new_AGEMA_signal_1082 ), .Q ( new_AGEMA_signal_9201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C ( clk ), .D ( new_AGEMA_signal_8988 ), .Q ( new_AGEMA_signal_9203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C ( clk ), .D ( new_AGEMA_signal_8990 ), .Q ( new_AGEMA_signal_9205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C ( clk ), .D ( new_AGEMA_signal_8992 ), .Q ( new_AGEMA_signal_9207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C ( clk ), .D ( new_AGEMA_signal_8994 ), .Q ( new_AGEMA_signal_9209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C ( clk ), .D ( n2815 ), .Q ( new_AGEMA_signal_9211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C ( clk ), .D ( new_AGEMA_signal_1065 ), .Q ( new_AGEMA_signal_9213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C ( clk ), .D ( new_AGEMA_signal_1066 ), .Q ( new_AGEMA_signal_9215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C ( clk ), .D ( new_AGEMA_signal_1067 ), .Q ( new_AGEMA_signal_9217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C ( clk ), .D ( n2723 ), .Q ( new_AGEMA_signal_9219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C ( clk ), .D ( new_AGEMA_signal_1059 ), .Q ( new_AGEMA_signal_9221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C ( clk ), .D ( new_AGEMA_signal_1060 ), .Q ( new_AGEMA_signal_9223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C ( clk ), .D ( new_AGEMA_signal_1061 ), .Q ( new_AGEMA_signal_9225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C ( clk ), .D ( n2709 ), .Q ( new_AGEMA_signal_9227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C ( clk ), .D ( new_AGEMA_signal_1320 ), .Q ( new_AGEMA_signal_9229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C ( clk ), .D ( new_AGEMA_signal_1321 ), .Q ( new_AGEMA_signal_9231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C ( clk ), .D ( new_AGEMA_signal_1322 ), .Q ( new_AGEMA_signal_9233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C ( clk ), .D ( n2753 ), .Q ( new_AGEMA_signal_9235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C ( clk ), .D ( new_AGEMA_signal_1077 ), .Q ( new_AGEMA_signal_9237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C ( clk ), .D ( new_AGEMA_signal_1078 ), .Q ( new_AGEMA_signal_9239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C ( clk ), .D ( new_AGEMA_signal_1079 ), .Q ( new_AGEMA_signal_9241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C ( clk ), .D ( n2401 ), .Q ( new_AGEMA_signal_9243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C ( clk ), .D ( new_AGEMA_signal_1140 ), .Q ( new_AGEMA_signal_9245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C ( clk ), .D ( new_AGEMA_signal_1141 ), .Q ( new_AGEMA_signal_9247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C ( clk ), .D ( new_AGEMA_signal_1142 ), .Q ( new_AGEMA_signal_9249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C ( clk ), .D ( new_AGEMA_signal_9036 ), .Q ( new_AGEMA_signal_9251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C ( clk ), .D ( new_AGEMA_signal_9038 ), .Q ( new_AGEMA_signal_9253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C ( clk ), .D ( new_AGEMA_signal_9040 ), .Q ( new_AGEMA_signal_9255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C ( clk ), .D ( new_AGEMA_signal_9042 ), .Q ( new_AGEMA_signal_9257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C ( clk ), .D ( new_AGEMA_signal_8996 ), .Q ( new_AGEMA_signal_9259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C ( clk ), .D ( new_AGEMA_signal_8998 ), .Q ( new_AGEMA_signal_9261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C ( clk ), .D ( new_AGEMA_signal_9000 ), .Q ( new_AGEMA_signal_9263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C ( clk ), .D ( new_AGEMA_signal_9002 ), .Q ( new_AGEMA_signal_9265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C ( clk ), .D ( n2615 ), .Q ( new_AGEMA_signal_9267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C ( clk ), .D ( new_AGEMA_signal_1035 ), .Q ( new_AGEMA_signal_9269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C ( clk ), .D ( new_AGEMA_signal_1036 ), .Q ( new_AGEMA_signal_9271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C ( clk ), .D ( new_AGEMA_signal_1037 ), .Q ( new_AGEMA_signal_9273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C ( clk ), .D ( n2643 ), .Q ( new_AGEMA_signal_9275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C ( clk ), .D ( new_AGEMA_signal_1098 ), .Q ( new_AGEMA_signal_9277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C ( clk ), .D ( new_AGEMA_signal_1099 ), .Q ( new_AGEMA_signal_9279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C ( clk ), .D ( new_AGEMA_signal_1100 ), .Q ( new_AGEMA_signal_9281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C ( clk ), .D ( n2563 ), .Q ( new_AGEMA_signal_9283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C ( clk ), .D ( new_AGEMA_signal_1137 ), .Q ( new_AGEMA_signal_9285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C ( clk ), .D ( new_AGEMA_signal_1138 ), .Q ( new_AGEMA_signal_9287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C ( clk ), .D ( new_AGEMA_signal_1139 ), .Q ( new_AGEMA_signal_9289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C ( clk ), .D ( n2612 ), .Q ( new_AGEMA_signal_9291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C ( clk ), .D ( new_AGEMA_signal_1275 ), .Q ( new_AGEMA_signal_9293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C ( clk ), .D ( new_AGEMA_signal_1276 ), .Q ( new_AGEMA_signal_9295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C ( clk ), .D ( new_AGEMA_signal_1277 ), .Q ( new_AGEMA_signal_9297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C ( clk ), .D ( n2824 ), .Q ( new_AGEMA_signal_9299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C ( clk ), .D ( new_AGEMA_signal_1119 ), .Q ( new_AGEMA_signal_9301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C ( clk ), .D ( new_AGEMA_signal_1120 ), .Q ( new_AGEMA_signal_9303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C ( clk ), .D ( new_AGEMA_signal_1121 ), .Q ( new_AGEMA_signal_9305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C ( clk ), .D ( n2816 ), .Q ( new_AGEMA_signal_9307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C ( clk ), .D ( new_AGEMA_signal_1041 ), .Q ( new_AGEMA_signal_9309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C ( clk ), .D ( new_AGEMA_signal_1042 ), .Q ( new_AGEMA_signal_9311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C ( clk ), .D ( new_AGEMA_signal_1043 ), .Q ( new_AGEMA_signal_9313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C ( clk ), .D ( n2073 ), .Q ( new_AGEMA_signal_9315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C ( clk ), .D ( new_AGEMA_signal_1053 ), .Q ( new_AGEMA_signal_9317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C ( clk ), .D ( new_AGEMA_signal_1054 ), .Q ( new_AGEMA_signal_9319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C ( clk ), .D ( new_AGEMA_signal_1055 ), .Q ( new_AGEMA_signal_9321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C ( clk ), .D ( n2519 ), .Q ( new_AGEMA_signal_9323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C ( clk ), .D ( new_AGEMA_signal_996 ), .Q ( new_AGEMA_signal_9325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C ( clk ), .D ( new_AGEMA_signal_997 ), .Q ( new_AGEMA_signal_9327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C ( clk ), .D ( new_AGEMA_signal_998 ), .Q ( new_AGEMA_signal_9329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C ( clk ), .D ( n2616 ), .Q ( new_AGEMA_signal_9331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C ( clk ), .D ( new_AGEMA_signal_1134 ), .Q ( new_AGEMA_signal_9333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C ( clk ), .D ( new_AGEMA_signal_1135 ), .Q ( new_AGEMA_signal_9335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C ( clk ), .D ( new_AGEMA_signal_1136 ), .Q ( new_AGEMA_signal_9337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C ( clk ), .D ( new_AGEMA_signal_9044 ), .Q ( new_AGEMA_signal_9339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C ( clk ), .D ( new_AGEMA_signal_9046 ), .Q ( new_AGEMA_signal_9341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C ( clk ), .D ( new_AGEMA_signal_9048 ), .Q ( new_AGEMA_signal_9343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C ( clk ), .D ( new_AGEMA_signal_9050 ), .Q ( new_AGEMA_signal_9345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C ( clk ), .D ( n2780 ), .Q ( new_AGEMA_signal_9347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C ( clk ), .D ( new_AGEMA_signal_1044 ), .Q ( new_AGEMA_signal_9349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C ( clk ), .D ( new_AGEMA_signal_1045 ), .Q ( new_AGEMA_signal_9351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C ( clk ), .D ( new_AGEMA_signal_1046 ), .Q ( new_AGEMA_signal_9353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C ( clk ), .D ( new_AGEMA_signal_9060 ), .Q ( new_AGEMA_signal_9355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C ( clk ), .D ( new_AGEMA_signal_9062 ), .Q ( new_AGEMA_signal_9357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C ( clk ), .D ( new_AGEMA_signal_9064 ), .Q ( new_AGEMA_signal_9359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C ( clk ), .D ( new_AGEMA_signal_9066 ), .Q ( new_AGEMA_signal_9361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C ( clk ), .D ( n2742 ), .Q ( new_AGEMA_signal_9363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C ( clk ), .D ( new_AGEMA_signal_1074 ), .Q ( new_AGEMA_signal_9365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C ( clk ), .D ( new_AGEMA_signal_1075 ), .Q ( new_AGEMA_signal_9367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C ( clk ), .D ( new_AGEMA_signal_1076 ), .Q ( new_AGEMA_signal_9369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C ( clk ), .D ( n2724 ), .Q ( new_AGEMA_signal_9371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C ( clk ), .D ( new_AGEMA_signal_1236 ), .Q ( new_AGEMA_signal_9373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C ( clk ), .D ( new_AGEMA_signal_1237 ), .Q ( new_AGEMA_signal_9375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C ( clk ), .D ( new_AGEMA_signal_1238 ), .Q ( new_AGEMA_signal_9377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C ( clk ), .D ( n2317 ), .Q ( new_AGEMA_signal_9379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C ( clk ), .D ( new_AGEMA_signal_1047 ), .Q ( new_AGEMA_signal_9381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C ( clk ), .D ( new_AGEMA_signal_1048 ), .Q ( new_AGEMA_signal_9383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C ( clk ), .D ( new_AGEMA_signal_1049 ), .Q ( new_AGEMA_signal_9385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C ( clk ), .D ( n2688 ), .Q ( new_AGEMA_signal_9387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C ( clk ), .D ( new_AGEMA_signal_1209 ), .Q ( new_AGEMA_signal_9389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C ( clk ), .D ( new_AGEMA_signal_1210 ), .Q ( new_AGEMA_signal_9391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C ( clk ), .D ( new_AGEMA_signal_1211 ), .Q ( new_AGEMA_signal_9393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C ( clk ), .D ( n2609 ), .Q ( new_AGEMA_signal_9395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C ( clk ), .D ( new_AGEMA_signal_1086 ), .Q ( new_AGEMA_signal_9397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C ( clk ), .D ( new_AGEMA_signal_1087 ), .Q ( new_AGEMA_signal_9399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C ( clk ), .D ( new_AGEMA_signal_1088 ), .Q ( new_AGEMA_signal_9401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C ( clk ), .D ( n2672 ), .Q ( new_AGEMA_signal_9403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C ( clk ), .D ( new_AGEMA_signal_1185 ), .Q ( new_AGEMA_signal_9405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C ( clk ), .D ( new_AGEMA_signal_1186 ), .Q ( new_AGEMA_signal_9407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C ( clk ), .D ( new_AGEMA_signal_1187 ), .Q ( new_AGEMA_signal_9409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C ( clk ), .D ( n2640 ), .Q ( new_AGEMA_signal_9411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C ( clk ), .D ( new_AGEMA_signal_1188 ), .Q ( new_AGEMA_signal_9413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C ( clk ), .D ( new_AGEMA_signal_1189 ), .Q ( new_AGEMA_signal_9415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C ( clk ), .D ( new_AGEMA_signal_1190 ), .Q ( new_AGEMA_signal_9417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C ( clk ), .D ( n2713 ), .Q ( new_AGEMA_signal_9419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C ( clk ), .D ( new_AGEMA_signal_1056 ), .Q ( new_AGEMA_signal_9421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C ( clk ), .D ( new_AGEMA_signal_1057 ), .Q ( new_AGEMA_signal_9423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C ( clk ), .D ( new_AGEMA_signal_1058 ), .Q ( new_AGEMA_signal_9425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C ( clk ), .D ( n2777 ), .Q ( new_AGEMA_signal_9427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C ( clk ), .D ( new_AGEMA_signal_1167 ), .Q ( new_AGEMA_signal_9429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C ( clk ), .D ( new_AGEMA_signal_1168 ), .Q ( new_AGEMA_signal_9431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C ( clk ), .D ( new_AGEMA_signal_1169 ), .Q ( new_AGEMA_signal_9433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C ( clk ), .D ( n2789 ), .Q ( new_AGEMA_signal_9435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C ( clk ), .D ( new_AGEMA_signal_1197 ), .Q ( new_AGEMA_signal_9437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C ( clk ), .D ( new_AGEMA_signal_1198 ), .Q ( new_AGEMA_signal_9439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C ( clk ), .D ( new_AGEMA_signal_1199 ), .Q ( new_AGEMA_signal_9441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C ( clk ), .D ( n2661 ), .Q ( new_AGEMA_signal_9443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C ( clk ), .D ( new_AGEMA_signal_1089 ), .Q ( new_AGEMA_signal_9445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C ( clk ), .D ( new_AGEMA_signal_1090 ), .Q ( new_AGEMA_signal_9447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C ( clk ), .D ( new_AGEMA_signal_1091 ), .Q ( new_AGEMA_signal_9449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C ( clk ), .D ( new_AGEMA_signal_9012 ), .Q ( new_AGEMA_signal_9451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C ( clk ), .D ( new_AGEMA_signal_9014 ), .Q ( new_AGEMA_signal_9453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C ( clk ), .D ( new_AGEMA_signal_9016 ), .Q ( new_AGEMA_signal_9455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C ( clk ), .D ( new_AGEMA_signal_9018 ), .Q ( new_AGEMA_signal_9457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C ( clk ), .D ( n2694 ), .Q ( new_AGEMA_signal_9459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C ( clk ), .D ( new_AGEMA_signal_1050 ), .Q ( new_AGEMA_signal_9461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C ( clk ), .D ( new_AGEMA_signal_1051 ), .Q ( new_AGEMA_signal_9463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C ( clk ), .D ( new_AGEMA_signal_1052 ), .Q ( new_AGEMA_signal_9465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C ( clk ), .D ( new_AGEMA_signal_9020 ), .Q ( new_AGEMA_signal_9467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C ( clk ), .D ( new_AGEMA_signal_9022 ), .Q ( new_AGEMA_signal_9469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C ( clk ), .D ( new_AGEMA_signal_9024 ), .Q ( new_AGEMA_signal_9471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C ( clk ), .D ( new_AGEMA_signal_9026 ), .Q ( new_AGEMA_signal_9473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C ( clk ), .D ( n2682 ), .Q ( new_AGEMA_signal_9475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C ( clk ), .D ( new_AGEMA_signal_1002 ), .Q ( new_AGEMA_signal_9477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C ( clk ), .D ( new_AGEMA_signal_1003 ), .Q ( new_AGEMA_signal_9479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C ( clk ), .D ( new_AGEMA_signal_1004 ), .Q ( new_AGEMA_signal_9481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C ( clk ), .D ( new_AGEMA_signal_9068 ), .Q ( new_AGEMA_signal_9483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C ( clk ), .D ( new_AGEMA_signal_9070 ), .Q ( new_AGEMA_signal_9485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C ( clk ), .D ( new_AGEMA_signal_9072 ), .Q ( new_AGEMA_signal_9487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C ( clk ), .D ( new_AGEMA_signal_9074 ), .Q ( new_AGEMA_signal_9489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C ( clk ), .D ( n2624 ), .Q ( new_AGEMA_signal_9491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C ( clk ), .D ( new_AGEMA_signal_1125 ), .Q ( new_AGEMA_signal_9493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C ( clk ), .D ( new_AGEMA_signal_1126 ), .Q ( new_AGEMA_signal_9495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C ( clk ), .D ( new_AGEMA_signal_1127 ), .Q ( new_AGEMA_signal_9497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C ( clk ), .D ( n2356 ), .Q ( new_AGEMA_signal_9499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C ( clk ), .D ( new_AGEMA_signal_1128 ), .Q ( new_AGEMA_signal_9501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C ( clk ), .D ( new_AGEMA_signal_1129 ), .Q ( new_AGEMA_signal_9503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C ( clk ), .D ( new_AGEMA_signal_1130 ), .Q ( new_AGEMA_signal_9505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C ( clk ), .D ( n2778 ), .Q ( new_AGEMA_signal_9507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C ( clk ), .D ( new_AGEMA_signal_1107 ), .Q ( new_AGEMA_signal_9509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C ( clk ), .D ( new_AGEMA_signal_1108 ), .Q ( new_AGEMA_signal_9511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C ( clk ), .D ( new_AGEMA_signal_1109 ), .Q ( new_AGEMA_signal_9513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C ( clk ), .D ( n2766 ), .Q ( new_AGEMA_signal_9515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C ( clk ), .D ( new_AGEMA_signal_1266 ), .Q ( new_AGEMA_signal_9517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C ( clk ), .D ( new_AGEMA_signal_1267 ), .Q ( new_AGEMA_signal_9519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C ( clk ), .D ( new_AGEMA_signal_1268 ), .Q ( new_AGEMA_signal_9521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C ( clk ), .D ( n2767 ), .Q ( new_AGEMA_signal_9523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C ( clk ), .D ( new_AGEMA_signal_1194 ), .Q ( new_AGEMA_signal_9525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C ( clk ), .D ( new_AGEMA_signal_1195 ), .Q ( new_AGEMA_signal_9527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C ( clk ), .D ( new_AGEMA_signal_1196 ), .Q ( new_AGEMA_signal_9529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C ( clk ), .D ( n2641 ), .Q ( new_AGEMA_signal_9531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C ( clk ), .D ( new_AGEMA_signal_1029 ), .Q ( new_AGEMA_signal_9533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C ( clk ), .D ( new_AGEMA_signal_1030 ), .Q ( new_AGEMA_signal_9535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C ( clk ), .D ( new_AGEMA_signal_1031 ), .Q ( new_AGEMA_signal_9537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C ( clk ), .D ( n2719 ), .Q ( new_AGEMA_signal_9539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C ( clk ), .D ( new_AGEMA_signal_1026 ), .Q ( new_AGEMA_signal_9541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C ( clk ), .D ( new_AGEMA_signal_1027 ), .Q ( new_AGEMA_signal_9543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C ( clk ), .D ( new_AGEMA_signal_1028 ), .Q ( new_AGEMA_signal_9545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C ( clk ), .D ( n2707 ), .Q ( new_AGEMA_signal_9547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C ( clk ), .D ( new_AGEMA_signal_1203 ), .Q ( new_AGEMA_signal_9549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C ( clk ), .D ( new_AGEMA_signal_1204 ), .Q ( new_AGEMA_signal_9551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C ( clk ), .D ( new_AGEMA_signal_1205 ), .Q ( new_AGEMA_signal_9553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C ( clk ), .D ( n2493 ), .Q ( new_AGEMA_signal_9555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C ( clk ), .D ( new_AGEMA_signal_1092 ), .Q ( new_AGEMA_signal_9557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C ( clk ), .D ( new_AGEMA_signal_1093 ), .Q ( new_AGEMA_signal_9559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C ( clk ), .D ( new_AGEMA_signal_1094 ), .Q ( new_AGEMA_signal_9561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C ( clk ), .D ( n2577 ), .Q ( new_AGEMA_signal_9563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C ( clk ), .D ( new_AGEMA_signal_1227 ), .Q ( new_AGEMA_signal_9565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C ( clk ), .D ( new_AGEMA_signal_1228 ), .Q ( new_AGEMA_signal_9567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C ( clk ), .D ( new_AGEMA_signal_1229 ), .Q ( new_AGEMA_signal_9569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C ( clk ), .D ( n2541 ), .Q ( new_AGEMA_signal_9571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C ( clk ), .D ( new_AGEMA_signal_1212 ), .Q ( new_AGEMA_signal_9573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C ( clk ), .D ( new_AGEMA_signal_1213 ), .Q ( new_AGEMA_signal_9575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C ( clk ), .D ( new_AGEMA_signal_1214 ), .Q ( new_AGEMA_signal_9577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C ( clk ), .D ( n2679 ), .Q ( new_AGEMA_signal_9579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C ( clk ), .D ( new_AGEMA_signal_1314 ), .Q ( new_AGEMA_signal_9581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C ( clk ), .D ( new_AGEMA_signal_1315 ), .Q ( new_AGEMA_signal_9583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C ( clk ), .D ( new_AGEMA_signal_1316 ), .Q ( new_AGEMA_signal_9585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C ( clk ), .D ( n2699 ), .Q ( new_AGEMA_signal_9587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C ( clk ), .D ( new_AGEMA_signal_1038 ), .Q ( new_AGEMA_signal_9589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C ( clk ), .D ( new_AGEMA_signal_1039 ), .Q ( new_AGEMA_signal_9591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C ( clk ), .D ( new_AGEMA_signal_1040 ), .Q ( new_AGEMA_signal_9593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C ( clk ), .D ( n2611 ), .Q ( new_AGEMA_signal_9595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C ( clk ), .D ( new_AGEMA_signal_1131 ), .Q ( new_AGEMA_signal_9597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C ( clk ), .D ( new_AGEMA_signal_1132 ), .Q ( new_AGEMA_signal_9599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C ( clk ), .D ( new_AGEMA_signal_1133 ), .Q ( new_AGEMA_signal_9601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C ( clk ), .D ( n2739 ), .Q ( new_AGEMA_signal_9603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C ( clk ), .D ( new_AGEMA_signal_1101 ), .Q ( new_AGEMA_signal_9605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C ( clk ), .D ( new_AGEMA_signal_1102 ), .Q ( new_AGEMA_signal_9607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C ( clk ), .D ( new_AGEMA_signal_1103 ), .Q ( new_AGEMA_signal_9609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C ( clk ), .D ( n2772 ), .Q ( new_AGEMA_signal_9611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C ( clk ), .D ( new_AGEMA_signal_1116 ), .Q ( new_AGEMA_signal_9613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C ( clk ), .D ( new_AGEMA_signal_1117 ), .Q ( new_AGEMA_signal_9615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C ( clk ), .D ( new_AGEMA_signal_1118 ), .Q ( new_AGEMA_signal_9617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C ( clk ), .D ( n2442 ), .Q ( new_AGEMA_signal_9635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C ( clk ), .D ( new_AGEMA_signal_1251 ), .Q ( new_AGEMA_signal_9639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C ( clk ), .D ( new_AGEMA_signal_1252 ), .Q ( new_AGEMA_signal_9643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C ( clk ), .D ( new_AGEMA_signal_1253 ), .Q ( new_AGEMA_signal_9647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C ( clk ), .D ( n2779 ), .Q ( new_AGEMA_signal_9739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C ( clk ), .D ( new_AGEMA_signal_1017 ), .Q ( new_AGEMA_signal_9743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C ( clk ), .D ( new_AGEMA_signal_1018 ), .Q ( new_AGEMA_signal_9747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C ( clk ), .D ( new_AGEMA_signal_1019 ), .Q ( new_AGEMA_signal_9751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C ( clk ), .D ( n2721 ), .Q ( new_AGEMA_signal_9811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C ( clk ), .D ( new_AGEMA_signal_1149 ), .Q ( new_AGEMA_signal_9815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C ( clk ), .D ( new_AGEMA_signal_1150 ), .Q ( new_AGEMA_signal_9819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C ( clk ), .D ( new_AGEMA_signal_1151 ), .Q ( new_AGEMA_signal_9823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C ( clk ), .D ( n2823 ), .Q ( new_AGEMA_signal_9867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C ( clk ), .D ( new_AGEMA_signal_1305 ), .Q ( new_AGEMA_signal_9871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C ( clk ), .D ( new_AGEMA_signal_1306 ), .Q ( new_AGEMA_signal_9875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C ( clk ), .D ( new_AGEMA_signal_1307 ), .Q ( new_AGEMA_signal_9879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C ( clk ), .D ( n2346 ), .Q ( new_AGEMA_signal_9907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C ( clk ), .D ( new_AGEMA_signal_1155 ), .Q ( new_AGEMA_signal_9911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C ( clk ), .D ( new_AGEMA_signal_1156 ), .Q ( new_AGEMA_signal_9915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C ( clk ), .D ( new_AGEMA_signal_1157 ), .Q ( new_AGEMA_signal_9919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C ( clk ), .D ( n2315 ), .Q ( new_AGEMA_signal_9947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C ( clk ), .D ( new_AGEMA_signal_999 ), .Q ( new_AGEMA_signal_9951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C ( clk ), .D ( new_AGEMA_signal_1000 ), .Q ( new_AGEMA_signal_9955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C ( clk ), .D ( new_AGEMA_signal_1001 ), .Q ( new_AGEMA_signal_9959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C ( clk ), .D ( new_AGEMA_signal_10100 ), .Q ( new_AGEMA_signal_10101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C ( clk ), .D ( new_AGEMA_signal_10106 ), .Q ( new_AGEMA_signal_10107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C ( clk ), .D ( new_AGEMA_signal_10112 ), .Q ( new_AGEMA_signal_10113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C ( clk ), .D ( new_AGEMA_signal_10118 ), .Q ( new_AGEMA_signal_10119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C ( clk ), .D ( new_AGEMA_signal_8972 ), .Q ( new_AGEMA_signal_10147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C ( clk ), .D ( new_AGEMA_signal_8974 ), .Q ( new_AGEMA_signal_10151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C ( clk ), .D ( new_AGEMA_signal_8976 ), .Q ( new_AGEMA_signal_10155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C ( clk ), .D ( new_AGEMA_signal_8978 ), .Q ( new_AGEMA_signal_10159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C ( clk ), .D ( n2600 ), .Q ( new_AGEMA_signal_10187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C ( clk ), .D ( new_AGEMA_signal_1068 ), .Q ( new_AGEMA_signal_10191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C ( clk ), .D ( new_AGEMA_signal_1069 ), .Q ( new_AGEMA_signal_10195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C ( clk ), .D ( new_AGEMA_signal_1070 ), .Q ( new_AGEMA_signal_10199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C ( clk ), .D ( n2750 ), .Q ( new_AGEMA_signal_10259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C ( clk ), .D ( new_AGEMA_signal_1032 ), .Q ( new_AGEMA_signal_10263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C ( clk ), .D ( new_AGEMA_signal_1033 ), .Q ( new_AGEMA_signal_10267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C ( clk ), .D ( new_AGEMA_signal_1034 ), .Q ( new_AGEMA_signal_10271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C ( clk ), .D ( new_AGEMA_signal_9028 ), .Q ( new_AGEMA_signal_10291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C ( clk ), .D ( new_AGEMA_signal_9030 ), .Q ( new_AGEMA_signal_10295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C ( clk ), .D ( new_AGEMA_signal_9032 ), .Q ( new_AGEMA_signal_10299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C ( clk ), .D ( new_AGEMA_signal_9034 ), .Q ( new_AGEMA_signal_10303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C ( clk ), .D ( n2737 ), .Q ( new_AGEMA_signal_10587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C ( clk ), .D ( new_AGEMA_signal_1191 ), .Q ( new_AGEMA_signal_10593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C ( clk ), .D ( new_AGEMA_signal_1192 ), .Q ( new_AGEMA_signal_10599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C ( clk ), .D ( new_AGEMA_signal_1193 ), .Q ( new_AGEMA_signal_10605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C ( clk ), .D ( n2785 ), .Q ( new_AGEMA_signal_10691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C ( clk ), .D ( new_AGEMA_signal_1083 ), .Q ( new_AGEMA_signal_10697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C ( clk ), .D ( new_AGEMA_signal_1084 ), .Q ( new_AGEMA_signal_10703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C ( clk ), .D ( new_AGEMA_signal_1085 ), .Q ( new_AGEMA_signal_10709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3127 ( .C ( clk ), .D ( n2595 ), .Q ( new_AGEMA_signal_11155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3135 ( .C ( clk ), .D ( new_AGEMA_signal_1005 ), .Q ( new_AGEMA_signal_11163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3143 ( .C ( clk ), .D ( new_AGEMA_signal_1006 ), .Q ( new_AGEMA_signal_11171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3151 ( .C ( clk ), .D ( new_AGEMA_signal_1007 ), .Q ( new_AGEMA_signal_11179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3167 ( .C ( clk ), .D ( n2437 ), .Q ( new_AGEMA_signal_11195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3175 ( .C ( clk ), .D ( new_AGEMA_signal_1104 ), .Q ( new_AGEMA_signal_11203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3183 ( .C ( clk ), .D ( new_AGEMA_signal_1105 ), .Q ( new_AGEMA_signal_11211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3191 ( .C ( clk ), .D ( new_AGEMA_signal_1106 ), .Q ( new_AGEMA_signal_11219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3471 ( .C ( clk ), .D ( n2828 ), .Q ( new_AGEMA_signal_11499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3479 ( .C ( clk ), .D ( new_AGEMA_signal_1311 ), .Q ( new_AGEMA_signal_11507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3487 ( .C ( clk ), .D ( new_AGEMA_signal_1312 ), .Q ( new_AGEMA_signal_11515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3495 ( .C ( clk ), .D ( new_AGEMA_signal_1313 ), .Q ( new_AGEMA_signal_11523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3815 ( .C ( clk ), .D ( n2538 ), .Q ( new_AGEMA_signal_11843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3823 ( .C ( clk ), .D ( new_AGEMA_signal_1071 ), .Q ( new_AGEMA_signal_11851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3831 ( .C ( clk ), .D ( new_AGEMA_signal_1072 ), .Q ( new_AGEMA_signal_11859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3839 ( .C ( clk ), .D ( new_AGEMA_signal_1073 ), .Q ( new_AGEMA_signal_11867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3935 ( .C ( clk ), .D ( n2809 ), .Q ( new_AGEMA_signal_11963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3943 ( .C ( clk ), .D ( new_AGEMA_signal_1317 ), .Q ( new_AGEMA_signal_11971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3951 ( .C ( clk ), .D ( new_AGEMA_signal_1318 ), .Q ( new_AGEMA_signal_11979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3959 ( .C ( clk ), .D ( new_AGEMA_signal_1319 ), .Q ( new_AGEMA_signal_11987 ) ) ;

    /* cells in depth 4 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1954 ( .a ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1959 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1964 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, n1922}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1974 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1977 ( .a ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n1926}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1980 ( .a ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .b ({new_AGEMA_signal_1214, new_AGEMA_signal_1213, new_AGEMA_signal_1212, n2541}), .clk ( clk ), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, new_AGEMA_signal_1509, n1925}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1986 ( .a ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1988 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .b ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U1989 ( .a ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1992 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1997 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1226, new_AGEMA_signal_1225, new_AGEMA_signal_1224, n1930}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2005 ( .a ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .b ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2006 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2010 ( .a ({new_AGEMA_signal_8962, new_AGEMA_signal_8960, new_AGEMA_signal_8958, new_AGEMA_signal_8956}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, n1937}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2022 ( .a ({new_AGEMA_signal_8970, new_AGEMA_signal_8968, new_AGEMA_signal_8966, new_AGEMA_signal_8964}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .clk ( clk ), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n1942}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(1)) U2026 ( .a ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2030 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .b ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, n1944}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2037 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, new_AGEMA_signal_1536, n1950}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2039 ( .a ({new_AGEMA_signal_8978, new_AGEMA_signal_8976, new_AGEMA_signal_8974, new_AGEMA_signal_8972}), .b ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .clk ( clk ), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n1949}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2042 ( .a ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .b ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2043 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .b ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2047 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2053 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}), .clk ( clk ), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, n1957}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2056 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .b ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .clk ( clk ), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2062 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1115, new_AGEMA_signal_1114, new_AGEMA_signal_1113, n1964}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2063 ( .a ({new_AGEMA_signal_8986, new_AGEMA_signal_8984, new_AGEMA_signal_8982, new_AGEMA_signal_8980}), .b ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2069 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .b ({new_AGEMA_signal_8994, new_AGEMA_signal_8992, new_AGEMA_signal_8990, new_AGEMA_signal_8988}), .clk ( clk ), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2072 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2073 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2075 ( .a ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .b ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2076 ( .a ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2079 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .b ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .clk ( clk ), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2080 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2081 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2083 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .b ({new_AGEMA_signal_8994, new_AGEMA_signal_8992, new_AGEMA_signal_8990, new_AGEMA_signal_8988}), .clk ( clk ), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2086 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2087 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2091 ( .a ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .b ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2095 ( .a ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1298, new_AGEMA_signal_1297, new_AGEMA_signal_1296, n1976}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2098 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .b ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2101 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .clk ( clk ), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, n1973}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2105 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .b ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2111 ( .a ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9000, new_AGEMA_signal_8998, new_AGEMA_signal_8996}), .clk ( clk ), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2113 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, n2741}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2118 ( .a ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n1992}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2120 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, new_AGEMA_signal_1581, n1991}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2123 ( .a ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .b ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1310, new_AGEMA_signal_1309, new_AGEMA_signal_1308, n1993}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2125 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, n1995}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2132 ( .a ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .b ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2135 ( .a ({new_AGEMA_signal_9010, new_AGEMA_signal_9008, new_AGEMA_signal_9006, new_AGEMA_signal_9004}), .b ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .clk ( clk ), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2003}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2140 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, n2008}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2141 ( .a ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .clk ( clk ), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2143 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .b ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .clk ( clk ), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, n2004}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2147 ( .a ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, n2009}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2151 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9000, new_AGEMA_signal_8998, new_AGEMA_signal_8996}), .clk ( clk ), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2157 ( .a ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .b ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, n2026}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2158 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .b ({new_AGEMA_signal_1094, new_AGEMA_signal_1093, new_AGEMA_signal_1092, n2493}), .clk ( clk ), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1610, new_AGEMA_signal_1609, new_AGEMA_signal_1608, n2022}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2159 ( .a ({new_AGEMA_signal_9018, new_AGEMA_signal_9016, new_AGEMA_signal_9014, new_AGEMA_signal_9012}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2167 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9000, new_AGEMA_signal_8998, new_AGEMA_signal_8996}), .clk ( clk ), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, n2027}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2171 ( .a ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2173 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2174 ( .a ({new_AGEMA_signal_8986, new_AGEMA_signal_8984, new_AGEMA_signal_8982, new_AGEMA_signal_8980}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2178 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .clk ( clk ), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1334, new_AGEMA_signal_1333, new_AGEMA_signal_1332, n2034}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2182 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .b ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2183 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2039}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2188 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, n2042}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2191 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .b ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2192 ( .a ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .b ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .clk ( clk ), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2044}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2198 ( .a ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .b ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .clk ( clk ), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2202 ( .a ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .b ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .clk ( clk ), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2055}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2205 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, n2057}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2208 ( .a ({new_AGEMA_signal_1316, new_AGEMA_signal_1315, new_AGEMA_signal_1314, n2679}), .b ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2212 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .b ({new_AGEMA_signal_1148, new_AGEMA_signal_1147, new_AGEMA_signal_1146, n2061}), .clk ( clk ), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1655, new_AGEMA_signal_1654, new_AGEMA_signal_1653, n2062}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2216 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .b ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2220 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, n2068}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2224 ( .a ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2225 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2228 ( .a ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, n2075}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(1)) U2233 ( .a ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .b ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, new_AGEMA_signal_1344, n2081}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2234 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .b ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, n2080}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2237 ( .a ({new_AGEMA_signal_1070, new_AGEMA_signal_1069, new_AGEMA_signal_1068, n2600}), .b ({new_AGEMA_signal_1028, new_AGEMA_signal_1027, new_AGEMA_signal_1026, n2719}), .clk ( clk ), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2238 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2239 ( .a ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, n2083}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2244 ( .a ({new_AGEMA_signal_9010, new_AGEMA_signal_9008, new_AGEMA_signal_9006, new_AGEMA_signal_9004}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, n2086}), .clk ( clk ), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2247 ( .a ({new_AGEMA_signal_8986, new_AGEMA_signal_8984, new_AGEMA_signal_8982, new_AGEMA_signal_8980}), .b ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2087}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2251 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .clk ( clk ), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2260 ( .a ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .b ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, new_AGEMA_signal_1680, n2100}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2277 ( .a ({new_AGEMA_signal_1103, new_AGEMA_signal_1102, new_AGEMA_signal_1101, n2739}), .b ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .clk ( clk ), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2279 ( .a ({new_AGEMA_signal_1130, new_AGEMA_signal_1129, new_AGEMA_signal_1128, n2356}), .b ({new_AGEMA_signal_1358, new_AGEMA_signal_1357, new_AGEMA_signal_1356, n2118}), .clk ( clk ), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_1691, new_AGEMA_signal_1690, new_AGEMA_signal_1689, n2121}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2284 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .b ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, n2122}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2286 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2294 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2297 ( .a ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .b ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2132}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2304 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2305 ( .a ({new_AGEMA_signal_8962, new_AGEMA_signal_8960, new_AGEMA_signal_8958, new_AGEMA_signal_8956}), .b ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .clk ( clk ), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, new_AGEMA_signal_1716, n2138}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2312 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .b ({new_AGEMA_signal_9026, new_AGEMA_signal_9024, new_AGEMA_signal_9022, new_AGEMA_signal_9020}), .clk ( clk ), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2322 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .b ({new_AGEMA_signal_9034, new_AGEMA_signal_9032, new_AGEMA_signal_9030, new_AGEMA_signal_9028}), .clk ( clk ), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2328 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9000, new_AGEMA_signal_8998, new_AGEMA_signal_8996}), .clk ( clk ), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, n2162}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2337 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .b ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2340 ( .a ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .b ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, n2178}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2342 ( .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2176}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2343 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, n2174}), .b ({new_AGEMA_signal_9010, new_AGEMA_signal_9008, new_AGEMA_signal_9006, new_AGEMA_signal_9004}), .clk ( clk ), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, n2175}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2348 ( .a ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .b ({new_AGEMA_signal_9034, new_AGEMA_signal_9032, new_AGEMA_signal_9030, new_AGEMA_signal_9028}), .clk ( clk ), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2182}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2353 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .b ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .clk ( clk ), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2188}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2355 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .clk ( clk ), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, n2189}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2357 ( .a ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2362 ( .a ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .b ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .clk ( clk ), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2363 ( .a ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9040, new_AGEMA_signal_9038, new_AGEMA_signal_9036}), .clk ( clk ), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) U2368 ( .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2378 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .b ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, n2213}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2380 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8984, new_AGEMA_signal_8982, new_AGEMA_signal_8980}), .clk ( clk ), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2215}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2384 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .b ({new_AGEMA_signal_1202, new_AGEMA_signal_1201, new_AGEMA_signal_1200, n2769}), .clk ( clk ), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, n2218}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2386 ( .a ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2219}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2405 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, n2240}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2407 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .b ({new_AGEMA_signal_1022, new_AGEMA_signal_1021, new_AGEMA_signal_1020, n2242}), .clk ( clk ), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2408 ( .a ({new_AGEMA_signal_9010, new_AGEMA_signal_9008, new_AGEMA_signal_9006, new_AGEMA_signal_9004}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, n2243}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2411 ( .a ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .clk ( clk ), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, n2245}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2422 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .b ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .clk ( clk ), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2423 ( .a ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2259}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2426 ( .a ({new_AGEMA_signal_1016, new_AGEMA_signal_1015, new_AGEMA_signal_1014, n2261}), .b ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .clk ( clk ), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, n2262}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2431 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_1394, new_AGEMA_signal_1393, new_AGEMA_signal_1392, n2266}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2432 ( .a ({new_AGEMA_signal_1118, new_AGEMA_signal_1117, new_AGEMA_signal_1116, n2772}), .b ({new_AGEMA_signal_9034, new_AGEMA_signal_9032, new_AGEMA_signal_9030, new_AGEMA_signal_9028}), .clk ( clk ), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2436 ( .a ({new_AGEMA_signal_8962, new_AGEMA_signal_8960, new_AGEMA_signal_8958, new_AGEMA_signal_8956}), .b ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .clk ( clk ), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2268}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2443 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .clk ( clk ), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, n2278}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2448 ( .a ({new_AGEMA_signal_9050, new_AGEMA_signal_9048, new_AGEMA_signal_9046, new_AGEMA_signal_9044}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2455 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .b ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2458 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .b ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .clk ( clk ), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, n2287}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2470 ( .a ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2471 ( .a ({new_AGEMA_signal_1154, new_AGEMA_signal_1153, new_AGEMA_signal_1152, n2298}), .b ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .clk ( clk ), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2299}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2481 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .b ({new_AGEMA_signal_1280, new_AGEMA_signal_1279, new_AGEMA_signal_1278, n2313}), .clk ( clk ), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2484 ( .a ({new_AGEMA_signal_1001, new_AGEMA_signal_1000, new_AGEMA_signal_999, n2315}), .b ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2316}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2486 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .b ({new_AGEMA_signal_1049, new_AGEMA_signal_1048, new_AGEMA_signal_1047, n2317}), .clk ( clk ), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_1412, new_AGEMA_signal_1411, new_AGEMA_signal_1410, n2318}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2492 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, n2325}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2494 ( .a ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2328}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2495 ( .a ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .b ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .clk ( clk ), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, n2327}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2505 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .b ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .clk ( clk ), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, n2343}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2510 ( .a ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_1835, new_AGEMA_signal_1834, new_AGEMA_signal_1833, n2344}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) U2512 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .b ({new_AGEMA_signal_1157, new_AGEMA_signal_1156, new_AGEMA_signal_1155, n2346}), .clk ( clk ), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2348}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2513 ( .a ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, n2347}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2520 ( .a ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .b ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_1424, new_AGEMA_signal_1423, new_AGEMA_signal_1422, n2363}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2521 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .b ({new_AGEMA_signal_8994, new_AGEMA_signal_8992, new_AGEMA_signal_8990, new_AGEMA_signal_8988}), .clk ( clk ), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, n2353}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2524 ( .a ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2355}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2530 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, n2672}), .clk ( clk ), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_1853, new_AGEMA_signal_1852, new_AGEMA_signal_1851, n2364}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2543 ( .a ({new_AGEMA_signal_8962, new_AGEMA_signal_8960, new_AGEMA_signal_8958, new_AGEMA_signal_8956}), .b ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .clk ( clk ), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2558 ( .a ({new_AGEMA_signal_1124, new_AGEMA_signal_1123, new_AGEMA_signal_1122, n2395}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2563 ( .a ({new_AGEMA_signal_9058, new_AGEMA_signal_9056, new_AGEMA_signal_9054, new_AGEMA_signal_9052}), .b ({new_AGEMA_signal_1082, new_AGEMA_signal_1081, new_AGEMA_signal_1080, n2400}), .clk ( clk ), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2564 ( .a ({new_AGEMA_signal_1142, new_AGEMA_signal_1141, new_AGEMA_signal_1140, n2401}), .b ({new_AGEMA_signal_9002, new_AGEMA_signal_9000, new_AGEMA_signal_8998, new_AGEMA_signal_8996}), .clk ( clk ), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2402}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2585 ( .a ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, n2428}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2588 ( .a ({new_AGEMA_signal_1163, new_AGEMA_signal_1162, new_AGEMA_signal_1161, n2430}), .b ({new_AGEMA_signal_1250, new_AGEMA_signal_1249, new_AGEMA_signal_1248, n2570}), .clk ( clk ), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, n2431}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2594 ( .a ({new_AGEMA_signal_1106, new_AGEMA_signal_1105, new_AGEMA_signal_1104, n2437}), .b ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2599 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, n2442}), .b ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .clk ( clk ), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2443}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2606 ( .a ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .b ({new_AGEMA_signal_1088, new_AGEMA_signal_1087, new_AGEMA_signal_1086, n2609}), .clk ( clk ), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2608 ( .a ({new_AGEMA_signal_1112, new_AGEMA_signal_1111, new_AGEMA_signal_1110, n2452}), .b ({new_AGEMA_signal_9066, new_AGEMA_signal_9064, new_AGEMA_signal_9062, new_AGEMA_signal_9060}), .clk ( clk ), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_1442, new_AGEMA_signal_1441, new_AGEMA_signal_1440, n2453}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2616 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, n2463}), .clk ( clk ), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, n2464}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2620 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1076, new_AGEMA_signal_1075, new_AGEMA_signal_1074, n2742}), .clk ( clk ), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_1448, new_AGEMA_signal_1447, new_AGEMA_signal_1446, n2468}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2624 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .b ({new_AGEMA_signal_8994, new_AGEMA_signal_8992, new_AGEMA_signal_8990, new_AGEMA_signal_8988}), .clk ( clk ), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, n2473}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2625 ( .a ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2472}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2628 ( .a ({new_AGEMA_signal_1091, new_AGEMA_signal_1090, new_AGEMA_signal_1089, n2661}), .b ({new_AGEMA_signal_1178, new_AGEMA_signal_1177, new_AGEMA_signal_1176, n2474}), .clk ( clk ), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_1457, new_AGEMA_signal_1456, new_AGEMA_signal_1455, n2475}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2632 ( .a ({new_AGEMA_signal_9074, new_AGEMA_signal_9072, new_AGEMA_signal_9070, new_AGEMA_signal_9068}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, n2828}), .clk ( clk ), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, new_AGEMA_signal_1905, n2480}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2638 ( .a ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, n2577}), .b ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, n2487}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2641 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .b ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .clk ( clk ), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2488}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2665 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .b ({new_AGEMA_signal_998, new_AGEMA_signal_997, new_AGEMA_signal_996, n2519}), .clk ( clk ), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2520}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2667 ( .a ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .b ({new_AGEMA_signal_1097, new_AGEMA_signal_1096, new_AGEMA_signal_1095, n2587}), .clk ( clk ), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, n2521}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2674 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .b ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .clk ( clk ), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, n2531}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2689 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, n2553}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2691 ( .a ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .clk ( clk ), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2554}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) U2695 ( .a ({new_AGEMA_signal_1013, new_AGEMA_signal_1012, new_AGEMA_signal_1011, n2559}), .b ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2560}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2698 ( .a ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .b ({new_AGEMA_signal_1139, new_AGEMA_signal_1138, new_AGEMA_signal_1137, n2563}), .clk ( clk ), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_1943, new_AGEMA_signal_1942, new_AGEMA_signal_1941, n2564}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2714 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, n2688}), .b ({new_AGEMA_signal_1052, new_AGEMA_signal_1051, new_AGEMA_signal_1050, n2694}), .clk ( clk ), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2586}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2720 ( .a ({new_AGEMA_signal_1007, new_AGEMA_signal_1006, new_AGEMA_signal_1005, n2595}), .b ({new_AGEMA_signal_1100, new_AGEMA_signal_1099, new_AGEMA_signal_1098, n2643}), .clk ( clk ), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, n2597}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2721 ( .a ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2596}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2723 ( .a ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .b ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .clk ( clk ), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, n2598}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2725 ( .a ({new_AGEMA_signal_992, new_AGEMA_signal_991, new_AGEMA_signal_990, n2635}), .b ({new_AGEMA_signal_8986, new_AGEMA_signal_8984, new_AGEMA_signal_8982, new_AGEMA_signal_8980}), .clk ( clk ), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, n2599}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2732 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .b ({new_AGEMA_signal_1292, new_AGEMA_signal_1291, new_AGEMA_signal_1290, n2818}), .clk ( clk ), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, n2610}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2734 ( .a ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .b ({new_AGEMA_signal_1133, new_AGEMA_signal_1132, new_AGEMA_signal_1131, n2611}), .clk ( clk ), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2614}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2735 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, n2612}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, n2613}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2737 ( .a ({new_AGEMA_signal_1136, new_AGEMA_signal_1135, new_AGEMA_signal_1134, n2616}), .b ({new_AGEMA_signal_1037, new_AGEMA_signal_1036, new_AGEMA_signal_1035, n2615}), .clk ( clk ), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_1475, new_AGEMA_signal_1474, new_AGEMA_signal_1473, n2617}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2742 ( .a ({new_AGEMA_signal_1127, new_AGEMA_signal_1126, new_AGEMA_signal_1125, n2624}), .b ({new_AGEMA_signal_1034, new_AGEMA_signal_1033, new_AGEMA_signal_1032, n2750}), .clk ( clk ), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, n2629}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2751 ( .a ({new_AGEMA_signal_1031, new_AGEMA_signal_1030, new_AGEMA_signal_1029, n2641}), .b ({new_AGEMA_signal_1190, new_AGEMA_signal_1189, new_AGEMA_signal_1188, n2640}), .clk ( clk ), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2757 ( .a ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, n2650}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2775 ( .a ({new_AGEMA_signal_9026, new_AGEMA_signal_9024, new_AGEMA_signal_9022, new_AGEMA_signal_9020}), .b ({new_AGEMA_signal_1004, new_AGEMA_signal_1003, new_AGEMA_signal_1002, n2682}), .clk ( clk ), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_1184, new_AGEMA_signal_1183, new_AGEMA_signal_1182, n2683}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2789 ( .a ({new_AGEMA_signal_1061, new_AGEMA_signal_1060, new_AGEMA_signal_1059, n2723}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, n2707}), .clk ( clk ), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2711}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2790 ( .a ({new_AGEMA_signal_1322, new_AGEMA_signal_1321, new_AGEMA_signal_1320, n2709}), .b ({new_AGEMA_signal_1010, new_AGEMA_signal_1009, new_AGEMA_signal_1008, n2708}), .clk ( clk ), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, n2710}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2792 ( .a ({new_AGEMA_signal_1058, new_AGEMA_signal_1057, new_AGEMA_signal_1056, n2713}), .b ({new_AGEMA_signal_1025, new_AGEMA_signal_1024, new_AGEMA_signal_1023, n2712}), .clk ( clk ), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_1484, new_AGEMA_signal_1483, new_AGEMA_signal_1482, n2714}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2797 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_1151, new_AGEMA_signal_1150, new_AGEMA_signal_1149, n2721}), .clk ( clk ), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, n2722}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2799 ( .a ({new_AGEMA_signal_1064, new_AGEMA_signal_1063, new_AGEMA_signal_1062, n2725}), .b ({new_AGEMA_signal_1238, new_AGEMA_signal_1237, new_AGEMA_signal_1236, n2724}), .clk ( clk ), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, n2726}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2806 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, n2737}), .b ({new_AGEMA_signal_1079, new_AGEMA_signal_1078, new_AGEMA_signal_1077, n2753}), .clk ( clk ), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2738}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2822 ( .a ({new_AGEMA_signal_1196, new_AGEMA_signal_1195, new_AGEMA_signal_1194, n2767}), .b ({new_AGEMA_signal_1268, new_AGEMA_signal_1267, new_AGEMA_signal_1266, n2766}), .clk ( clk ), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, n2768}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2828 ( .a ({new_AGEMA_signal_1109, new_AGEMA_signal_1108, new_AGEMA_signal_1107, n2778}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, n2777}), .clk ( clk ), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2782}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2829 ( .a ({new_AGEMA_signal_1046, new_AGEMA_signal_1045, new_AGEMA_signal_1044, n2780}), .b ({new_AGEMA_signal_1019, new_AGEMA_signal_1018, new_AGEMA_signal_1017, n2779}), .clk ( clk ), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, n2781}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2832 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, n2786}), .b ({new_AGEMA_signal_1085, new_AGEMA_signal_1084, new_AGEMA_signal_1083, n2785}), .clk ( clk ), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, n2787}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2834 ( .a ({new_AGEMA_signal_995, new_AGEMA_signal_994, new_AGEMA_signal_993, n2790}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, n2789}), .clk ( clk ), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, new_AGEMA_signal_2028, n2794}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2835 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, n2792}), .b ({new_AGEMA_signal_9050, new_AGEMA_signal_9048, new_AGEMA_signal_9046, new_AGEMA_signal_9044}), .clk ( clk ), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, n2793}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2844 ( .a ({new_AGEMA_signal_9074, new_AGEMA_signal_9072, new_AGEMA_signal_9070, new_AGEMA_signal_9068}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, n2809}), .clk ( clk ), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2812}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2847 ( .a ({new_AGEMA_signal_1043, new_AGEMA_signal_1042, new_AGEMA_signal_1041, n2816}), .b ({new_AGEMA_signal_1067, new_AGEMA_signal_1066, new_AGEMA_signal_1065, n2815}), .clk ( clk ), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, n2820}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2851 ( .a ({new_AGEMA_signal_1121, new_AGEMA_signal_1120, new_AGEMA_signal_1119, n2824}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, n2823}), .clk ( clk ), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, n2825}) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C ( clk ), .D ( new_AGEMA_signal_9075 ), .Q ( new_AGEMA_signal_9076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C ( clk ), .D ( new_AGEMA_signal_9077 ), .Q ( new_AGEMA_signal_9078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C ( clk ), .D ( new_AGEMA_signal_9079 ), .Q ( new_AGEMA_signal_9080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C ( clk ), .D ( new_AGEMA_signal_9081 ), .Q ( new_AGEMA_signal_9082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C ( clk ), .D ( new_AGEMA_signal_9083 ), .Q ( new_AGEMA_signal_9084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C ( clk ), .D ( new_AGEMA_signal_9085 ), .Q ( new_AGEMA_signal_9086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C ( clk ), .D ( new_AGEMA_signal_9087 ), .Q ( new_AGEMA_signal_9088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C ( clk ), .D ( new_AGEMA_signal_9089 ), .Q ( new_AGEMA_signal_9090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C ( clk ), .D ( new_AGEMA_signal_9091 ), .Q ( new_AGEMA_signal_9092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C ( clk ), .D ( new_AGEMA_signal_9093 ), .Q ( new_AGEMA_signal_9094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C ( clk ), .D ( new_AGEMA_signal_9095 ), .Q ( new_AGEMA_signal_9096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C ( clk ), .D ( new_AGEMA_signal_9097 ), .Q ( new_AGEMA_signal_9098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C ( clk ), .D ( new_AGEMA_signal_9099 ), .Q ( new_AGEMA_signal_9100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C ( clk ), .D ( new_AGEMA_signal_9101 ), .Q ( new_AGEMA_signal_9102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C ( clk ), .D ( new_AGEMA_signal_9103 ), .Q ( new_AGEMA_signal_9104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C ( clk ), .D ( new_AGEMA_signal_9105 ), .Q ( new_AGEMA_signal_9106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C ( clk ), .D ( new_AGEMA_signal_9107 ), .Q ( new_AGEMA_signal_9108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C ( clk ), .D ( new_AGEMA_signal_9109 ), .Q ( new_AGEMA_signal_9110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C ( clk ), .D ( new_AGEMA_signal_9111 ), .Q ( new_AGEMA_signal_9112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C ( clk ), .D ( new_AGEMA_signal_9113 ), .Q ( new_AGEMA_signal_9114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C ( clk ), .D ( new_AGEMA_signal_9115 ), .Q ( new_AGEMA_signal_9116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C ( clk ), .D ( new_AGEMA_signal_9117 ), .Q ( new_AGEMA_signal_9118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C ( clk ), .D ( new_AGEMA_signal_9119 ), .Q ( new_AGEMA_signal_9120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C ( clk ), .D ( new_AGEMA_signal_9121 ), .Q ( new_AGEMA_signal_9122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C ( clk ), .D ( new_AGEMA_signal_9123 ), .Q ( new_AGEMA_signal_9124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C ( clk ), .D ( new_AGEMA_signal_9125 ), .Q ( new_AGEMA_signal_9126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C ( clk ), .D ( new_AGEMA_signal_9127 ), .Q ( new_AGEMA_signal_9128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C ( clk ), .D ( new_AGEMA_signal_9129 ), .Q ( new_AGEMA_signal_9130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C ( clk ), .D ( new_AGEMA_signal_9131 ), .Q ( new_AGEMA_signal_9132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C ( clk ), .D ( new_AGEMA_signal_9133 ), .Q ( new_AGEMA_signal_9134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C ( clk ), .D ( new_AGEMA_signal_9135 ), .Q ( new_AGEMA_signal_9136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C ( clk ), .D ( new_AGEMA_signal_9137 ), .Q ( new_AGEMA_signal_9138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C ( clk ), .D ( new_AGEMA_signal_9139 ), .Q ( new_AGEMA_signal_9140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C ( clk ), .D ( new_AGEMA_signal_9141 ), .Q ( new_AGEMA_signal_9142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C ( clk ), .D ( new_AGEMA_signal_9143 ), .Q ( new_AGEMA_signal_9144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C ( clk ), .D ( new_AGEMA_signal_9145 ), .Q ( new_AGEMA_signal_9146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C ( clk ), .D ( new_AGEMA_signal_9147 ), .Q ( new_AGEMA_signal_9148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C ( clk ), .D ( new_AGEMA_signal_9149 ), .Q ( new_AGEMA_signal_9150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C ( clk ), .D ( new_AGEMA_signal_9151 ), .Q ( new_AGEMA_signal_9152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C ( clk ), .D ( new_AGEMA_signal_9153 ), .Q ( new_AGEMA_signal_9154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C ( clk ), .D ( new_AGEMA_signal_9155 ), .Q ( new_AGEMA_signal_9156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C ( clk ), .D ( new_AGEMA_signal_9157 ), .Q ( new_AGEMA_signal_9158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C ( clk ), .D ( new_AGEMA_signal_9159 ), .Q ( new_AGEMA_signal_9160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C ( clk ), .D ( new_AGEMA_signal_9161 ), .Q ( new_AGEMA_signal_9162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C ( clk ), .D ( new_AGEMA_signal_9163 ), .Q ( new_AGEMA_signal_9164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C ( clk ), .D ( new_AGEMA_signal_9165 ), .Q ( new_AGEMA_signal_9166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C ( clk ), .D ( new_AGEMA_signal_9167 ), .Q ( new_AGEMA_signal_9168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C ( clk ), .D ( new_AGEMA_signal_9169 ), .Q ( new_AGEMA_signal_9170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C ( clk ), .D ( new_AGEMA_signal_9171 ), .Q ( new_AGEMA_signal_9172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C ( clk ), .D ( new_AGEMA_signal_9173 ), .Q ( new_AGEMA_signal_9174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C ( clk ), .D ( new_AGEMA_signal_9175 ), .Q ( new_AGEMA_signal_9176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C ( clk ), .D ( new_AGEMA_signal_9177 ), .Q ( new_AGEMA_signal_9178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C ( clk ), .D ( new_AGEMA_signal_9179 ), .Q ( new_AGEMA_signal_9180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C ( clk ), .D ( new_AGEMA_signal_9181 ), .Q ( new_AGEMA_signal_9182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C ( clk ), .D ( new_AGEMA_signal_9183 ), .Q ( new_AGEMA_signal_9184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C ( clk ), .D ( new_AGEMA_signal_9185 ), .Q ( new_AGEMA_signal_9186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C ( clk ), .D ( new_AGEMA_signal_9187 ), .Q ( new_AGEMA_signal_9188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C ( clk ), .D ( new_AGEMA_signal_9189 ), .Q ( new_AGEMA_signal_9190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C ( clk ), .D ( new_AGEMA_signal_9191 ), .Q ( new_AGEMA_signal_9192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C ( clk ), .D ( new_AGEMA_signal_9193 ), .Q ( new_AGEMA_signal_9194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C ( clk ), .D ( new_AGEMA_signal_9195 ), .Q ( new_AGEMA_signal_9196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C ( clk ), .D ( new_AGEMA_signal_9197 ), .Q ( new_AGEMA_signal_9198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C ( clk ), .D ( new_AGEMA_signal_9199 ), .Q ( new_AGEMA_signal_9200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C ( clk ), .D ( new_AGEMA_signal_9201 ), .Q ( new_AGEMA_signal_9202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C ( clk ), .D ( new_AGEMA_signal_9203 ), .Q ( new_AGEMA_signal_9204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C ( clk ), .D ( new_AGEMA_signal_9205 ), .Q ( new_AGEMA_signal_9206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C ( clk ), .D ( new_AGEMA_signal_9207 ), .Q ( new_AGEMA_signal_9208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C ( clk ), .D ( new_AGEMA_signal_9209 ), .Q ( new_AGEMA_signal_9210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C ( clk ), .D ( new_AGEMA_signal_9211 ), .Q ( new_AGEMA_signal_9212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C ( clk ), .D ( new_AGEMA_signal_9213 ), .Q ( new_AGEMA_signal_9214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C ( clk ), .D ( new_AGEMA_signal_9215 ), .Q ( new_AGEMA_signal_9216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C ( clk ), .D ( new_AGEMA_signal_9217 ), .Q ( new_AGEMA_signal_9218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C ( clk ), .D ( new_AGEMA_signal_9219 ), .Q ( new_AGEMA_signal_9220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C ( clk ), .D ( new_AGEMA_signal_9221 ), .Q ( new_AGEMA_signal_9222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C ( clk ), .D ( new_AGEMA_signal_9223 ), .Q ( new_AGEMA_signal_9224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C ( clk ), .D ( new_AGEMA_signal_9225 ), .Q ( new_AGEMA_signal_9226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C ( clk ), .D ( new_AGEMA_signal_9227 ), .Q ( new_AGEMA_signal_9228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C ( clk ), .D ( new_AGEMA_signal_9229 ), .Q ( new_AGEMA_signal_9230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C ( clk ), .D ( new_AGEMA_signal_9231 ), .Q ( new_AGEMA_signal_9232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C ( clk ), .D ( new_AGEMA_signal_9233 ), .Q ( new_AGEMA_signal_9234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C ( clk ), .D ( new_AGEMA_signal_9235 ), .Q ( new_AGEMA_signal_9236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C ( clk ), .D ( new_AGEMA_signal_9237 ), .Q ( new_AGEMA_signal_9238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C ( clk ), .D ( new_AGEMA_signal_9239 ), .Q ( new_AGEMA_signal_9240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C ( clk ), .D ( new_AGEMA_signal_9241 ), .Q ( new_AGEMA_signal_9242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C ( clk ), .D ( new_AGEMA_signal_9243 ), .Q ( new_AGEMA_signal_9244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C ( clk ), .D ( new_AGEMA_signal_9245 ), .Q ( new_AGEMA_signal_9246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C ( clk ), .D ( new_AGEMA_signal_9247 ), .Q ( new_AGEMA_signal_9248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C ( clk ), .D ( new_AGEMA_signal_9249 ), .Q ( new_AGEMA_signal_9250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C ( clk ), .D ( new_AGEMA_signal_9251 ), .Q ( new_AGEMA_signal_9252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C ( clk ), .D ( new_AGEMA_signal_9253 ), .Q ( new_AGEMA_signal_9254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C ( clk ), .D ( new_AGEMA_signal_9255 ), .Q ( new_AGEMA_signal_9256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C ( clk ), .D ( new_AGEMA_signal_9257 ), .Q ( new_AGEMA_signal_9258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C ( clk ), .D ( new_AGEMA_signal_9259 ), .Q ( new_AGEMA_signal_9260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C ( clk ), .D ( new_AGEMA_signal_9261 ), .Q ( new_AGEMA_signal_9262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C ( clk ), .D ( new_AGEMA_signal_9263 ), .Q ( new_AGEMA_signal_9264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C ( clk ), .D ( new_AGEMA_signal_9265 ), .Q ( new_AGEMA_signal_9266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C ( clk ), .D ( new_AGEMA_signal_9267 ), .Q ( new_AGEMA_signal_9268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C ( clk ), .D ( new_AGEMA_signal_9269 ), .Q ( new_AGEMA_signal_9270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C ( clk ), .D ( new_AGEMA_signal_9271 ), .Q ( new_AGEMA_signal_9272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C ( clk ), .D ( new_AGEMA_signal_9273 ), .Q ( new_AGEMA_signal_9274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C ( clk ), .D ( new_AGEMA_signal_9275 ), .Q ( new_AGEMA_signal_9276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C ( clk ), .D ( new_AGEMA_signal_9277 ), .Q ( new_AGEMA_signal_9278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C ( clk ), .D ( new_AGEMA_signal_9279 ), .Q ( new_AGEMA_signal_9280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C ( clk ), .D ( new_AGEMA_signal_9281 ), .Q ( new_AGEMA_signal_9282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C ( clk ), .D ( new_AGEMA_signal_9283 ), .Q ( new_AGEMA_signal_9284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C ( clk ), .D ( new_AGEMA_signal_9285 ), .Q ( new_AGEMA_signal_9286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C ( clk ), .D ( new_AGEMA_signal_9287 ), .Q ( new_AGEMA_signal_9288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C ( clk ), .D ( new_AGEMA_signal_9289 ), .Q ( new_AGEMA_signal_9290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C ( clk ), .D ( new_AGEMA_signal_9291 ), .Q ( new_AGEMA_signal_9292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C ( clk ), .D ( new_AGEMA_signal_9293 ), .Q ( new_AGEMA_signal_9294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C ( clk ), .D ( new_AGEMA_signal_9295 ), .Q ( new_AGEMA_signal_9296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C ( clk ), .D ( new_AGEMA_signal_9297 ), .Q ( new_AGEMA_signal_9298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C ( clk ), .D ( new_AGEMA_signal_9299 ), .Q ( new_AGEMA_signal_9300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C ( clk ), .D ( new_AGEMA_signal_9301 ), .Q ( new_AGEMA_signal_9302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C ( clk ), .D ( new_AGEMA_signal_9303 ), .Q ( new_AGEMA_signal_9304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C ( clk ), .D ( new_AGEMA_signal_9305 ), .Q ( new_AGEMA_signal_9306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C ( clk ), .D ( new_AGEMA_signal_9307 ), .Q ( new_AGEMA_signal_9308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C ( clk ), .D ( new_AGEMA_signal_9309 ), .Q ( new_AGEMA_signal_9310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C ( clk ), .D ( new_AGEMA_signal_9311 ), .Q ( new_AGEMA_signal_9312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C ( clk ), .D ( new_AGEMA_signal_9313 ), .Q ( new_AGEMA_signal_9314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C ( clk ), .D ( new_AGEMA_signal_9315 ), .Q ( new_AGEMA_signal_9316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C ( clk ), .D ( new_AGEMA_signal_9317 ), .Q ( new_AGEMA_signal_9318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C ( clk ), .D ( new_AGEMA_signal_9319 ), .Q ( new_AGEMA_signal_9320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C ( clk ), .D ( new_AGEMA_signal_9321 ), .Q ( new_AGEMA_signal_9322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C ( clk ), .D ( new_AGEMA_signal_9323 ), .Q ( new_AGEMA_signal_9324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C ( clk ), .D ( new_AGEMA_signal_9325 ), .Q ( new_AGEMA_signal_9326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C ( clk ), .D ( new_AGEMA_signal_9327 ), .Q ( new_AGEMA_signal_9328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C ( clk ), .D ( new_AGEMA_signal_9329 ), .Q ( new_AGEMA_signal_9330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C ( clk ), .D ( new_AGEMA_signal_9331 ), .Q ( new_AGEMA_signal_9332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C ( clk ), .D ( new_AGEMA_signal_9333 ), .Q ( new_AGEMA_signal_9334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C ( clk ), .D ( new_AGEMA_signal_9335 ), .Q ( new_AGEMA_signal_9336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C ( clk ), .D ( new_AGEMA_signal_9337 ), .Q ( new_AGEMA_signal_9338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C ( clk ), .D ( new_AGEMA_signal_9339 ), .Q ( new_AGEMA_signal_9340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C ( clk ), .D ( new_AGEMA_signal_9341 ), .Q ( new_AGEMA_signal_9342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C ( clk ), .D ( new_AGEMA_signal_9343 ), .Q ( new_AGEMA_signal_9344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C ( clk ), .D ( new_AGEMA_signal_9345 ), .Q ( new_AGEMA_signal_9346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C ( clk ), .D ( new_AGEMA_signal_9347 ), .Q ( new_AGEMA_signal_9348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C ( clk ), .D ( new_AGEMA_signal_9349 ), .Q ( new_AGEMA_signal_9350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C ( clk ), .D ( new_AGEMA_signal_9351 ), .Q ( new_AGEMA_signal_9352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C ( clk ), .D ( new_AGEMA_signal_9353 ), .Q ( new_AGEMA_signal_9354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C ( clk ), .D ( new_AGEMA_signal_9355 ), .Q ( new_AGEMA_signal_9356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C ( clk ), .D ( new_AGEMA_signal_9357 ), .Q ( new_AGEMA_signal_9358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C ( clk ), .D ( new_AGEMA_signal_9359 ), .Q ( new_AGEMA_signal_9360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C ( clk ), .D ( new_AGEMA_signal_9361 ), .Q ( new_AGEMA_signal_9362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C ( clk ), .D ( new_AGEMA_signal_9363 ), .Q ( new_AGEMA_signal_9364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C ( clk ), .D ( new_AGEMA_signal_9365 ), .Q ( new_AGEMA_signal_9366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C ( clk ), .D ( new_AGEMA_signal_9367 ), .Q ( new_AGEMA_signal_9368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C ( clk ), .D ( new_AGEMA_signal_9369 ), .Q ( new_AGEMA_signal_9370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C ( clk ), .D ( new_AGEMA_signal_9371 ), .Q ( new_AGEMA_signal_9372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C ( clk ), .D ( new_AGEMA_signal_9373 ), .Q ( new_AGEMA_signal_9374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C ( clk ), .D ( new_AGEMA_signal_9375 ), .Q ( new_AGEMA_signal_9376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C ( clk ), .D ( new_AGEMA_signal_9377 ), .Q ( new_AGEMA_signal_9378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C ( clk ), .D ( new_AGEMA_signal_9379 ), .Q ( new_AGEMA_signal_9380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C ( clk ), .D ( new_AGEMA_signal_9381 ), .Q ( new_AGEMA_signal_9382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C ( clk ), .D ( new_AGEMA_signal_9383 ), .Q ( new_AGEMA_signal_9384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C ( clk ), .D ( new_AGEMA_signal_9385 ), .Q ( new_AGEMA_signal_9386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C ( clk ), .D ( new_AGEMA_signal_9387 ), .Q ( new_AGEMA_signal_9388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C ( clk ), .D ( new_AGEMA_signal_9389 ), .Q ( new_AGEMA_signal_9390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C ( clk ), .D ( new_AGEMA_signal_9391 ), .Q ( new_AGEMA_signal_9392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C ( clk ), .D ( new_AGEMA_signal_9393 ), .Q ( new_AGEMA_signal_9394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C ( clk ), .D ( new_AGEMA_signal_9395 ), .Q ( new_AGEMA_signal_9396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C ( clk ), .D ( new_AGEMA_signal_9397 ), .Q ( new_AGEMA_signal_9398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C ( clk ), .D ( new_AGEMA_signal_9399 ), .Q ( new_AGEMA_signal_9400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C ( clk ), .D ( new_AGEMA_signal_9401 ), .Q ( new_AGEMA_signal_9402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C ( clk ), .D ( new_AGEMA_signal_9403 ), .Q ( new_AGEMA_signal_9404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C ( clk ), .D ( new_AGEMA_signal_9405 ), .Q ( new_AGEMA_signal_9406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C ( clk ), .D ( new_AGEMA_signal_9407 ), .Q ( new_AGEMA_signal_9408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C ( clk ), .D ( new_AGEMA_signal_9409 ), .Q ( new_AGEMA_signal_9410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C ( clk ), .D ( new_AGEMA_signal_9411 ), .Q ( new_AGEMA_signal_9412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C ( clk ), .D ( new_AGEMA_signal_9413 ), .Q ( new_AGEMA_signal_9414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C ( clk ), .D ( new_AGEMA_signal_9415 ), .Q ( new_AGEMA_signal_9416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C ( clk ), .D ( new_AGEMA_signal_9417 ), .Q ( new_AGEMA_signal_9418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C ( clk ), .D ( new_AGEMA_signal_9419 ), .Q ( new_AGEMA_signal_9420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C ( clk ), .D ( new_AGEMA_signal_9421 ), .Q ( new_AGEMA_signal_9422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C ( clk ), .D ( new_AGEMA_signal_9423 ), .Q ( new_AGEMA_signal_9424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C ( clk ), .D ( new_AGEMA_signal_9425 ), .Q ( new_AGEMA_signal_9426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C ( clk ), .D ( new_AGEMA_signal_9427 ), .Q ( new_AGEMA_signal_9428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C ( clk ), .D ( new_AGEMA_signal_9429 ), .Q ( new_AGEMA_signal_9430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C ( clk ), .D ( new_AGEMA_signal_9431 ), .Q ( new_AGEMA_signal_9432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C ( clk ), .D ( new_AGEMA_signal_9433 ), .Q ( new_AGEMA_signal_9434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C ( clk ), .D ( new_AGEMA_signal_9435 ), .Q ( new_AGEMA_signal_9436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C ( clk ), .D ( new_AGEMA_signal_9437 ), .Q ( new_AGEMA_signal_9438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C ( clk ), .D ( new_AGEMA_signal_9439 ), .Q ( new_AGEMA_signal_9440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C ( clk ), .D ( new_AGEMA_signal_9441 ), .Q ( new_AGEMA_signal_9442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C ( clk ), .D ( new_AGEMA_signal_9443 ), .Q ( new_AGEMA_signal_9444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C ( clk ), .D ( new_AGEMA_signal_9445 ), .Q ( new_AGEMA_signal_9446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C ( clk ), .D ( new_AGEMA_signal_9447 ), .Q ( new_AGEMA_signal_9448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C ( clk ), .D ( new_AGEMA_signal_9449 ), .Q ( new_AGEMA_signal_9450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C ( clk ), .D ( new_AGEMA_signal_9451 ), .Q ( new_AGEMA_signal_9452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C ( clk ), .D ( new_AGEMA_signal_9453 ), .Q ( new_AGEMA_signal_9454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C ( clk ), .D ( new_AGEMA_signal_9455 ), .Q ( new_AGEMA_signal_9456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C ( clk ), .D ( new_AGEMA_signal_9457 ), .Q ( new_AGEMA_signal_9458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C ( clk ), .D ( new_AGEMA_signal_9459 ), .Q ( new_AGEMA_signal_9460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C ( clk ), .D ( new_AGEMA_signal_9461 ), .Q ( new_AGEMA_signal_9462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C ( clk ), .D ( new_AGEMA_signal_9463 ), .Q ( new_AGEMA_signal_9464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C ( clk ), .D ( new_AGEMA_signal_9465 ), .Q ( new_AGEMA_signal_9466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C ( clk ), .D ( new_AGEMA_signal_9467 ), .Q ( new_AGEMA_signal_9468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C ( clk ), .D ( new_AGEMA_signal_9469 ), .Q ( new_AGEMA_signal_9470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C ( clk ), .D ( new_AGEMA_signal_9471 ), .Q ( new_AGEMA_signal_9472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C ( clk ), .D ( new_AGEMA_signal_9473 ), .Q ( new_AGEMA_signal_9474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C ( clk ), .D ( new_AGEMA_signal_9475 ), .Q ( new_AGEMA_signal_9476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C ( clk ), .D ( new_AGEMA_signal_9477 ), .Q ( new_AGEMA_signal_9478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C ( clk ), .D ( new_AGEMA_signal_9479 ), .Q ( new_AGEMA_signal_9480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C ( clk ), .D ( new_AGEMA_signal_9481 ), .Q ( new_AGEMA_signal_9482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C ( clk ), .D ( new_AGEMA_signal_9483 ), .Q ( new_AGEMA_signal_9484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C ( clk ), .D ( new_AGEMA_signal_9485 ), .Q ( new_AGEMA_signal_9486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C ( clk ), .D ( new_AGEMA_signal_9487 ), .Q ( new_AGEMA_signal_9488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C ( clk ), .D ( new_AGEMA_signal_9489 ), .Q ( new_AGEMA_signal_9490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C ( clk ), .D ( new_AGEMA_signal_9491 ), .Q ( new_AGEMA_signal_9492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C ( clk ), .D ( new_AGEMA_signal_9493 ), .Q ( new_AGEMA_signal_9494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C ( clk ), .D ( new_AGEMA_signal_9495 ), .Q ( new_AGEMA_signal_9496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C ( clk ), .D ( new_AGEMA_signal_9497 ), .Q ( new_AGEMA_signal_9498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C ( clk ), .D ( new_AGEMA_signal_9499 ), .Q ( new_AGEMA_signal_9500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C ( clk ), .D ( new_AGEMA_signal_9501 ), .Q ( new_AGEMA_signal_9502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C ( clk ), .D ( new_AGEMA_signal_9503 ), .Q ( new_AGEMA_signal_9504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C ( clk ), .D ( new_AGEMA_signal_9505 ), .Q ( new_AGEMA_signal_9506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C ( clk ), .D ( new_AGEMA_signal_9507 ), .Q ( new_AGEMA_signal_9508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C ( clk ), .D ( new_AGEMA_signal_9509 ), .Q ( new_AGEMA_signal_9510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C ( clk ), .D ( new_AGEMA_signal_9511 ), .Q ( new_AGEMA_signal_9512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C ( clk ), .D ( new_AGEMA_signal_9513 ), .Q ( new_AGEMA_signal_9514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C ( clk ), .D ( new_AGEMA_signal_9515 ), .Q ( new_AGEMA_signal_9516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C ( clk ), .D ( new_AGEMA_signal_9517 ), .Q ( new_AGEMA_signal_9518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C ( clk ), .D ( new_AGEMA_signal_9519 ), .Q ( new_AGEMA_signal_9520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C ( clk ), .D ( new_AGEMA_signal_9521 ), .Q ( new_AGEMA_signal_9522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C ( clk ), .D ( new_AGEMA_signal_9523 ), .Q ( new_AGEMA_signal_9524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C ( clk ), .D ( new_AGEMA_signal_9525 ), .Q ( new_AGEMA_signal_9526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C ( clk ), .D ( new_AGEMA_signal_9527 ), .Q ( new_AGEMA_signal_9528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C ( clk ), .D ( new_AGEMA_signal_9529 ), .Q ( new_AGEMA_signal_9530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C ( clk ), .D ( new_AGEMA_signal_9531 ), .Q ( new_AGEMA_signal_9532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C ( clk ), .D ( new_AGEMA_signal_9533 ), .Q ( new_AGEMA_signal_9534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C ( clk ), .D ( new_AGEMA_signal_9535 ), .Q ( new_AGEMA_signal_9536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C ( clk ), .D ( new_AGEMA_signal_9537 ), .Q ( new_AGEMA_signal_9538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C ( clk ), .D ( new_AGEMA_signal_9539 ), .Q ( new_AGEMA_signal_9540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C ( clk ), .D ( new_AGEMA_signal_9541 ), .Q ( new_AGEMA_signal_9542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C ( clk ), .D ( new_AGEMA_signal_9543 ), .Q ( new_AGEMA_signal_9544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C ( clk ), .D ( new_AGEMA_signal_9545 ), .Q ( new_AGEMA_signal_9546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C ( clk ), .D ( new_AGEMA_signal_9547 ), .Q ( new_AGEMA_signal_9548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C ( clk ), .D ( new_AGEMA_signal_9549 ), .Q ( new_AGEMA_signal_9550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C ( clk ), .D ( new_AGEMA_signal_9551 ), .Q ( new_AGEMA_signal_9552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C ( clk ), .D ( new_AGEMA_signal_9553 ), .Q ( new_AGEMA_signal_9554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C ( clk ), .D ( new_AGEMA_signal_9555 ), .Q ( new_AGEMA_signal_9556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C ( clk ), .D ( new_AGEMA_signal_9557 ), .Q ( new_AGEMA_signal_9558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C ( clk ), .D ( new_AGEMA_signal_9559 ), .Q ( new_AGEMA_signal_9560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C ( clk ), .D ( new_AGEMA_signal_9561 ), .Q ( new_AGEMA_signal_9562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C ( clk ), .D ( new_AGEMA_signal_9563 ), .Q ( new_AGEMA_signal_9564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C ( clk ), .D ( new_AGEMA_signal_9565 ), .Q ( new_AGEMA_signal_9566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C ( clk ), .D ( new_AGEMA_signal_9567 ), .Q ( new_AGEMA_signal_9568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C ( clk ), .D ( new_AGEMA_signal_9569 ), .Q ( new_AGEMA_signal_9570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C ( clk ), .D ( new_AGEMA_signal_9571 ), .Q ( new_AGEMA_signal_9572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C ( clk ), .D ( new_AGEMA_signal_9573 ), .Q ( new_AGEMA_signal_9574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C ( clk ), .D ( new_AGEMA_signal_9575 ), .Q ( new_AGEMA_signal_9576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C ( clk ), .D ( new_AGEMA_signal_9577 ), .Q ( new_AGEMA_signal_9578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C ( clk ), .D ( new_AGEMA_signal_9579 ), .Q ( new_AGEMA_signal_9580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C ( clk ), .D ( new_AGEMA_signal_9581 ), .Q ( new_AGEMA_signal_9582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C ( clk ), .D ( new_AGEMA_signal_9583 ), .Q ( new_AGEMA_signal_9584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C ( clk ), .D ( new_AGEMA_signal_9585 ), .Q ( new_AGEMA_signal_9586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C ( clk ), .D ( new_AGEMA_signal_9587 ), .Q ( new_AGEMA_signal_9588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C ( clk ), .D ( new_AGEMA_signal_9589 ), .Q ( new_AGEMA_signal_9590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C ( clk ), .D ( new_AGEMA_signal_9591 ), .Q ( new_AGEMA_signal_9592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C ( clk ), .D ( new_AGEMA_signal_9593 ), .Q ( new_AGEMA_signal_9594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C ( clk ), .D ( new_AGEMA_signal_9595 ), .Q ( new_AGEMA_signal_9596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C ( clk ), .D ( new_AGEMA_signal_9597 ), .Q ( new_AGEMA_signal_9598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C ( clk ), .D ( new_AGEMA_signal_9599 ), .Q ( new_AGEMA_signal_9600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C ( clk ), .D ( new_AGEMA_signal_9601 ), .Q ( new_AGEMA_signal_9602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C ( clk ), .D ( new_AGEMA_signal_9603 ), .Q ( new_AGEMA_signal_9604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C ( clk ), .D ( new_AGEMA_signal_9605 ), .Q ( new_AGEMA_signal_9606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C ( clk ), .D ( new_AGEMA_signal_9607 ), .Q ( new_AGEMA_signal_9608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C ( clk ), .D ( new_AGEMA_signal_9609 ), .Q ( new_AGEMA_signal_9610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C ( clk ), .D ( new_AGEMA_signal_9611 ), .Q ( new_AGEMA_signal_9612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C ( clk ), .D ( new_AGEMA_signal_9613 ), .Q ( new_AGEMA_signal_9614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C ( clk ), .D ( new_AGEMA_signal_9615 ), .Q ( new_AGEMA_signal_9616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C ( clk ), .D ( new_AGEMA_signal_9617 ), .Q ( new_AGEMA_signal_9618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C ( clk ), .D ( new_AGEMA_signal_9635 ), .Q ( new_AGEMA_signal_9636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C ( clk ), .D ( new_AGEMA_signal_9639 ), .Q ( new_AGEMA_signal_9640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C ( clk ), .D ( new_AGEMA_signal_9643 ), .Q ( new_AGEMA_signal_9644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C ( clk ), .D ( new_AGEMA_signal_9647 ), .Q ( new_AGEMA_signal_9648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C ( clk ), .D ( new_AGEMA_signal_9739 ), .Q ( new_AGEMA_signal_9740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C ( clk ), .D ( new_AGEMA_signal_9743 ), .Q ( new_AGEMA_signal_9744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C ( clk ), .D ( new_AGEMA_signal_9747 ), .Q ( new_AGEMA_signal_9748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C ( clk ), .D ( new_AGEMA_signal_9751 ), .Q ( new_AGEMA_signal_9752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C ( clk ), .D ( new_AGEMA_signal_9811 ), .Q ( new_AGEMA_signal_9812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C ( clk ), .D ( new_AGEMA_signal_9815 ), .Q ( new_AGEMA_signal_9816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C ( clk ), .D ( new_AGEMA_signal_9819 ), .Q ( new_AGEMA_signal_9820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C ( clk ), .D ( new_AGEMA_signal_9823 ), .Q ( new_AGEMA_signal_9824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C ( clk ), .D ( new_AGEMA_signal_9867 ), .Q ( new_AGEMA_signal_9868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C ( clk ), .D ( new_AGEMA_signal_9871 ), .Q ( new_AGEMA_signal_9872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C ( clk ), .D ( new_AGEMA_signal_9875 ), .Q ( new_AGEMA_signal_9876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C ( clk ), .D ( new_AGEMA_signal_9879 ), .Q ( new_AGEMA_signal_9880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C ( clk ), .D ( new_AGEMA_signal_9907 ), .Q ( new_AGEMA_signal_9908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C ( clk ), .D ( new_AGEMA_signal_9911 ), .Q ( new_AGEMA_signal_9912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C ( clk ), .D ( new_AGEMA_signal_9915 ), .Q ( new_AGEMA_signal_9916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C ( clk ), .D ( new_AGEMA_signal_9919 ), .Q ( new_AGEMA_signal_9920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C ( clk ), .D ( new_AGEMA_signal_9947 ), .Q ( new_AGEMA_signal_9948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C ( clk ), .D ( new_AGEMA_signal_9951 ), .Q ( new_AGEMA_signal_9952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C ( clk ), .D ( new_AGEMA_signal_9955 ), .Q ( new_AGEMA_signal_9956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C ( clk ), .D ( new_AGEMA_signal_9959 ), .Q ( new_AGEMA_signal_9960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C ( clk ), .D ( new_AGEMA_signal_10101 ), .Q ( new_AGEMA_signal_10102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C ( clk ), .D ( new_AGEMA_signal_10107 ), .Q ( new_AGEMA_signal_10108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C ( clk ), .D ( new_AGEMA_signal_10113 ), .Q ( new_AGEMA_signal_10114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C ( clk ), .D ( new_AGEMA_signal_10119 ), .Q ( new_AGEMA_signal_10120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C ( clk ), .D ( new_AGEMA_signal_10147 ), .Q ( new_AGEMA_signal_10148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C ( clk ), .D ( new_AGEMA_signal_10151 ), .Q ( new_AGEMA_signal_10152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C ( clk ), .D ( new_AGEMA_signal_10155 ), .Q ( new_AGEMA_signal_10156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C ( clk ), .D ( new_AGEMA_signal_10159 ), .Q ( new_AGEMA_signal_10160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C ( clk ), .D ( new_AGEMA_signal_10187 ), .Q ( new_AGEMA_signal_10188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C ( clk ), .D ( new_AGEMA_signal_10191 ), .Q ( new_AGEMA_signal_10192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C ( clk ), .D ( new_AGEMA_signal_10195 ), .Q ( new_AGEMA_signal_10196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C ( clk ), .D ( new_AGEMA_signal_10199 ), .Q ( new_AGEMA_signal_10200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C ( clk ), .D ( new_AGEMA_signal_10259 ), .Q ( new_AGEMA_signal_10260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C ( clk ), .D ( new_AGEMA_signal_10263 ), .Q ( new_AGEMA_signal_10264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C ( clk ), .D ( new_AGEMA_signal_10267 ), .Q ( new_AGEMA_signal_10268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C ( clk ), .D ( new_AGEMA_signal_10271 ), .Q ( new_AGEMA_signal_10272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C ( clk ), .D ( new_AGEMA_signal_10291 ), .Q ( new_AGEMA_signal_10292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C ( clk ), .D ( new_AGEMA_signal_10295 ), .Q ( new_AGEMA_signal_10296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C ( clk ), .D ( new_AGEMA_signal_10299 ), .Q ( new_AGEMA_signal_10300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C ( clk ), .D ( new_AGEMA_signal_10303 ), .Q ( new_AGEMA_signal_10304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C ( clk ), .D ( new_AGEMA_signal_10587 ), .Q ( new_AGEMA_signal_10588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C ( clk ), .D ( new_AGEMA_signal_10593 ), .Q ( new_AGEMA_signal_10594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C ( clk ), .D ( new_AGEMA_signal_10599 ), .Q ( new_AGEMA_signal_10600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C ( clk ), .D ( new_AGEMA_signal_10605 ), .Q ( new_AGEMA_signal_10606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C ( clk ), .D ( new_AGEMA_signal_10691 ), .Q ( new_AGEMA_signal_10692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C ( clk ), .D ( new_AGEMA_signal_10697 ), .Q ( new_AGEMA_signal_10698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C ( clk ), .D ( new_AGEMA_signal_10703 ), .Q ( new_AGEMA_signal_10704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C ( clk ), .D ( new_AGEMA_signal_10709 ), .Q ( new_AGEMA_signal_10710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3128 ( .C ( clk ), .D ( new_AGEMA_signal_11155 ), .Q ( new_AGEMA_signal_11156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3136 ( .C ( clk ), .D ( new_AGEMA_signal_11163 ), .Q ( new_AGEMA_signal_11164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3144 ( .C ( clk ), .D ( new_AGEMA_signal_11171 ), .Q ( new_AGEMA_signal_11172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3152 ( .C ( clk ), .D ( new_AGEMA_signal_11179 ), .Q ( new_AGEMA_signal_11180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3168 ( .C ( clk ), .D ( new_AGEMA_signal_11195 ), .Q ( new_AGEMA_signal_11196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3176 ( .C ( clk ), .D ( new_AGEMA_signal_11203 ), .Q ( new_AGEMA_signal_11204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3184 ( .C ( clk ), .D ( new_AGEMA_signal_11211 ), .Q ( new_AGEMA_signal_11212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3192 ( .C ( clk ), .D ( new_AGEMA_signal_11219 ), .Q ( new_AGEMA_signal_11220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3472 ( .C ( clk ), .D ( new_AGEMA_signal_11499 ), .Q ( new_AGEMA_signal_11500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3480 ( .C ( clk ), .D ( new_AGEMA_signal_11507 ), .Q ( new_AGEMA_signal_11508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3488 ( .C ( clk ), .D ( new_AGEMA_signal_11515 ), .Q ( new_AGEMA_signal_11516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3496 ( .C ( clk ), .D ( new_AGEMA_signal_11523 ), .Q ( new_AGEMA_signal_11524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3816 ( .C ( clk ), .D ( new_AGEMA_signal_11843 ), .Q ( new_AGEMA_signal_11844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3824 ( .C ( clk ), .D ( new_AGEMA_signal_11851 ), .Q ( new_AGEMA_signal_11852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3832 ( .C ( clk ), .D ( new_AGEMA_signal_11859 ), .Q ( new_AGEMA_signal_11860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3840 ( .C ( clk ), .D ( new_AGEMA_signal_11867 ), .Q ( new_AGEMA_signal_11868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3936 ( .C ( clk ), .D ( new_AGEMA_signal_11963 ), .Q ( new_AGEMA_signal_11964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3944 ( .C ( clk ), .D ( new_AGEMA_signal_11971 ), .Q ( new_AGEMA_signal_11972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3952 ( .C ( clk ), .D ( new_AGEMA_signal_11979 ), .Q ( new_AGEMA_signal_11980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3960 ( .C ( clk ), .D ( new_AGEMA_signal_11987 ), .Q ( new_AGEMA_signal_11988 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_1591 ( .C ( clk ), .D ( n2755 ), .Q ( new_AGEMA_signal_9619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C ( clk ), .D ( new_AGEMA_signal_1206 ), .Q ( new_AGEMA_signal_9621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C ( clk ), .D ( new_AGEMA_signal_1207 ), .Q ( new_AGEMA_signal_9623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C ( clk ), .D ( new_AGEMA_signal_1208 ), .Q ( new_AGEMA_signal_9625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C ( clk ), .D ( n2151 ), .Q ( new_AGEMA_signal_9627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C ( clk ), .D ( new_AGEMA_signal_1512 ), .Q ( new_AGEMA_signal_9629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C ( clk ), .D ( new_AGEMA_signal_1513 ), .Q ( new_AGEMA_signal_9631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C ( clk ), .D ( new_AGEMA_signal_1514 ), .Q ( new_AGEMA_signal_9633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C ( clk ), .D ( new_AGEMA_signal_9636 ), .Q ( new_AGEMA_signal_9637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C ( clk ), .D ( new_AGEMA_signal_9640 ), .Q ( new_AGEMA_signal_9641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C ( clk ), .D ( new_AGEMA_signal_9644 ), .Q ( new_AGEMA_signal_9645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C ( clk ), .D ( new_AGEMA_signal_9648 ), .Q ( new_AGEMA_signal_9649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C ( clk ), .D ( new_AGEMA_signal_9140 ), .Q ( new_AGEMA_signal_9651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C ( clk ), .D ( new_AGEMA_signal_9142 ), .Q ( new_AGEMA_signal_9653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C ( clk ), .D ( new_AGEMA_signal_9144 ), .Q ( new_AGEMA_signal_9655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C ( clk ), .D ( new_AGEMA_signal_9146 ), .Q ( new_AGEMA_signal_9657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C ( clk ), .D ( new_AGEMA_signal_9116 ), .Q ( new_AGEMA_signal_9659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C ( clk ), .D ( new_AGEMA_signal_9118 ), .Q ( new_AGEMA_signal_9661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C ( clk ), .D ( new_AGEMA_signal_9120 ), .Q ( new_AGEMA_signal_9663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C ( clk ), .D ( new_AGEMA_signal_9122 ), .Q ( new_AGEMA_signal_9665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C ( clk ), .D ( n1964 ), .Q ( new_AGEMA_signal_9667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C ( clk ), .D ( new_AGEMA_signal_1113 ), .Q ( new_AGEMA_signal_9669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C ( clk ), .D ( new_AGEMA_signal_1114 ), .Q ( new_AGEMA_signal_9671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C ( clk ), .D ( new_AGEMA_signal_1115 ), .Q ( new_AGEMA_signal_9673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C ( clk ), .D ( n2673 ), .Q ( new_AGEMA_signal_9675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C ( clk ), .D ( new_AGEMA_signal_1272 ), .Q ( new_AGEMA_signal_9677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C ( clk ), .D ( new_AGEMA_signal_1273 ), .Q ( new_AGEMA_signal_9679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C ( clk ), .D ( new_AGEMA_signal_1274 ), .Q ( new_AGEMA_signal_9681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C ( clk ), .D ( n2359 ), .Q ( new_AGEMA_signal_9683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C ( clk ), .D ( new_AGEMA_signal_1557 ), .Q ( new_AGEMA_signal_9685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C ( clk ), .D ( new_AGEMA_signal_1558 ), .Q ( new_AGEMA_signal_9687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C ( clk ), .D ( new_AGEMA_signal_1559 ), .Q ( new_AGEMA_signal_9689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C ( clk ), .D ( n1973 ), .Q ( new_AGEMA_signal_9691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C ( clk ), .D ( new_AGEMA_signal_1569 ), .Q ( new_AGEMA_signal_9693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C ( clk ), .D ( new_AGEMA_signal_1570 ), .Q ( new_AGEMA_signal_9695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C ( clk ), .D ( new_AGEMA_signal_1571 ), .Q ( new_AGEMA_signal_9697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C ( clk ), .D ( n2690 ), .Q ( new_AGEMA_signal_9699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C ( clk ), .D ( new_AGEMA_signal_1299 ), .Q ( new_AGEMA_signal_9701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C ( clk ), .D ( new_AGEMA_signal_1300 ), .Q ( new_AGEMA_signal_9703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C ( clk ), .D ( new_AGEMA_signal_1301 ), .Q ( new_AGEMA_signal_9705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C ( clk ), .D ( n2741 ), .Q ( new_AGEMA_signal_9707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C ( clk ), .D ( new_AGEMA_signal_1575 ), .Q ( new_AGEMA_signal_9709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C ( clk ), .D ( new_AGEMA_signal_1576 ), .Q ( new_AGEMA_signal_9711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C ( clk ), .D ( new_AGEMA_signal_1577 ), .Q ( new_AGEMA_signal_9713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C ( clk ), .D ( n1993 ), .Q ( new_AGEMA_signal_9715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C ( clk ), .D ( new_AGEMA_signal_1308 ), .Q ( new_AGEMA_signal_9717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C ( clk ), .D ( new_AGEMA_signal_1309 ), .Q ( new_AGEMA_signal_9719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C ( clk ), .D ( new_AGEMA_signal_1310 ), .Q ( new_AGEMA_signal_9721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C ( clk ), .D ( n2241 ), .Q ( new_AGEMA_signal_9723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C ( clk ), .D ( new_AGEMA_signal_1587 ), .Q ( new_AGEMA_signal_9725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C ( clk ), .D ( new_AGEMA_signal_1588 ), .Q ( new_AGEMA_signal_9727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C ( clk ), .D ( new_AGEMA_signal_1589 ), .Q ( new_AGEMA_signal_9729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C ( clk ), .D ( new_AGEMA_signal_9356 ), .Q ( new_AGEMA_signal_9731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C ( clk ), .D ( new_AGEMA_signal_9358 ), .Q ( new_AGEMA_signal_9733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C ( clk ), .D ( new_AGEMA_signal_9360 ), .Q ( new_AGEMA_signal_9735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C ( clk ), .D ( new_AGEMA_signal_9362 ), .Q ( new_AGEMA_signal_9737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C ( clk ), .D ( new_AGEMA_signal_9740 ), .Q ( new_AGEMA_signal_9741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C ( clk ), .D ( new_AGEMA_signal_9744 ), .Q ( new_AGEMA_signal_9745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C ( clk ), .D ( new_AGEMA_signal_9748 ), .Q ( new_AGEMA_signal_9749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C ( clk ), .D ( new_AGEMA_signal_9752 ), .Q ( new_AGEMA_signal_9753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C ( clk ), .D ( n2290 ), .Q ( new_AGEMA_signal_9755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C ( clk ), .D ( new_AGEMA_signal_1620 ), .Q ( new_AGEMA_signal_9757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C ( clk ), .D ( new_AGEMA_signal_1621 ), .Q ( new_AGEMA_signal_9759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C ( clk ), .D ( new_AGEMA_signal_1622 ), .Q ( new_AGEMA_signal_9761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C ( clk ), .D ( n2171 ), .Q ( new_AGEMA_signal_9763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C ( clk ), .D ( new_AGEMA_signal_1335 ), .Q ( new_AGEMA_signal_9765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C ( clk ), .D ( new_AGEMA_signal_1336 ), .Q ( new_AGEMA_signal_9767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C ( clk ), .D ( new_AGEMA_signal_1337 ), .Q ( new_AGEMA_signal_9769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C ( clk ), .D ( n2042 ), .Q ( new_AGEMA_signal_9771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C ( clk ), .D ( new_AGEMA_signal_1632 ), .Q ( new_AGEMA_signal_9773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C ( clk ), .D ( new_AGEMA_signal_1633 ), .Q ( new_AGEMA_signal_9775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C ( clk ), .D ( new_AGEMA_signal_1634 ), .Q ( new_AGEMA_signal_9777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C ( clk ), .D ( n2754 ), .Q ( new_AGEMA_signal_9779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C ( clk ), .D ( new_AGEMA_signal_1635 ), .Q ( new_AGEMA_signal_9781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C ( clk ), .D ( new_AGEMA_signal_1636 ), .Q ( new_AGEMA_signal_9783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C ( clk ), .D ( new_AGEMA_signal_1637 ), .Q ( new_AGEMA_signal_9785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C ( clk ), .D ( new_AGEMA_signal_9076 ), .Q ( new_AGEMA_signal_9787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C ( clk ), .D ( new_AGEMA_signal_9078 ), .Q ( new_AGEMA_signal_9789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C ( clk ), .D ( new_AGEMA_signal_9080 ), .Q ( new_AGEMA_signal_9791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C ( clk ), .D ( new_AGEMA_signal_9082 ), .Q ( new_AGEMA_signal_9793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C ( clk ), .D ( n2535 ), .Q ( new_AGEMA_signal_9795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C ( clk ), .D ( new_AGEMA_signal_1566 ), .Q ( new_AGEMA_signal_9797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C ( clk ), .D ( new_AGEMA_signal_1567 ), .Q ( new_AGEMA_signal_9799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C ( clk ), .D ( new_AGEMA_signal_1568 ), .Q ( new_AGEMA_signal_9801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C ( clk ), .D ( n2642 ), .Q ( new_AGEMA_signal_9803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C ( clk ), .D ( new_AGEMA_signal_1338 ), .Q ( new_AGEMA_signal_9805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C ( clk ), .D ( new_AGEMA_signal_1339 ), .Q ( new_AGEMA_signal_9807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C ( clk ), .D ( new_AGEMA_signal_1340 ), .Q ( new_AGEMA_signal_9809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C ( clk ), .D ( new_AGEMA_signal_9812 ), .Q ( new_AGEMA_signal_9813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C ( clk ), .D ( new_AGEMA_signal_9816 ), .Q ( new_AGEMA_signal_9817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C ( clk ), .D ( new_AGEMA_signal_9820 ), .Q ( new_AGEMA_signal_9821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C ( clk ), .D ( new_AGEMA_signal_9824 ), .Q ( new_AGEMA_signal_9825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C ( clk ), .D ( n2773 ), .Q ( new_AGEMA_signal_9827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C ( clk ), .D ( new_AGEMA_signal_1668 ), .Q ( new_AGEMA_signal_9829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C ( clk ), .D ( new_AGEMA_signal_1669 ), .Q ( new_AGEMA_signal_9831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C ( clk ), .D ( new_AGEMA_signal_1670 ), .Q ( new_AGEMA_signal_9833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C ( clk ), .D ( n2627 ), .Q ( new_AGEMA_signal_9835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C ( clk ), .D ( new_AGEMA_signal_1260 ), .Q ( new_AGEMA_signal_9837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C ( clk ), .D ( new_AGEMA_signal_1261 ), .Q ( new_AGEMA_signal_9839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C ( clk ), .D ( new_AGEMA_signal_1262 ), .Q ( new_AGEMA_signal_9841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C ( clk ), .D ( new_AGEMA_signal_9236 ), .Q ( new_AGEMA_signal_9843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C ( clk ), .D ( new_AGEMA_signal_9238 ), .Q ( new_AGEMA_signal_9845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C ( clk ), .D ( new_AGEMA_signal_9240 ), .Q ( new_AGEMA_signal_9847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C ( clk ), .D ( new_AGEMA_signal_9242 ), .Q ( new_AGEMA_signal_9849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C ( clk ), .D ( n2631 ), .Q ( new_AGEMA_signal_9851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C ( clk ), .D ( new_AGEMA_signal_1218 ), .Q ( new_AGEMA_signal_9853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C ( clk ), .D ( new_AGEMA_signal_1219 ), .Q ( new_AGEMA_signal_9855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C ( clk ), .D ( new_AGEMA_signal_1220 ), .Q ( new_AGEMA_signal_9857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C ( clk ), .D ( n2376 ), .Q ( new_AGEMA_signal_9859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C ( clk ), .D ( new_AGEMA_signal_1623 ), .Q ( new_AGEMA_signal_9861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C ( clk ), .D ( new_AGEMA_signal_1624 ), .Q ( new_AGEMA_signal_9863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C ( clk ), .D ( new_AGEMA_signal_1625 ), .Q ( new_AGEMA_signal_9865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C ( clk ), .D ( new_AGEMA_signal_9868 ), .Q ( new_AGEMA_signal_9869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C ( clk ), .D ( new_AGEMA_signal_9872 ), .Q ( new_AGEMA_signal_9873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C ( clk ), .D ( new_AGEMA_signal_9876 ), .Q ( new_AGEMA_signal_9877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C ( clk ), .D ( new_AGEMA_signal_9880 ), .Q ( new_AGEMA_signal_9881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C ( clk ), .D ( new_AGEMA_signal_9420 ), .Q ( new_AGEMA_signal_9883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C ( clk ), .D ( new_AGEMA_signal_9422 ), .Q ( new_AGEMA_signal_9885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C ( clk ), .D ( new_AGEMA_signal_9424 ), .Q ( new_AGEMA_signal_9887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C ( clk ), .D ( new_AGEMA_signal_9426 ), .Q ( new_AGEMA_signal_9889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C ( clk ), .D ( new_AGEMA_signal_9276 ), .Q ( new_AGEMA_signal_9891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C ( clk ), .D ( new_AGEMA_signal_9278 ), .Q ( new_AGEMA_signal_9893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C ( clk ), .D ( new_AGEMA_signal_9280 ), .Q ( new_AGEMA_signal_9895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C ( clk ), .D ( new_AGEMA_signal_9282 ), .Q ( new_AGEMA_signal_9897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C ( clk ), .D ( new_AGEMA_signal_9308 ), .Q ( new_AGEMA_signal_9899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C ( clk ), .D ( new_AGEMA_signal_9310 ), .Q ( new_AGEMA_signal_9901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C ( clk ), .D ( new_AGEMA_signal_9312 ), .Q ( new_AGEMA_signal_9903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C ( clk ), .D ( new_AGEMA_signal_9314 ), .Q ( new_AGEMA_signal_9905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C ( clk ), .D ( new_AGEMA_signal_9908 ), .Q ( new_AGEMA_signal_9909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C ( clk ), .D ( new_AGEMA_signal_9912 ), .Q ( new_AGEMA_signal_9913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C ( clk ), .D ( new_AGEMA_signal_9916 ), .Q ( new_AGEMA_signal_9917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C ( clk ), .D ( new_AGEMA_signal_9920 ), .Q ( new_AGEMA_signal_9921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C ( clk ), .D ( new_AGEMA_signal_9580 ), .Q ( new_AGEMA_signal_9923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C ( clk ), .D ( new_AGEMA_signal_9582 ), .Q ( new_AGEMA_signal_9925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C ( clk ), .D ( new_AGEMA_signal_9584 ), .Q ( new_AGEMA_signal_9927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C ( clk ), .D ( new_AGEMA_signal_9586 ), .Q ( new_AGEMA_signal_9929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C ( clk ), .D ( n2498 ), .Q ( new_AGEMA_signal_9931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C ( clk ), .D ( new_AGEMA_signal_1347 ), .Q ( new_AGEMA_signal_9933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C ( clk ), .D ( new_AGEMA_signal_1348 ), .Q ( new_AGEMA_signal_9935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C ( clk ), .D ( new_AGEMA_signal_1349 ), .Q ( new_AGEMA_signal_9937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C ( clk ), .D ( n2178 ), .Q ( new_AGEMA_signal_9939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C ( clk ), .D ( new_AGEMA_signal_1371 ), .Q ( new_AGEMA_signal_9941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C ( clk ), .D ( new_AGEMA_signal_1372 ), .Q ( new_AGEMA_signal_9943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C ( clk ), .D ( new_AGEMA_signal_1373 ), .Q ( new_AGEMA_signal_9945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C ( clk ), .D ( new_AGEMA_signal_9948 ), .Q ( new_AGEMA_signal_9949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C ( clk ), .D ( new_AGEMA_signal_9952 ), .Q ( new_AGEMA_signal_9953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C ( clk ), .D ( new_AGEMA_signal_9956 ), .Q ( new_AGEMA_signal_9957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C ( clk ), .D ( new_AGEMA_signal_9960 ), .Q ( new_AGEMA_signal_9961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C ( clk ), .D ( n2505 ), .Q ( new_AGEMA_signal_9963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C ( clk ), .D ( new_AGEMA_signal_1554 ), .Q ( new_AGEMA_signal_9965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C ( clk ), .D ( new_AGEMA_signal_1555 ), .Q ( new_AGEMA_signal_9967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C ( clk ), .D ( new_AGEMA_signal_1556 ), .Q ( new_AGEMA_signal_9969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C ( clk ), .D ( n2540 ), .Q ( new_AGEMA_signal_9971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C ( clk ), .D ( new_AGEMA_signal_1779 ), .Q ( new_AGEMA_signal_9973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C ( clk ), .D ( new_AGEMA_signal_1780 ), .Q ( new_AGEMA_signal_9975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C ( clk ), .D ( new_AGEMA_signal_1781 ), .Q ( new_AGEMA_signal_9977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C ( clk ), .D ( n2266 ), .Q ( new_AGEMA_signal_9979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C ( clk ), .D ( new_AGEMA_signal_1392 ), .Q ( new_AGEMA_signal_9981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C ( clk ), .D ( new_AGEMA_signal_1393 ), .Q ( new_AGEMA_signal_9983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C ( clk ), .D ( new_AGEMA_signal_1394 ), .Q ( new_AGEMA_signal_9985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C ( clk ), .D ( n2278 ), .Q ( new_AGEMA_signal_9987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C ( clk ), .D ( new_AGEMA_signal_1791 ), .Q ( new_AGEMA_signal_9989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C ( clk ), .D ( new_AGEMA_signal_1792 ), .Q ( new_AGEMA_signal_9991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C ( clk ), .D ( new_AGEMA_signal_1793 ), .Q ( new_AGEMA_signal_9993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C ( clk ), .D ( new_AGEMA_signal_9404 ), .Q ( new_AGEMA_signal_9995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C ( clk ), .D ( new_AGEMA_signal_9406 ), .Q ( new_AGEMA_signal_9997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C ( clk ), .D ( new_AGEMA_signal_9408 ), .Q ( new_AGEMA_signal_9999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C ( clk ), .D ( new_AGEMA_signal_9410 ), .Q ( new_AGEMA_signal_10001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C ( clk ), .D ( new_AGEMA_signal_9492 ), .Q ( new_AGEMA_signal_10003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C ( clk ), .D ( new_AGEMA_signal_9494 ), .Q ( new_AGEMA_signal_10005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C ( clk ), .D ( new_AGEMA_signal_9496 ), .Q ( new_AGEMA_signal_10007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C ( clk ), .D ( new_AGEMA_signal_9498 ), .Q ( new_AGEMA_signal_10009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C ( clk ), .D ( new_AGEMA_signal_9220 ), .Q ( new_AGEMA_signal_10011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C ( clk ), .D ( new_AGEMA_signal_9222 ), .Q ( new_AGEMA_signal_10013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C ( clk ), .D ( new_AGEMA_signal_9224 ), .Q ( new_AGEMA_signal_10015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C ( clk ), .D ( new_AGEMA_signal_9226 ), .Q ( new_AGEMA_signal_10017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C ( clk ), .D ( new_AGEMA_signal_9204 ), .Q ( new_AGEMA_signal_10019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C ( clk ), .D ( new_AGEMA_signal_9206 ), .Q ( new_AGEMA_signal_10021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C ( clk ), .D ( new_AGEMA_signal_9208 ), .Q ( new_AGEMA_signal_10023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C ( clk ), .D ( new_AGEMA_signal_9210 ), .Q ( new_AGEMA_signal_10025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C ( clk ), .D ( n2318 ), .Q ( new_AGEMA_signal_10027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C ( clk ), .D ( new_AGEMA_signal_1410 ), .Q ( new_AGEMA_signal_10029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C ( clk ), .D ( new_AGEMA_signal_1411 ), .Q ( new_AGEMA_signal_10031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C ( clk ), .D ( new_AGEMA_signal_1412 ), .Q ( new_AGEMA_signal_10033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C ( clk ), .D ( n2325 ), .Q ( new_AGEMA_signal_10035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C ( clk ), .D ( new_AGEMA_signal_1821 ), .Q ( new_AGEMA_signal_10037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C ( clk ), .D ( new_AGEMA_signal_1822 ), .Q ( new_AGEMA_signal_10039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C ( clk ), .D ( new_AGEMA_signal_1823 ), .Q ( new_AGEMA_signal_10041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C ( clk ), .D ( n2677 ), .Q ( new_AGEMA_signal_10043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C ( clk ), .D ( new_AGEMA_signal_1257 ), .Q ( new_AGEMA_signal_10045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C ( clk ), .D ( new_AGEMA_signal_1258 ), .Q ( new_AGEMA_signal_10047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C ( clk ), .D ( new_AGEMA_signal_1259 ), .Q ( new_AGEMA_signal_10049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C ( clk ), .D ( new_AGEMA_signal_9564 ), .Q ( new_AGEMA_signal_10051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C ( clk ), .D ( new_AGEMA_signal_9566 ), .Q ( new_AGEMA_signal_10053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C ( clk ), .D ( new_AGEMA_signal_9568 ), .Q ( new_AGEMA_signal_10055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C ( clk ), .D ( new_AGEMA_signal_9570 ), .Q ( new_AGEMA_signal_10057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C ( clk ), .D ( new_AGEMA_signal_9596 ), .Q ( new_AGEMA_signal_10059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C ( clk ), .D ( new_AGEMA_signal_9598 ), .Q ( new_AGEMA_signal_10061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C ( clk ), .D ( new_AGEMA_signal_9600 ), .Q ( new_AGEMA_signal_10063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C ( clk ), .D ( new_AGEMA_signal_9602 ), .Q ( new_AGEMA_signal_10065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C ( clk ), .D ( new_AGEMA_signal_9292 ), .Q ( new_AGEMA_signal_10067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C ( clk ), .D ( new_AGEMA_signal_9294 ), .Q ( new_AGEMA_signal_10069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C ( clk ), .D ( new_AGEMA_signal_9296 ), .Q ( new_AGEMA_signal_10071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C ( clk ), .D ( new_AGEMA_signal_9298 ), .Q ( new_AGEMA_signal_10073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C ( clk ), .D ( new_AGEMA_signal_9092 ), .Q ( new_AGEMA_signal_10075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C ( clk ), .D ( new_AGEMA_signal_9094 ), .Q ( new_AGEMA_signal_10077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C ( clk ), .D ( new_AGEMA_signal_9096 ), .Q ( new_AGEMA_signal_10079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C ( clk ), .D ( new_AGEMA_signal_9098 ), .Q ( new_AGEMA_signal_10081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C ( clk ), .D ( n2625 ), .Q ( new_AGEMA_signal_10083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C ( clk ), .D ( new_AGEMA_signal_1560 ), .Q ( new_AGEMA_signal_10085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C ( clk ), .D ( new_AGEMA_signal_1561 ), .Q ( new_AGEMA_signal_10087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C ( clk ), .D ( new_AGEMA_signal_1562 ), .Q ( new_AGEMA_signal_10089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C ( clk ), .D ( n2431 ), .Q ( new_AGEMA_signal_10091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C ( clk ), .D ( new_AGEMA_signal_1884 ), .Q ( new_AGEMA_signal_10093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C ( clk ), .D ( new_AGEMA_signal_1885 ), .Q ( new_AGEMA_signal_10095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C ( clk ), .D ( new_AGEMA_signal_1886 ), .Q ( new_AGEMA_signal_10097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C ( clk ), .D ( new_AGEMA_signal_10102 ), .Q ( new_AGEMA_signal_10103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C ( clk ), .D ( new_AGEMA_signal_10108 ), .Q ( new_AGEMA_signal_10109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C ( clk ), .D ( new_AGEMA_signal_10114 ), .Q ( new_AGEMA_signal_10115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C ( clk ), .D ( new_AGEMA_signal_10120 ), .Q ( new_AGEMA_signal_10121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C ( clk ), .D ( n2453 ), .Q ( new_AGEMA_signal_10123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C ( clk ), .D ( new_AGEMA_signal_1440 ), .Q ( new_AGEMA_signal_10125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C ( clk ), .D ( new_AGEMA_signal_1441 ), .Q ( new_AGEMA_signal_10127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C ( clk ), .D ( new_AGEMA_signal_1442 ), .Q ( new_AGEMA_signal_10129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C ( clk ), .D ( n2475 ), .Q ( new_AGEMA_signal_10131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C ( clk ), .D ( new_AGEMA_signal_1455 ), .Q ( new_AGEMA_signal_10133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C ( clk ), .D ( new_AGEMA_signal_1456 ), .Q ( new_AGEMA_signal_10135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C ( clk ), .D ( new_AGEMA_signal_1457 ), .Q ( new_AGEMA_signal_10137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C ( clk ), .D ( n2487 ), .Q ( new_AGEMA_signal_10139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C ( clk ), .D ( new_AGEMA_signal_1908 ), .Q ( new_AGEMA_signal_10141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C ( clk ), .D ( new_AGEMA_signal_1909 ), .Q ( new_AGEMA_signal_10143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C ( clk ), .D ( new_AGEMA_signal_1910 ), .Q ( new_AGEMA_signal_10145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C ( clk ), .D ( new_AGEMA_signal_10148 ), .Q ( new_AGEMA_signal_10149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C ( clk ), .D ( new_AGEMA_signal_10152 ), .Q ( new_AGEMA_signal_10153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C ( clk ), .D ( new_AGEMA_signal_10156 ), .Q ( new_AGEMA_signal_10157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C ( clk ), .D ( new_AGEMA_signal_10160 ), .Q ( new_AGEMA_signal_10161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C ( clk ), .D ( new_AGEMA_signal_9372 ), .Q ( new_AGEMA_signal_10163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C ( clk ), .D ( new_AGEMA_signal_9374 ), .Q ( new_AGEMA_signal_10165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C ( clk ), .D ( new_AGEMA_signal_9376 ), .Q ( new_AGEMA_signal_10167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C ( clk ), .D ( new_AGEMA_signal_9378 ), .Q ( new_AGEMA_signal_10169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C ( clk ), .D ( new_AGEMA_signal_9388 ), .Q ( new_AGEMA_signal_10171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C ( clk ), .D ( new_AGEMA_signal_9390 ), .Q ( new_AGEMA_signal_10173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C ( clk ), .D ( new_AGEMA_signal_9392 ), .Q ( new_AGEMA_signal_10175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C ( clk ), .D ( new_AGEMA_signal_9394 ), .Q ( new_AGEMA_signal_10177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C ( clk ), .D ( n2564 ), .Q ( new_AGEMA_signal_10179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C ( clk ), .D ( new_AGEMA_signal_1941 ), .Q ( new_AGEMA_signal_10181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C ( clk ), .D ( new_AGEMA_signal_1942 ), .Q ( new_AGEMA_signal_10183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C ( clk ), .D ( new_AGEMA_signal_1943 ), .Q ( new_AGEMA_signal_10185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C ( clk ), .D ( new_AGEMA_signal_10188 ), .Q ( new_AGEMA_signal_10189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C ( clk ), .D ( new_AGEMA_signal_10192 ), .Q ( new_AGEMA_signal_10193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C ( clk ), .D ( new_AGEMA_signal_10196 ), .Q ( new_AGEMA_signal_10197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C ( clk ), .D ( new_AGEMA_signal_10200 ), .Q ( new_AGEMA_signal_10201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C ( clk ), .D ( n2617 ), .Q ( new_AGEMA_signal_10203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C ( clk ), .D ( new_AGEMA_signal_1473 ), .Q ( new_AGEMA_signal_10205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C ( clk ), .D ( new_AGEMA_signal_1474 ), .Q ( new_AGEMA_signal_10207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C ( clk ), .D ( new_AGEMA_signal_1475 ), .Q ( new_AGEMA_signal_10209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C ( clk ), .D ( n2647 ), .Q ( new_AGEMA_signal_10211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C ( clk ), .D ( new_AGEMA_signal_1359 ), .Q ( new_AGEMA_signal_10213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C ( clk ), .D ( new_AGEMA_signal_1360 ), .Q ( new_AGEMA_signal_10215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C ( clk ), .D ( new_AGEMA_signal_1361 ), .Q ( new_AGEMA_signal_10217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C ( clk ), .D ( n2674 ), .Q ( new_AGEMA_signal_10219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C ( clk ), .D ( new_AGEMA_signal_2241 ), .Q ( new_AGEMA_signal_10221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C ( clk ), .D ( new_AGEMA_signal_2242 ), .Q ( new_AGEMA_signal_10223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C ( clk ), .D ( new_AGEMA_signal_2243 ), .Q ( new_AGEMA_signal_10225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C ( clk ), .D ( n2683 ), .Q ( new_AGEMA_signal_10227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C ( clk ), .D ( new_AGEMA_signal_1182 ), .Q ( new_AGEMA_signal_10229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C ( clk ), .D ( new_AGEMA_signal_1183 ), .Q ( new_AGEMA_signal_10231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C ( clk ), .D ( new_AGEMA_signal_1184 ), .Q ( new_AGEMA_signal_10233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C ( clk ), .D ( n2714 ), .Q ( new_AGEMA_signal_10235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C ( clk ), .D ( new_AGEMA_signal_1482 ), .Q ( new_AGEMA_signal_10237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C ( clk ), .D ( new_AGEMA_signal_1483 ), .Q ( new_AGEMA_signal_10239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C ( clk ), .D ( new_AGEMA_signal_1484 ), .Q ( new_AGEMA_signal_10241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C ( clk ), .D ( n2726 ), .Q ( new_AGEMA_signal_10243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C ( clk ), .D ( new_AGEMA_signal_2007 ), .Q ( new_AGEMA_signal_10245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C ( clk ), .D ( new_AGEMA_signal_2008 ), .Q ( new_AGEMA_signal_10247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C ( clk ), .D ( new_AGEMA_signal_2009 ), .Q ( new_AGEMA_signal_10249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C ( clk ), .D ( n2734 ), .Q ( new_AGEMA_signal_10251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C ( clk ), .D ( new_AGEMA_signal_1515 ), .Q ( new_AGEMA_signal_10253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C ( clk ), .D ( new_AGEMA_signal_1516 ), .Q ( new_AGEMA_signal_10255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C ( clk ), .D ( new_AGEMA_signal_1517 ), .Q ( new_AGEMA_signal_10257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C ( clk ), .D ( new_AGEMA_signal_10260 ), .Q ( new_AGEMA_signal_10261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C ( clk ), .D ( new_AGEMA_signal_10264 ), .Q ( new_AGEMA_signal_10265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C ( clk ), .D ( new_AGEMA_signal_10268 ), .Q ( new_AGEMA_signal_10269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C ( clk ), .D ( new_AGEMA_signal_10272 ), .Q ( new_AGEMA_signal_10273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C ( clk ), .D ( n2763 ), .Q ( new_AGEMA_signal_10275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C ( clk ), .D ( new_AGEMA_signal_1518 ), .Q ( new_AGEMA_signal_10277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C ( clk ), .D ( new_AGEMA_signal_1519 ), .Q ( new_AGEMA_signal_10279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C ( clk ), .D ( new_AGEMA_signal_1520 ), .Q ( new_AGEMA_signal_10281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C ( clk ), .D ( n2784 ), .Q ( new_AGEMA_signal_10283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C ( clk ), .D ( new_AGEMA_signal_1977 ), .Q ( new_AGEMA_signal_10285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C ( clk ), .D ( new_AGEMA_signal_1978 ), .Q ( new_AGEMA_signal_10287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C ( clk ), .D ( new_AGEMA_signal_1979 ), .Q ( new_AGEMA_signal_10289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C ( clk ), .D ( new_AGEMA_signal_10292 ), .Q ( new_AGEMA_signal_10293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C ( clk ), .D ( new_AGEMA_signal_10296 ), .Q ( new_AGEMA_signal_10297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C ( clk ), .D ( new_AGEMA_signal_10300 ), .Q ( new_AGEMA_signal_10301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C ( clk ), .D ( new_AGEMA_signal_10304 ), .Q ( new_AGEMA_signal_10305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C ( clk ), .D ( n2820 ), .Q ( new_AGEMA_signal_10307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C ( clk ), .D ( new_AGEMA_signal_1494 ), .Q ( new_AGEMA_signal_10309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C ( clk ), .D ( new_AGEMA_signal_1495 ), .Q ( new_AGEMA_signal_10311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C ( clk ), .D ( new_AGEMA_signal_1496 ), .Q ( new_AGEMA_signal_10313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C ( clk ), .D ( new_AGEMA_signal_9548 ), .Q ( new_AGEMA_signal_10315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C ( clk ), .D ( new_AGEMA_signal_9550 ), .Q ( new_AGEMA_signal_10319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C ( clk ), .D ( new_AGEMA_signal_9552 ), .Q ( new_AGEMA_signal_10323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C ( clk ), .D ( new_AGEMA_signal_9554 ), .Q ( new_AGEMA_signal_10327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C ( clk ), .D ( n1930 ), .Q ( new_AGEMA_signal_10331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C ( clk ), .D ( new_AGEMA_signal_1224 ), .Q ( new_AGEMA_signal_10335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C ( clk ), .D ( new_AGEMA_signal_1225 ), .Q ( new_AGEMA_signal_10339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C ( clk ), .D ( new_AGEMA_signal_1226 ), .Q ( new_AGEMA_signal_10343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C ( clk ), .D ( n1976 ), .Q ( new_AGEMA_signal_10363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C ( clk ), .D ( new_AGEMA_signal_1296 ), .Q ( new_AGEMA_signal_10367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C ( clk ), .D ( new_AGEMA_signal_1297 ), .Q ( new_AGEMA_signal_10371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C ( clk ), .D ( new_AGEMA_signal_1298 ), .Q ( new_AGEMA_signal_10375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C ( clk ), .D ( new_AGEMA_signal_9212 ), .Q ( new_AGEMA_signal_10387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C ( clk ), .D ( new_AGEMA_signal_9214 ), .Q ( new_AGEMA_signal_10391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C ( clk ), .D ( new_AGEMA_signal_9216 ), .Q ( new_AGEMA_signal_10395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C ( clk ), .D ( new_AGEMA_signal_9218 ), .Q ( new_AGEMA_signal_10399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C ( clk ), .D ( n2008 ), .Q ( new_AGEMA_signal_10411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C ( clk ), .D ( new_AGEMA_signal_1593 ), .Q ( new_AGEMA_signal_10415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C ( clk ), .D ( new_AGEMA_signal_1594 ), .Q ( new_AGEMA_signal_10419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C ( clk ), .D ( new_AGEMA_signal_1595 ), .Q ( new_AGEMA_signal_10423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C ( clk ), .D ( n2022 ), .Q ( new_AGEMA_signal_10427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C ( clk ), .D ( new_AGEMA_signal_1608 ), .Q ( new_AGEMA_signal_10431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C ( clk ), .D ( new_AGEMA_signal_1609 ), .Q ( new_AGEMA_signal_10435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C ( clk ), .D ( new_AGEMA_signal_1610 ), .Q ( new_AGEMA_signal_10439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C ( clk ), .D ( n2057 ), .Q ( new_AGEMA_signal_10475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C ( clk ), .D ( new_AGEMA_signal_1647 ), .Q ( new_AGEMA_signal_10479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C ( clk ), .D ( new_AGEMA_signal_1648 ), .Q ( new_AGEMA_signal_10483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C ( clk ), .D ( new_AGEMA_signal_1649 ), .Q ( new_AGEMA_signal_10487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C ( clk ), .D ( n2062 ), .Q ( new_AGEMA_signal_10491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C ( clk ), .D ( new_AGEMA_signal_1653 ), .Q ( new_AGEMA_signal_10495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C ( clk ), .D ( new_AGEMA_signal_1654 ), .Q ( new_AGEMA_signal_10499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C ( clk ), .D ( new_AGEMA_signal_1655 ), .Q ( new_AGEMA_signal_10503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C ( clk ), .D ( n2075 ), .Q ( new_AGEMA_signal_10507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C ( clk ), .D ( new_AGEMA_signal_1341 ), .Q ( new_AGEMA_signal_10511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C ( clk ), .D ( new_AGEMA_signal_1342 ), .Q ( new_AGEMA_signal_10515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C ( clk ), .D ( new_AGEMA_signal_1343 ), .Q ( new_AGEMA_signal_10519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C ( clk ), .D ( n2121 ), .Q ( new_AGEMA_signal_10547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C ( clk ), .D ( new_AGEMA_signal_1689 ), .Q ( new_AGEMA_signal_10551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C ( clk ), .D ( new_AGEMA_signal_1690 ), .Q ( new_AGEMA_signal_10555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C ( clk ), .D ( new_AGEMA_signal_1691 ), .Q ( new_AGEMA_signal_10559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C ( clk ), .D ( new_AGEMA_signal_9172 ), .Q ( new_AGEMA_signal_10571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C ( clk ), .D ( new_AGEMA_signal_9174 ), .Q ( new_AGEMA_signal_10575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C ( clk ), .D ( new_AGEMA_signal_9176 ), .Q ( new_AGEMA_signal_10579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C ( clk ), .D ( new_AGEMA_signal_9178 ), .Q ( new_AGEMA_signal_10583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C ( clk ), .D ( new_AGEMA_signal_10588 ), .Q ( new_AGEMA_signal_10589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C ( clk ), .D ( new_AGEMA_signal_10594 ), .Q ( new_AGEMA_signal_10595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C ( clk ), .D ( new_AGEMA_signal_10600 ), .Q ( new_AGEMA_signal_10601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C ( clk ), .D ( new_AGEMA_signal_10606 ), .Q ( new_AGEMA_signal_10607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C ( clk ), .D ( new_AGEMA_signal_9460 ), .Q ( new_AGEMA_signal_10611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C ( clk ), .D ( new_AGEMA_signal_9462 ), .Q ( new_AGEMA_signal_10615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C ( clk ), .D ( new_AGEMA_signal_9464 ), .Q ( new_AGEMA_signal_10619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C ( clk ), .D ( new_AGEMA_signal_9466 ), .Q ( new_AGEMA_signal_10623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C ( clk ), .D ( new_AGEMA_signal_9516 ), .Q ( new_AGEMA_signal_10627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C ( clk ), .D ( new_AGEMA_signal_9518 ), .Q ( new_AGEMA_signal_10631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C ( clk ), .D ( new_AGEMA_signal_9520 ), .Q ( new_AGEMA_signal_10635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C ( clk ), .D ( new_AGEMA_signal_9522 ), .Q ( new_AGEMA_signal_10639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C ( clk ), .D ( n2245 ), .Q ( new_AGEMA_signal_10675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C ( clk ), .D ( new_AGEMA_signal_1776 ), .Q ( new_AGEMA_signal_10679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C ( clk ), .D ( new_AGEMA_signal_1777 ), .Q ( new_AGEMA_signal_10683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C ( clk ), .D ( new_AGEMA_signal_1778 ), .Q ( new_AGEMA_signal_10687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C ( clk ), .D ( new_AGEMA_signal_10692 ), .Q ( new_AGEMA_signal_10693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C ( clk ), .D ( new_AGEMA_signal_10698 ), .Q ( new_AGEMA_signal_10699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C ( clk ), .D ( new_AGEMA_signal_10704 ), .Q ( new_AGEMA_signal_10705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C ( clk ), .D ( new_AGEMA_signal_10710 ), .Q ( new_AGEMA_signal_10711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C ( clk ), .D ( n2262 ), .Q ( new_AGEMA_signal_10715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C ( clk ), .D ( new_AGEMA_signal_1389 ), .Q ( new_AGEMA_signal_10719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C ( clk ), .D ( new_AGEMA_signal_1390 ), .Q ( new_AGEMA_signal_10723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C ( clk ), .D ( new_AGEMA_signal_1391 ), .Q ( new_AGEMA_signal_10727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C ( clk ), .D ( n2343 ), .Q ( new_AGEMA_signal_10755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C ( clk ), .D ( new_AGEMA_signal_1827 ), .Q ( new_AGEMA_signal_10759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C ( clk ), .D ( new_AGEMA_signal_1828 ), .Q ( new_AGEMA_signal_10763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C ( clk ), .D ( new_AGEMA_signal_1829 ), .Q ( new_AGEMA_signal_10767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C ( clk ), .D ( new_AGEMA_signal_9468 ), .Q ( new_AGEMA_signal_10787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C ( clk ), .D ( new_AGEMA_signal_9470 ), .Q ( new_AGEMA_signal_10791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C ( clk ), .D ( new_AGEMA_signal_9472 ), .Q ( new_AGEMA_signal_10795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C ( clk ), .D ( new_AGEMA_signal_9474 ), .Q ( new_AGEMA_signal_10799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C ( clk ), .D ( new_AGEMA_signal_9436 ), .Q ( new_AGEMA_signal_10803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C ( clk ), .D ( new_AGEMA_signal_9438 ), .Q ( new_AGEMA_signal_10807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C ( clk ), .D ( new_AGEMA_signal_9440 ), .Q ( new_AGEMA_signal_10811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C ( clk ), .D ( new_AGEMA_signal_9442 ), .Q ( new_AGEMA_signal_10815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C ( clk ), .D ( new_AGEMA_signal_9156 ), .Q ( new_AGEMA_signal_10819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C ( clk ), .D ( new_AGEMA_signal_9158 ), .Q ( new_AGEMA_signal_10823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C ( clk ), .D ( new_AGEMA_signal_9160 ), .Q ( new_AGEMA_signal_10827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C ( clk ), .D ( new_AGEMA_signal_9162 ), .Q ( new_AGEMA_signal_10831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C ( clk ), .D ( new_AGEMA_signal_9260 ), .Q ( new_AGEMA_signal_10835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C ( clk ), .D ( new_AGEMA_signal_9262 ), .Q ( new_AGEMA_signal_10839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C ( clk ), .D ( new_AGEMA_signal_9264 ), .Q ( new_AGEMA_signal_10843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C ( clk ), .D ( new_AGEMA_signal_9266 ), .Q ( new_AGEMA_signal_10847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C ( clk ), .D ( n2417 ), .Q ( new_AGEMA_signal_10851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C ( clk ), .D ( new_AGEMA_signal_2088 ), .Q ( new_AGEMA_signal_10855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C ( clk ), .D ( new_AGEMA_signal_2089 ), .Q ( new_AGEMA_signal_10859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C ( clk ), .D ( new_AGEMA_signal_2090 ), .Q ( new_AGEMA_signal_10863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C ( clk ), .D ( new_AGEMA_signal_9540 ), .Q ( new_AGEMA_signal_10899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C ( clk ), .D ( new_AGEMA_signal_9542 ), .Q ( new_AGEMA_signal_10903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C ( clk ), .D ( new_AGEMA_signal_9544 ), .Q ( new_AGEMA_signal_10907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C ( clk ), .D ( new_AGEMA_signal_9546 ), .Q ( new_AGEMA_signal_10911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C ( clk ), .D ( n2483 ), .Q ( new_AGEMA_signal_10915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C ( clk ), .D ( new_AGEMA_signal_1437 ), .Q ( new_AGEMA_signal_10919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C ( clk ), .D ( new_AGEMA_signal_1438 ), .Q ( new_AGEMA_signal_10923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C ( clk ), .D ( new_AGEMA_signal_1439 ), .Q ( new_AGEMA_signal_10927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2975 ( .C ( clk ), .D ( n2629 ), .Q ( new_AGEMA_signal_11003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2979 ( .C ( clk ), .D ( new_AGEMA_signal_1476 ), .Q ( new_AGEMA_signal_11007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2983 ( .C ( clk ), .D ( new_AGEMA_signal_1477 ), .Q ( new_AGEMA_signal_11011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2987 ( .C ( clk ), .D ( new_AGEMA_signal_1478 ), .Q ( new_AGEMA_signal_11015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3031 ( .C ( clk ), .D ( n2736 ), .Q ( new_AGEMA_signal_11059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3035 ( .C ( clk ), .D ( new_AGEMA_signal_1269 ), .Q ( new_AGEMA_signal_11063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3039 ( .C ( clk ), .D ( new_AGEMA_signal_1270 ), .Q ( new_AGEMA_signal_11067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3043 ( .C ( clk ), .D ( new_AGEMA_signal_1271 ), .Q ( new_AGEMA_signal_11071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3047 ( .C ( clk ), .D ( new_AGEMA_signal_9364 ), .Q ( new_AGEMA_signal_11075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3051 ( .C ( clk ), .D ( new_AGEMA_signal_9366 ), .Q ( new_AGEMA_signal_11079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3055 ( .C ( clk ), .D ( new_AGEMA_signal_9368 ), .Q ( new_AGEMA_signal_11083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3059 ( .C ( clk ), .D ( new_AGEMA_signal_9370 ), .Q ( new_AGEMA_signal_11087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3063 ( .C ( clk ), .D ( new_AGEMA_signal_9252 ), .Q ( new_AGEMA_signal_11091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3067 ( .C ( clk ), .D ( new_AGEMA_signal_9254 ), .Q ( new_AGEMA_signal_11095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3071 ( .C ( clk ), .D ( new_AGEMA_signal_9256 ), .Q ( new_AGEMA_signal_11099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3075 ( .C ( clk ), .D ( new_AGEMA_signal_9258 ), .Q ( new_AGEMA_signal_11103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3079 ( .C ( clk ), .D ( n2787 ), .Q ( new_AGEMA_signal_11107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3083 ( .C ( clk ), .D ( new_AGEMA_signal_2025 ), .Q ( new_AGEMA_signal_11111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3087 ( .C ( clk ), .D ( new_AGEMA_signal_2026 ), .Q ( new_AGEMA_signal_11115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3091 ( .C ( clk ), .D ( new_AGEMA_signal_2027 ), .Q ( new_AGEMA_signal_11119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3129 ( .C ( clk ), .D ( new_AGEMA_signal_11156 ), .Q ( new_AGEMA_signal_11157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3137 ( .C ( clk ), .D ( new_AGEMA_signal_11164 ), .Q ( new_AGEMA_signal_11165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3145 ( .C ( clk ), .D ( new_AGEMA_signal_11172 ), .Q ( new_AGEMA_signal_11173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3153 ( .C ( clk ), .D ( new_AGEMA_signal_11180 ), .Q ( new_AGEMA_signal_11181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3169 ( .C ( clk ), .D ( new_AGEMA_signal_11196 ), .Q ( new_AGEMA_signal_11197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3177 ( .C ( clk ), .D ( new_AGEMA_signal_11204 ), .Q ( new_AGEMA_signal_11205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3185 ( .C ( clk ), .D ( new_AGEMA_signal_11212 ), .Q ( new_AGEMA_signal_11213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3193 ( .C ( clk ), .D ( new_AGEMA_signal_11220 ), .Q ( new_AGEMA_signal_11221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3199 ( .C ( clk ), .D ( n2009 ), .Q ( new_AGEMA_signal_11227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3205 ( .C ( clk ), .D ( new_AGEMA_signal_1602 ), .Q ( new_AGEMA_signal_11233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3211 ( .C ( clk ), .D ( new_AGEMA_signal_1603 ), .Q ( new_AGEMA_signal_11239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3217 ( .C ( clk ), .D ( new_AGEMA_signal_1604 ), .Q ( new_AGEMA_signal_11245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3239 ( .C ( clk ), .D ( n2034 ), .Q ( new_AGEMA_signal_11267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3245 ( .C ( clk ), .D ( new_AGEMA_signal_1332 ), .Q ( new_AGEMA_signal_11273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3251 ( .C ( clk ), .D ( new_AGEMA_signal_1333 ), .Q ( new_AGEMA_signal_11279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3257 ( .C ( clk ), .D ( new_AGEMA_signal_1334 ), .Q ( new_AGEMA_signal_11285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3271 ( .C ( clk ), .D ( new_AGEMA_signal_9532 ), .Q ( new_AGEMA_signal_11299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3277 ( .C ( clk ), .D ( new_AGEMA_signal_9534 ), .Q ( new_AGEMA_signal_11305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3283 ( .C ( clk ), .D ( new_AGEMA_signal_9536 ), .Q ( new_AGEMA_signal_11311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3289 ( .C ( clk ), .D ( new_AGEMA_signal_9538 ), .Q ( new_AGEMA_signal_11317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3295 ( .C ( clk ), .D ( new_AGEMA_signal_9588 ), .Q ( new_AGEMA_signal_11323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3301 ( .C ( clk ), .D ( new_AGEMA_signal_9590 ), .Q ( new_AGEMA_signal_11329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3307 ( .C ( clk ), .D ( new_AGEMA_signal_9592 ), .Q ( new_AGEMA_signal_11335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3313 ( .C ( clk ), .D ( new_AGEMA_signal_9594 ), .Q ( new_AGEMA_signal_11341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3343 ( .C ( clk ), .D ( new_AGEMA_signal_9084 ), .Q ( new_AGEMA_signal_11371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3349 ( .C ( clk ), .D ( new_AGEMA_signal_9086 ), .Q ( new_AGEMA_signal_11377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3355 ( .C ( clk ), .D ( new_AGEMA_signal_9088 ), .Q ( new_AGEMA_signal_11383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3361 ( .C ( clk ), .D ( new_AGEMA_signal_9090 ), .Q ( new_AGEMA_signal_11389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3367 ( .C ( clk ), .D ( n2122 ), .Q ( new_AGEMA_signal_11395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3373 ( .C ( clk ), .D ( new_AGEMA_signal_1695 ), .Q ( new_AGEMA_signal_11401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3379 ( .C ( clk ), .D ( new_AGEMA_signal_1696 ), .Q ( new_AGEMA_signal_11407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3385 ( .C ( clk ), .D ( new_AGEMA_signal_1697 ), .Q ( new_AGEMA_signal_11413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3399 ( .C ( clk ), .D ( n2220 ), .Q ( new_AGEMA_signal_11427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3405 ( .C ( clk ), .D ( new_AGEMA_signal_1713 ), .Q ( new_AGEMA_signal_11433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3411 ( .C ( clk ), .D ( new_AGEMA_signal_1714 ), .Q ( new_AGEMA_signal_11439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3417 ( .C ( clk ), .D ( new_AGEMA_signal_1715 ), .Q ( new_AGEMA_signal_11445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3473 ( .C ( clk ), .D ( new_AGEMA_signal_11500 ), .Q ( new_AGEMA_signal_11501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3481 ( .C ( clk ), .D ( new_AGEMA_signal_11508 ), .Q ( new_AGEMA_signal_11509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3489 ( .C ( clk ), .D ( new_AGEMA_signal_11516 ), .Q ( new_AGEMA_signal_11517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3497 ( .C ( clk ), .D ( new_AGEMA_signal_11524 ), .Q ( new_AGEMA_signal_11525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3503 ( .C ( clk ), .D ( new_AGEMA_signal_9284 ), .Q ( new_AGEMA_signal_11531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3509 ( .C ( clk ), .D ( new_AGEMA_signal_9286 ), .Q ( new_AGEMA_signal_11537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3515 ( .C ( clk ), .D ( new_AGEMA_signal_9288 ), .Q ( new_AGEMA_signal_11543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3521 ( .C ( clk ), .D ( new_AGEMA_signal_9290 ), .Q ( new_AGEMA_signal_11549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3615 ( .C ( clk ), .D ( n2344 ), .Q ( new_AGEMA_signal_11643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3621 ( .C ( clk ), .D ( new_AGEMA_signal_1833 ), .Q ( new_AGEMA_signal_11649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3627 ( .C ( clk ), .D ( new_AGEMA_signal_1834 ), .Q ( new_AGEMA_signal_11655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3633 ( .C ( clk ), .D ( new_AGEMA_signal_1835 ), .Q ( new_AGEMA_signal_11661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3743 ( .C ( clk ), .D ( n2468 ), .Q ( new_AGEMA_signal_11771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3749 ( .C ( clk ), .D ( new_AGEMA_signal_1446 ), .Q ( new_AGEMA_signal_11777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3755 ( .C ( clk ), .D ( new_AGEMA_signal_1447 ), .Q ( new_AGEMA_signal_11783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3761 ( .C ( clk ), .D ( new_AGEMA_signal_1448 ), .Q ( new_AGEMA_signal_11789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3767 ( .C ( clk ), .D ( n2761 ), .Q ( new_AGEMA_signal_11795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3773 ( .C ( clk ), .D ( new_AGEMA_signal_1548 ), .Q ( new_AGEMA_signal_11801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3779 ( .C ( clk ), .D ( new_AGEMA_signal_1549 ), .Q ( new_AGEMA_signal_11807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3785 ( .C ( clk ), .D ( new_AGEMA_signal_1550 ), .Q ( new_AGEMA_signal_11813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3817 ( .C ( clk ), .D ( new_AGEMA_signal_11844 ), .Q ( new_AGEMA_signal_11845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3825 ( .C ( clk ), .D ( new_AGEMA_signal_11852 ), .Q ( new_AGEMA_signal_11853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3833 ( .C ( clk ), .D ( new_AGEMA_signal_11860 ), .Q ( new_AGEMA_signal_11861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3841 ( .C ( clk ), .D ( new_AGEMA_signal_11868 ), .Q ( new_AGEMA_signal_11869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3937 ( .C ( clk ), .D ( new_AGEMA_signal_11964 ), .Q ( new_AGEMA_signal_11965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3945 ( .C ( clk ), .D ( new_AGEMA_signal_11972 ), .Q ( new_AGEMA_signal_11973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3953 ( .C ( clk ), .D ( new_AGEMA_signal_11980 ), .Q ( new_AGEMA_signal_11981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3961 ( .C ( clk ), .D ( new_AGEMA_signal_11988 ), .Q ( new_AGEMA_signal_11989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3999 ( .C ( clk ), .D ( n2825 ), .Q ( new_AGEMA_signal_12027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4005 ( .C ( clk ), .D ( new_AGEMA_signal_2040 ), .Q ( new_AGEMA_signal_12033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4011 ( .C ( clk ), .D ( new_AGEMA_signal_2041 ), .Q ( new_AGEMA_signal_12039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4017 ( .C ( clk ), .D ( new_AGEMA_signal_2042 ), .Q ( new_AGEMA_signal_12045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4031 ( .C ( clk ), .D ( n1957 ), .Q ( new_AGEMA_signal_12059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4039 ( .C ( clk ), .D ( new_AGEMA_signal_1263 ), .Q ( new_AGEMA_signal_12067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4047 ( .C ( clk ), .D ( new_AGEMA_signal_1264 ), .Q ( new_AGEMA_signal_12075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4055 ( .C ( clk ), .D ( new_AGEMA_signal_1265 ), .Q ( new_AGEMA_signal_12083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4087 ( .C ( clk ), .D ( n2026 ), .Q ( new_AGEMA_signal_12115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4095 ( .C ( clk ), .D ( new_AGEMA_signal_1323 ), .Q ( new_AGEMA_signal_12123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4103 ( .C ( clk ), .D ( new_AGEMA_signal_1324 ), .Q ( new_AGEMA_signal_12131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4111 ( .C ( clk ), .D ( new_AGEMA_signal_1325 ), .Q ( new_AGEMA_signal_12139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4167 ( .C ( clk ), .D ( n2811 ), .Q ( new_AGEMA_signal_12195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4175 ( .C ( clk ), .D ( new_AGEMA_signal_1698 ), .Q ( new_AGEMA_signal_12203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4183 ( .C ( clk ), .D ( new_AGEMA_signal_1699 ), .Q ( new_AGEMA_signal_12211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4191 ( .C ( clk ), .D ( new_AGEMA_signal_1700 ), .Q ( new_AGEMA_signal_12219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4351 ( .C ( clk ), .D ( new_AGEMA_signal_9612 ), .Q ( new_AGEMA_signal_12379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4359 ( .C ( clk ), .D ( new_AGEMA_signal_9614 ), .Q ( new_AGEMA_signal_12387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4367 ( .C ( clk ), .D ( new_AGEMA_signal_9616 ), .Q ( new_AGEMA_signal_12395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4375 ( .C ( clk ), .D ( new_AGEMA_signal_9618 ), .Q ( new_AGEMA_signal_12403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4423 ( .C ( clk ), .D ( n2363 ), .Q ( new_AGEMA_signal_12451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4431 ( .C ( clk ), .D ( new_AGEMA_signal_1422 ), .Q ( new_AGEMA_signal_12459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4439 ( .C ( clk ), .D ( new_AGEMA_signal_1423 ), .Q ( new_AGEMA_signal_12467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4447 ( .C ( clk ), .D ( new_AGEMA_signal_1424 ), .Q ( new_AGEMA_signal_12475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4551 ( .C ( clk ), .D ( new_AGEMA_signal_9524 ), .Q ( new_AGEMA_signal_12579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4559 ( .C ( clk ), .D ( new_AGEMA_signal_9526 ), .Q ( new_AGEMA_signal_12587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4567 ( .C ( clk ), .D ( new_AGEMA_signal_9528 ), .Q ( new_AGEMA_signal_12595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4575 ( .C ( clk ), .D ( new_AGEMA_signal_9530 ), .Q ( new_AGEMA_signal_12603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4583 ( .C ( clk ), .D ( new_AGEMA_signal_9124 ), .Q ( new_AGEMA_signal_12611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4591 ( .C ( clk ), .D ( new_AGEMA_signal_9126 ), .Q ( new_AGEMA_signal_12619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4599 ( .C ( clk ), .D ( new_AGEMA_signal_9128 ), .Q ( new_AGEMA_signal_12627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4607 ( .C ( clk ), .D ( new_AGEMA_signal_9130 ), .Q ( new_AGEMA_signal_12635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4927 ( .C ( clk ), .D ( n2544 ), .Q ( new_AGEMA_signal_12955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4937 ( .C ( clk ), .D ( new_AGEMA_signal_1353 ), .Q ( new_AGEMA_signal_12965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4947 ( .C ( clk ), .D ( new_AGEMA_signal_1354 ), .Q ( new_AGEMA_signal_12975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4957 ( .C ( clk ), .D ( new_AGEMA_signal_1355 ), .Q ( new_AGEMA_signal_12985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5127 ( .C ( clk ), .D ( n2364 ), .Q ( new_AGEMA_signal_13155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5137 ( .C ( clk ), .D ( new_AGEMA_signal_1851 ), .Q ( new_AGEMA_signal_13165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5147 ( .C ( clk ), .D ( new_AGEMA_signal_1852 ), .Q ( new_AGEMA_signal_13175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5157 ( .C ( clk ), .D ( new_AGEMA_signal_1853 ), .Q ( new_AGEMA_signal_13185 ) ) ;

    /* cells in depth 6 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1960 ( .a ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}), .b ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}), .clk ( clk ), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, n1924}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1967 ( .a ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, n1922}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9080, new_AGEMA_signal_9078, new_AGEMA_signal_9076}), .clk ( clk ), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n1923}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1981 ( .a ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, n1926}), .b ({new_AGEMA_signal_1511, new_AGEMA_signal_1510, new_AGEMA_signal_1509, n1925}), .clk ( clk ), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, n1927}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1993 ( .a ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .b ({new_AGEMA_signal_1520, new_AGEMA_signal_1519, new_AGEMA_signal_1518, n2763}), .clk ( clk ), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, n1929}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2007 ( .a ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2011 ( .a ({new_AGEMA_signal_9098, new_AGEMA_signal_9096, new_AGEMA_signal_9094, new_AGEMA_signal_9092}), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, n1937}), .clk ( clk ), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n1938}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2019 ( .a ({new_AGEMA_signal_9106, new_AGEMA_signal_9104, new_AGEMA_signal_9102, new_AGEMA_signal_9100}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2023 ( .a ({new_AGEMA_signal_9114, new_AGEMA_signal_9112, new_AGEMA_signal_9110, new_AGEMA_signal_9108}), .b ({new_AGEMA_signal_1244, new_AGEMA_signal_1243, new_AGEMA_signal_1242, n1942}), .clk ( clk ), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, n1943}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2027 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}), .b ({new_AGEMA_signal_9122, new_AGEMA_signal_9120, new_AGEMA_signal_9118, new_AGEMA_signal_9116}), .clk ( clk ), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n1946}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2031 ( .a ({new_AGEMA_signal_9130, new_AGEMA_signal_9128, new_AGEMA_signal_9126, new_AGEMA_signal_9124}), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, n1944}), .clk ( clk ), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, new_AGEMA_signal_2064, n1945}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2034 ( .a ({new_AGEMA_signal_9138, new_AGEMA_signal_9136, new_AGEMA_signal_9134, new_AGEMA_signal_9132}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .clk ( clk ), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, n1956}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2040 ( .a ({new_AGEMA_signal_1538, new_AGEMA_signal_1537, new_AGEMA_signal_1536, n1950}), .b ({new_AGEMA_signal_1256, new_AGEMA_signal_1255, new_AGEMA_signal_1254, n1949}), .clk ( clk ), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n1951}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2048 ( .a ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .b ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, n1952}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2057 ( .a ({new_AGEMA_signal_9146, new_AGEMA_signal_9144, new_AGEMA_signal_9142, new_AGEMA_signal_9140}), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}), .clk ( clk ), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(1)) U2061 ( .a ({new_AGEMA_signal_1502, new_AGEMA_signal_1501, new_AGEMA_signal_1500, n1962}), .b ({new_AGEMA_signal_9154, new_AGEMA_signal_9152, new_AGEMA_signal_9150, new_AGEMA_signal_9148}), .clk ( clk ), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, n1966}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2064 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9160, new_AGEMA_signal_9158, new_AGEMA_signal_9156}), .clk ( clk ), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, new_AGEMA_signal_1545, n1963}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2077 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, n1968}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2082 ( .a ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .b ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2088 ( .a ({new_AGEMA_signal_9170, new_AGEMA_signal_9168, new_AGEMA_signal_9166, new_AGEMA_signal_9164}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n1972}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2092 ( .a ({new_AGEMA_signal_9178, new_AGEMA_signal_9176, new_AGEMA_signal_9174, new_AGEMA_signal_9172}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}), .clk ( clk ), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, n1971}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2099 ( .a ({new_AGEMA_signal_9186, new_AGEMA_signal_9184, new_AGEMA_signal_9182, new_AGEMA_signal_9180}), .b ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, n2535}), .clk ( clk ), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, n1974}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2106 ( .a ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .b ({new_AGEMA_signal_9146, new_AGEMA_signal_9144, new_AGEMA_signal_9142, new_AGEMA_signal_9140}), .clk ( clk ), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, new_AGEMA_signal_2100, n1979}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2112 ( .a ({new_AGEMA_signal_9194, new_AGEMA_signal_9192, new_AGEMA_signal_9190, new_AGEMA_signal_9188}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, new_AGEMA_signal_1572, n1985}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2121 ( .a ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, n1992}), .b ({new_AGEMA_signal_1583, new_AGEMA_signal_1582, new_AGEMA_signal_1581, n1991}), .clk ( clk ), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n1994}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2126 ( .a ({new_AGEMA_signal_9202, new_AGEMA_signal_9200, new_AGEMA_signal_9198, new_AGEMA_signal_9196}), .b ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, n1995}), .clk ( clk ), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, n1996}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2136 ( .a ({new_AGEMA_signal_9210, new_AGEMA_signal_9208, new_AGEMA_signal_9206, new_AGEMA_signal_9204}), .b ({new_AGEMA_signal_1592, new_AGEMA_signal_1591, new_AGEMA_signal_1590, n2003}), .clk ( clk ), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2142 ( .a ({new_AGEMA_signal_9218, new_AGEMA_signal_9216, new_AGEMA_signal_9214, new_AGEMA_signal_9212}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .clk ( clk ), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, n2006}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2144 ( .a ({new_AGEMA_signal_9226, new_AGEMA_signal_9224, new_AGEMA_signal_9222, new_AGEMA_signal_9220}), .b ({new_AGEMA_signal_1601, new_AGEMA_signal_1600, new_AGEMA_signal_1599, n2004}), .clk ( clk ), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2005}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2152 ( .a ({new_AGEMA_signal_9234, new_AGEMA_signal_9232, new_AGEMA_signal_9230, new_AGEMA_signal_9228}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, n2013}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2160 ( .a ({new_AGEMA_signal_9242, new_AGEMA_signal_9240, new_AGEMA_signal_9238, new_AGEMA_signal_9236}), .b ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}), .clk ( clk ), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, n2020}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2164 ( .a ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .b ({new_AGEMA_signal_9250, new_AGEMA_signal_9248, new_AGEMA_signal_9246, new_AGEMA_signal_9244}), .clk ( clk ), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, n2023}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2168 ( .a ({new_AGEMA_signal_1145, new_AGEMA_signal_1144, new_AGEMA_signal_1143, n2027}), .b ({new_AGEMA_signal_9258, new_AGEMA_signal_9256, new_AGEMA_signal_9254, new_AGEMA_signal_9252}), .clk ( clk ), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, n2028}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2172 ( .a ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, n2033}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2175 ( .a ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .b ({new_AGEMA_signal_9274, new_AGEMA_signal_9272, new_AGEMA_signal_9270, new_AGEMA_signal_9268}), .clk ( clk ), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2031}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2184 ( .a ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .b ({new_AGEMA_signal_1628, new_AGEMA_signal_1627, new_AGEMA_signal_1626, n2039}), .clk ( clk ), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, n2040}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2187 ( .a ({new_AGEMA_signal_9282, new_AGEMA_signal_9280, new_AGEMA_signal_9278, new_AGEMA_signal_9276}), .b ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, n2050}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2193 ( .a ({new_AGEMA_signal_9290, new_AGEMA_signal_9288, new_AGEMA_signal_9286, new_AGEMA_signal_9284}), .b ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, n2044}), .clk ( clk ), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2045}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2199 ( .a ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .b ({new_AGEMA_signal_9146, new_AGEMA_signal_9144, new_AGEMA_signal_9142, new_AGEMA_signal_9140}), .clk ( clk ), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, n2051}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2203 ( .a ({new_AGEMA_signal_9298, new_AGEMA_signal_9296, new_AGEMA_signal_9294, new_AGEMA_signal_9292}), .b ({new_AGEMA_signal_1646, new_AGEMA_signal_1645, new_AGEMA_signal_1644, n2055}), .clk ( clk ), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2056}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2209 ( .a ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9304, new_AGEMA_signal_9302, new_AGEMA_signal_9300}), .clk ( clk ), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, n2060}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2215 ( .a ({new_AGEMA_signal_9314, new_AGEMA_signal_9312, new_AGEMA_signal_9310, new_AGEMA_signal_9308}), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .clk ( clk ), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2066}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2217 ( .a ({new_AGEMA_signal_9258, new_AGEMA_signal_9256, new_AGEMA_signal_9254, new_AGEMA_signal_9252}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, n2065}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2221 ( .a ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, n2068}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_2156, new_AGEMA_signal_2155, new_AGEMA_signal_2154, n2069}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2226 ( .a ({new_AGEMA_signal_9322, new_AGEMA_signal_9320, new_AGEMA_signal_9318, new_AGEMA_signal_9316}), .b ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}), .clk ( clk ), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, n2074}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2235 ( .a ({new_AGEMA_signal_1346, new_AGEMA_signal_1345, new_AGEMA_signal_1344, n2081}), .b ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, n2080}), .clk ( clk ), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2082}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2240 ( .a ({new_AGEMA_signal_9226, new_AGEMA_signal_9224, new_AGEMA_signal_9222, new_AGEMA_signal_9220}), .b ({new_AGEMA_signal_1673, new_AGEMA_signal_1672, new_AGEMA_signal_1671, n2083}), .clk ( clk ), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, n2084}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2242 ( .a ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .b ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .clk ( clk ), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2085}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2245 ( .a ({new_AGEMA_signal_9330, new_AGEMA_signal_9328, new_AGEMA_signal_9326, new_AGEMA_signal_9324}), .b ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}), .clk ( clk ), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2248 ( .a ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, n2088}), .b ({new_AGEMA_signal_1352, new_AGEMA_signal_1351, new_AGEMA_signal_1350, n2087}), .clk ( clk ), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_2174, new_AGEMA_signal_2173, new_AGEMA_signal_2172, n2089}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2252 ( .a ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}), .clk ( clk ), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2254 ( .a ({new_AGEMA_signal_9338, new_AGEMA_signal_9336, new_AGEMA_signal_9334, new_AGEMA_signal_9332}), .b ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .clk ( clk ), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, n2092}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(1)) U2256 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .b ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .clk ( clk ), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, n2094}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2261 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, n2101}), .b ({new_AGEMA_signal_1682, new_AGEMA_signal_1681, new_AGEMA_signal_1680, n2100}), .clk ( clk ), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2265 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2271 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .b ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2114}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2273 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .b ({new_AGEMA_signal_9226, new_AGEMA_signal_9224, new_AGEMA_signal_9222, new_AGEMA_signal_9220}), .clk ( clk ), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, n2115}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2280 ( .a ({new_AGEMA_signal_9346, new_AGEMA_signal_9344, new_AGEMA_signal_9342, new_AGEMA_signal_9340}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2281 ( .a ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, n2119}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2291 ( .a ({new_AGEMA_signal_9354, new_AGEMA_signal_9352, new_AGEMA_signal_9350, new_AGEMA_signal_9348}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, n2130}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2292 ( .a ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .b ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .clk ( clk ), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2129}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2295 ( .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .b ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .clk ( clk ), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_1709, new_AGEMA_signal_1708, new_AGEMA_signal_1707, n2150}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2298 ( .a ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .b ({new_AGEMA_signal_1364, new_AGEMA_signal_1363, new_AGEMA_signal_1362, n2132}), .clk ( clk ), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2133}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2302 ( .a ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .b ({new_AGEMA_signal_9370, new_AGEMA_signal_9368, new_AGEMA_signal_9366, new_AGEMA_signal_9364}), .clk ( clk ), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, n2136}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2306 ( .a ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .b ({new_AGEMA_signal_1718, new_AGEMA_signal_1717, new_AGEMA_signal_1716, n2138}), .clk ( clk ), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2139}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2313 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9376, new_AGEMA_signal_9374, new_AGEMA_signal_9372}), .b ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}), .clk ( clk ), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, n2144}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2318 ( .a ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, n2151}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_2210, new_AGEMA_signal_2209, new_AGEMA_signal_2208, n2152}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2321 ( .a ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, n2156}), .clk ( clk ), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, n2170}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2323 ( .a ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2157}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2329 ( .a ({new_AGEMA_signal_9386, new_AGEMA_signal_9384, new_AGEMA_signal_9382, new_AGEMA_signal_9380}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, n2162}), .clk ( clk ), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, new_AGEMA_signal_1725, n2163}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2335 ( .a ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, n2171}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, n2172}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2338 ( .a ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .b ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}), .clk ( clk ), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_1370, new_AGEMA_signal_1369, new_AGEMA_signal_1368, n2186}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2339 ( .a ({new_AGEMA_signal_9186, new_AGEMA_signal_9184, new_AGEMA_signal_9182, new_AGEMA_signal_9180}), .b ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .clk ( clk ), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, n2181}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2344 ( .a ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, n2176}), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, n2175}), .clk ( clk ), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2177}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2349 ( .a ({new_AGEMA_signal_9146, new_AGEMA_signal_9144, new_AGEMA_signal_9142, new_AGEMA_signal_9140}), .b ({new_AGEMA_signal_1166, new_AGEMA_signal_1165, new_AGEMA_signal_1164, n2182}), .clk ( clk ), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_1376, new_AGEMA_signal_1375, new_AGEMA_signal_1374, n2183}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2354 ( .a ({new_AGEMA_signal_9394, new_AGEMA_signal_9392, new_AGEMA_signal_9390, new_AGEMA_signal_9388}), .b ({new_AGEMA_signal_1736, new_AGEMA_signal_1735, new_AGEMA_signal_1734, n2188}), .clk ( clk ), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, n2195}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2356 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, n2190}), .b ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, n2189}), .clk ( clk ), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, n2193}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2358 ( .a ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}), .clk ( clk ), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, n2191}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2364 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .b ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}), .clk ( clk ), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_1745, new_AGEMA_signal_1744, new_AGEMA_signal_1743, n2196}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2367 ( .a ({new_AGEMA_signal_9122, new_AGEMA_signal_9120, new_AGEMA_signal_9118, new_AGEMA_signal_9116}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .clk ( clk ), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2201}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2369 ( .a ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .b ({new_AGEMA_signal_9410, new_AGEMA_signal_9408, new_AGEMA_signal_9406, new_AGEMA_signal_9404}), .clk ( clk ), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, n2200}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2371 ( .s ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .clk ( clk ), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, n2202}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2379 ( .a ({new_AGEMA_signal_1619, new_AGEMA_signal_1618, new_AGEMA_signal_1617, n2214}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, n2213}), .clk ( clk ), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, new_AGEMA_signal_2244, n2217}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2381 ( .a ({new_AGEMA_signal_9418, new_AGEMA_signal_9416, new_AGEMA_signal_9414, new_AGEMA_signal_9412}), .b ({new_AGEMA_signal_1388, new_AGEMA_signal_1387, new_AGEMA_signal_1386, n2215}), .clk ( clk ), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2216}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2385 ( .a ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, n2218}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .clk ( clk ), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, n2222}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2387 ( .a ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, n2220}), .b ({new_AGEMA_signal_1754, new_AGEMA_signal_1753, new_AGEMA_signal_1752, n2219}), .clk ( clk ), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2221}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2391 ( .a ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .b ({new_AGEMA_signal_9426, new_AGEMA_signal_9424, new_AGEMA_signal_9422, new_AGEMA_signal_9420}), .clk ( clk ), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, n2226}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2393 ( .s ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .b ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .a ({new_AGEMA_signal_1328, new_AGEMA_signal_1327, new_AGEMA_signal_1326, n2227}), .clk ( clk ), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, n2228}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2397 ( .a ({new_AGEMA_signal_9242, new_AGEMA_signal_9240, new_AGEMA_signal_9238, new_AGEMA_signal_9236}), .b ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_1763, new_AGEMA_signal_1762, new_AGEMA_signal_1761, n2237}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2398 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .b ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .clk ( clk ), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2233}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2403 ( .a ({new_AGEMA_signal_9434, new_AGEMA_signal_9432, new_AGEMA_signal_9430, new_AGEMA_signal_9428}), .b ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .clk ( clk ), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, n2238}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2406 ( .a ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, n2241}), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, n2240}), .clk ( clk ), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, n2248}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2409 ( .a ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}), .b ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, n2243}), .clk ( clk ), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, n2244}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2414 ( .a ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9080, new_AGEMA_signal_9078, new_AGEMA_signal_9076}), .clk ( clk ), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_2264, new_AGEMA_signal_2263, new_AGEMA_signal_2262, n2249}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2417 ( .s ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .b ({new_AGEMA_signal_1664, new_AGEMA_signal_1663, new_AGEMA_signal_1662, n2252}), .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, n2253}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2424 ( .a ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .b ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, n2259}), .clk ( clk ), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2260}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2429 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .b ({new_AGEMA_signal_9442, new_AGEMA_signal_9440, new_AGEMA_signal_9438, new_AGEMA_signal_9436}), .clk ( clk ), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, n2273}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2430 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9448, new_AGEMA_signal_9446, new_AGEMA_signal_9444}), .b ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .clk ( clk ), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, n2752}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2433 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}), .b ({new_AGEMA_signal_9346, new_AGEMA_signal_9344, new_AGEMA_signal_9342, new_AGEMA_signal_9340}), .clk ( clk ), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, n2265}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2437 ( .a ({new_AGEMA_signal_9458, new_AGEMA_signal_9456, new_AGEMA_signal_9454, new_AGEMA_signal_9452}), .b ({new_AGEMA_signal_1400, new_AGEMA_signal_1399, new_AGEMA_signal_1398, n2268}), .clk ( clk ), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2269}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2444 ( .a ({new_AGEMA_signal_9162, new_AGEMA_signal_9160, new_AGEMA_signal_9158, new_AGEMA_signal_9156}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2277}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2449 ( .a ({new_AGEMA_signal_9466, new_AGEMA_signal_9464, new_AGEMA_signal_9462, new_AGEMA_signal_9460}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}), .clk ( clk ), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, new_AGEMA_signal_1797, n2282}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2452 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, n2284}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2456 ( .a ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .b ({new_AGEMA_signal_9474, new_AGEMA_signal_9472, new_AGEMA_signal_9470, new_AGEMA_signal_9468}), .clk ( clk ), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2459 ( .a ({new_AGEMA_signal_9098, new_AGEMA_signal_9096, new_AGEMA_signal_9094, new_AGEMA_signal_9092}), .b ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, n2287}), .clk ( clk ), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, n2288}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2462 ( .a ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .b ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .clk ( clk ), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2464 ( .a ({new_AGEMA_signal_9386, new_AGEMA_signal_9384, new_AGEMA_signal_9382, new_AGEMA_signal_9380}), .b ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, n2290}), .clk ( clk ), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, n2293}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2467 ( .a ({new_AGEMA_signal_9338, new_AGEMA_signal_9336, new_AGEMA_signal_9334, new_AGEMA_signal_9332}), .b ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .clk ( clk ), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_1808, new_AGEMA_signal_1807, new_AGEMA_signal_1806, n2294}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2472 ( .a ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .b ({new_AGEMA_signal_1406, new_AGEMA_signal_1405, new_AGEMA_signal_1404, n2299}), .clk ( clk ), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2300}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2480 ( .a ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, n2734}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .clk ( clk ), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, n2323}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) U2482 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .b ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}), .clk ( clk ), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2314}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2485 ( .a ({new_AGEMA_signal_1172, new_AGEMA_signal_1171, new_AGEMA_signal_1170, n2316}), .b ({new_AGEMA_signal_9482, new_AGEMA_signal_9480, new_AGEMA_signal_9478, new_AGEMA_signal_9476}), .clk ( clk ), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, n2319}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2491 ( .a ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .clk ( clk ), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2326}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2496 ( .a ({new_AGEMA_signal_1826, new_AGEMA_signal_1825, new_AGEMA_signal_1824, n2328}), .b ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, n2327}), .clk ( clk ), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2329}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2501 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, n2417}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, n2335}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2506 ( .a ({new_AGEMA_signal_9234, new_AGEMA_signal_9232, new_AGEMA_signal_9230, new_AGEMA_signal_9228}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, n2341}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2507 ( .a ({new_AGEMA_signal_9490, new_AGEMA_signal_9488, new_AGEMA_signal_9486, new_AGEMA_signal_9484}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .clk ( clk ), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2340}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2514 ( .a ({new_AGEMA_signal_1418, new_AGEMA_signal_1417, new_AGEMA_signal_1416, n2348}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, n2347}), .clk ( clk ), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, n2349}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2517 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9496, new_AGEMA_signal_9494, new_AGEMA_signal_9492}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .clk ( clk ), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, n2375}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2518 ( .a ({new_AGEMA_signal_9378, new_AGEMA_signal_9376, new_AGEMA_signal_9374, new_AGEMA_signal_9372}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, n2736}), .clk ( clk ), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2352}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2522 ( .a ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, n2353}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, n2354}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2525 ( .a ({new_AGEMA_signal_9506, new_AGEMA_signal_9504, new_AGEMA_signal_9502, new_AGEMA_signal_9500}), .b ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, n2355}), .clk ( clk ), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, n2357}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2527 ( .a ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, n2359}), .b ({new_AGEMA_signal_9514, new_AGEMA_signal_9512, new_AGEMA_signal_9510, new_AGEMA_signal_9508}), .clk ( clk ), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, n2360}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2534 ( .a ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, n2369}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2536 ( .a ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, n2371}), .b ({new_AGEMA_signal_9426, new_AGEMA_signal_9424, new_AGEMA_signal_9422, new_AGEMA_signal_9420}), .clk ( clk ), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, n2372}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2539 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, n2376}), .clk ( clk ), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, n2377}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2544 ( .a ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .b ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}), .clk ( clk ), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, n2467}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2545 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9520, new_AGEMA_signal_9518, new_AGEMA_signal_9516}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, n2383}), .clk ( clk ), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, n2385}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2546 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2384}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2548 ( .a ({new_AGEMA_signal_9226, new_AGEMA_signal_9224, new_AGEMA_signal_9222, new_AGEMA_signal_9220}), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .clk ( clk ), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, n2386}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2552 ( .a ({new_AGEMA_signal_9394, new_AGEMA_signal_9392, new_AGEMA_signal_9390, new_AGEMA_signal_9388}), .b ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .clk ( clk ), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, n2394}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2553 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .clk ( clk ), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2391}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2554 ( .a ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2390}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2559 ( .a ({new_AGEMA_signal_9338, new_AGEMA_signal_9336, new_AGEMA_signal_9334, new_AGEMA_signal_9332}), .b ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .clk ( clk ), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_1871, new_AGEMA_signal_1870, new_AGEMA_signal_1869, n2396}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2562 ( .a ({new_AGEMA_signal_9530, new_AGEMA_signal_9528, new_AGEMA_signal_9526, new_AGEMA_signal_9524}), .b ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .clk ( clk ), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, n2406}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2565 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}), .b ({new_AGEMA_signal_1436, new_AGEMA_signal_1435, new_AGEMA_signal_1434, n2402}), .clk ( clk ), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2403}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2569 ( .a ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, n2407}), .b ({new_AGEMA_signal_9370, new_AGEMA_signal_9368, new_AGEMA_signal_9366, new_AGEMA_signal_9364}), .clk ( clk ), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, n2408}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2573 ( .a ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, n2412}), .b ({new_AGEMA_signal_9434, new_AGEMA_signal_9432, new_AGEMA_signal_9430, new_AGEMA_signal_9428}), .clk ( clk ), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2574 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .b ({new_AGEMA_signal_9290, new_AGEMA_signal_9288, new_AGEMA_signal_9286, new_AGEMA_signal_9284}), .clk ( clk ), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, n2413}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2577 ( .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, n2415}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2416}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2586 ( .a ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, n2428}), .b ({new_AGEMA_signal_9538, new_AGEMA_signal_9536, new_AGEMA_signal_9534, new_AGEMA_signal_9532}), .clk ( clk ), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, n2433}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2587 ( .a ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, n2429}), .clk ( clk ), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2591 ( .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, n2647}), .b ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .clk ( clk ), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, n2434}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2595 ( .a ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, n2438}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, n2483}), .clk ( clk ), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, n2439}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2598 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9520, new_AGEMA_signal_9518, new_AGEMA_signal_9516}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .clk ( clk ), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2445}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2600 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .b ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, n2443}), .clk ( clk ), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, n2444}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2602 ( .a ({new_AGEMA_signal_9186, new_AGEMA_signal_9184, new_AGEMA_signal_9182, new_AGEMA_signal_9180}), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, n2446}), .clk ( clk ), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2447}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2607 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}), .clk ( clk ), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, n2454}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2617 ( .a ({new_AGEMA_signal_9346, new_AGEMA_signal_9344, new_AGEMA_signal_9342, new_AGEMA_signal_9340}), .b ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, n2464}), .clk ( clk ), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2465}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2622 ( .a ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .b ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .clk ( clk ), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, n2470}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2626 ( .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, n2473}), .b ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, n2472}), .clk ( clk ), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2476}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2633 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9544, new_AGEMA_signal_9542, new_AGEMA_signal_9540}), .b ({new_AGEMA_signal_1907, new_AGEMA_signal_1906, new_AGEMA_signal_1905, n2480}), .clk ( clk ), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2481}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2639 ( .a ({new_AGEMA_signal_9554, new_AGEMA_signal_9552, new_AGEMA_signal_9550, new_AGEMA_signal_9548}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, n2486}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2642 ( .a ({new_AGEMA_signal_9450, new_AGEMA_signal_9448, new_AGEMA_signal_9446, new_AGEMA_signal_9444}), .b ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, n2488}), .clk ( clk ), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_1916, new_AGEMA_signal_1915, new_AGEMA_signal_1914, n2489}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2645 ( .a ({new_AGEMA_signal_9562, new_AGEMA_signal_9560, new_AGEMA_signal_9558, new_AGEMA_signal_9556}), .b ({new_AGEMA_signal_1232, new_AGEMA_signal_1231, new_AGEMA_signal_1230, n2492}), .clk ( clk ), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, n2497}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2646 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9568, new_AGEMA_signal_9566, new_AGEMA_signal_9564}), .b ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .clk ( clk ), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2495}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2647 ( .a ({new_AGEMA_signal_9354, new_AGEMA_signal_9352, new_AGEMA_signal_9350, new_AGEMA_signal_9348}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2494}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2650 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, n2498}), .b ({new_AGEMA_signal_9122, new_AGEMA_signal_9120, new_AGEMA_signal_9118, new_AGEMA_signal_9116}), .clk ( clk ), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_1925, new_AGEMA_signal_1924, new_AGEMA_signal_1923, n2499}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2653 ( .a ({new_AGEMA_signal_9122, new_AGEMA_signal_9120, new_AGEMA_signal_9118, new_AGEMA_signal_9116}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, n2674}), .clk ( clk ), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, n2503}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2655 ( .s ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .b ({new_AGEMA_signal_1556, new_AGEMA_signal_1555, new_AGEMA_signal_1554, n2505}), .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .clk ( clk ), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, n2506}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2662 ( .a ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .b ({new_AGEMA_signal_9210, new_AGEMA_signal_9208, new_AGEMA_signal_9206, new_AGEMA_signal_9204}), .clk ( clk ), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, n2518}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2663 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2517}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2666 ( .a ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, n2520}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .clk ( clk ), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, n2523}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2668 ( .a ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, n2521}), .clk ( clk ), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2522}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2675 ( .a ({new_AGEMA_signal_9210, new_AGEMA_signal_9208, new_AGEMA_signal_9206, new_AGEMA_signal_9204}), .b ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, n2531}), .clk ( clk ), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, n2532}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2677 ( .a ({new_AGEMA_signal_9082, new_AGEMA_signal_9080, new_AGEMA_signal_9078, new_AGEMA_signal_9076}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, n2533}), .clk ( clk ), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2534}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2681 ( .a ({new_AGEMA_signal_9578, new_AGEMA_signal_9576, new_AGEMA_signal_9574, new_AGEMA_signal_9572}), .b ({new_AGEMA_signal_1781, new_AGEMA_signal_1780, new_AGEMA_signal_1779, n2540}), .clk ( clk ), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, n2542}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2683 ( .a ({new_AGEMA_signal_1160, new_AGEMA_signal_1159, new_AGEMA_signal_1158, n2545}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, n2544}), .clk ( clk ), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2546}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2687 ( .a ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .clk ( clk ), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, n2551}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2690 ( .a ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, n2553}), .b ({new_AGEMA_signal_9586, new_AGEMA_signal_9584, new_AGEMA_signal_9582, new_AGEMA_signal_9580}), .clk ( clk ), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, n2558}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2692 ( .a ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, n2555}), .b ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, n2554}), .clk ( clk ), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, n2556}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2696 ( .a ({new_AGEMA_signal_1772, new_AGEMA_signal_1771, new_AGEMA_signal_1770, n2561}), .b ({new_AGEMA_signal_1466, new_AGEMA_signal_1465, new_AGEMA_signal_1464, n2560}), .clk ( clk ), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, n2566}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2697 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9592, new_AGEMA_signal_9590, new_AGEMA_signal_9588}), .b ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, n2562}), .clk ( clk ), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2703 ( .a ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, n2572}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, n2571}), .clk ( clk ), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2573}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2705 ( .a ({new_AGEMA_signal_9530, new_AGEMA_signal_9528, new_AGEMA_signal_9526, new_AGEMA_signal_9524}), .b ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .clk ( clk ), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, n2585}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2706 ( .a ({new_AGEMA_signal_9442, new_AGEMA_signal_9440, new_AGEMA_signal_9438, new_AGEMA_signal_9436}), .b ({new_AGEMA_signal_1262, new_AGEMA_signal_1261, new_AGEMA_signal_1260, n2627}), .clk ( clk ), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, n2581}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2707 ( .a ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, n2575}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2579}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2708 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9568, new_AGEMA_signal_9566, new_AGEMA_signal_9564}), .b ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, n2576}), .clk ( clk ), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, n2578}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2711 ( .a ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .b ({new_AGEMA_signal_9410, new_AGEMA_signal_9408, new_AGEMA_signal_9406, new_AGEMA_signal_9404}), .clk ( clk ), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, n2582}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2715 ( .a ({new_AGEMA_signal_9154, new_AGEMA_signal_9152, new_AGEMA_signal_9150, new_AGEMA_signal_9148}), .b ({new_AGEMA_signal_1952, new_AGEMA_signal_1951, new_AGEMA_signal_1950, n2586}), .clk ( clk ), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, n2588}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2719 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, n2594}), .b ({new_AGEMA_signal_9530, new_AGEMA_signal_9528, new_AGEMA_signal_9526, new_AGEMA_signal_9524}), .clk ( clk ), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, n2607}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2722 ( .a ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, n2597}), .b ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, n2596}), .clk ( clk ), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, n2605}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2724 ( .a ({new_AGEMA_signal_1961, new_AGEMA_signal_1960, new_AGEMA_signal_1959, n2598}), .b ({new_AGEMA_signal_9602, new_AGEMA_signal_9600, new_AGEMA_signal_9598, new_AGEMA_signal_9596}), .clk ( clk ), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, n2603}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2726 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, n2599}), .b ({new_AGEMA_signal_9434, new_AGEMA_signal_9432, new_AGEMA_signal_9430, new_AGEMA_signal_9428}), .clk ( clk ), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2601}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2733 ( .a ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, n2610}), .b ({new_AGEMA_signal_9402, new_AGEMA_signal_9400, new_AGEMA_signal_9398, new_AGEMA_signal_9396}), .clk ( clk ), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, n2620}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2736 ( .a ({new_AGEMA_signal_1970, new_AGEMA_signal_1969, new_AGEMA_signal_1968, n2614}), .b ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, n2613}), .clk ( clk ), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2618}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2743 ( .a ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, n2625}), .clk ( clk ), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, n2626}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2746 ( .a ({new_AGEMA_signal_1220, new_AGEMA_signal_1219, new_AGEMA_signal_1218, n2631}), .b ({new_AGEMA_signal_9266, new_AGEMA_signal_9264, new_AGEMA_signal_9262, new_AGEMA_signal_9260}), .clk ( clk ), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, n2632}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2752 ( .a ({new_AGEMA_signal_1979, new_AGEMA_signal_1978, new_AGEMA_signal_1977, n2784}), .b ({new_AGEMA_signal_1340, new_AGEMA_signal_1339, new_AGEMA_signal_1338, n2642}), .clk ( clk ), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2644}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2754 ( .a ({new_AGEMA_signal_9114, new_AGEMA_signal_9112, new_AGEMA_signal_9110, new_AGEMA_signal_9108}), .b ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, n2645}), .clk ( clk ), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2646}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2758 ( .a ({new_AGEMA_signal_1286, new_AGEMA_signal_1285, new_AGEMA_signal_1284, n2651}), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, n2650}), .clk ( clk ), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, n2653}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2760 ( .a ({new_AGEMA_signal_9434, new_AGEMA_signal_9432, new_AGEMA_signal_9430, new_AGEMA_signal_9428}), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, n2654}), .clk ( clk ), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, n2655}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2764 ( .a ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, n2662}), .b ({new_AGEMA_signal_9450, new_AGEMA_signal_9448, new_AGEMA_signal_9446, new_AGEMA_signal_9444}), .clk ( clk ), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, n2663}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2770 ( .a ({new_AGEMA_signal_1274, new_AGEMA_signal_1273, new_AGEMA_signal_1272, n2673}), .b ({new_AGEMA_signal_9410, new_AGEMA_signal_9408, new_AGEMA_signal_9406, new_AGEMA_signal_9404}), .clk ( clk ), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2675}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2772 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, n2677}), .b ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, n2676}), .clk ( clk ), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, n2678}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2780 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, n2690}), .b ({new_AGEMA_signal_9442, new_AGEMA_signal_9440, new_AGEMA_signal_9438, new_AGEMA_signal_9436}), .clk ( clk ), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, n2691}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2782 ( .a ({new_AGEMA_signal_9466, new_AGEMA_signal_9464, new_AGEMA_signal_9462, new_AGEMA_signal_9460}), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, n2693}), .clk ( clk ), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, n2695}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2785 ( .a ({new_AGEMA_signal_1430, new_AGEMA_signal_1429, new_AGEMA_signal_1428, n2700}), .b ({new_AGEMA_signal_9594, new_AGEMA_signal_9592, new_AGEMA_signal_9590, new_AGEMA_signal_9588}), .clk ( clk ), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, new_AGEMA_signal_1995, n2701}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2791 ( .a ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, n2711}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, n2710}), .clk ( clk ), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, n2717}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2796 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, n2720}), .b ({new_AGEMA_signal_9362, new_AGEMA_signal_9360, new_AGEMA_signal_9358, new_AGEMA_signal_9356}), .clk ( clk ), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, n2729}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2798 ( .a ({new_AGEMA_signal_9226, new_AGEMA_signal_9224, new_AGEMA_signal_9222, new_AGEMA_signal_9220}), .b ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, n2722}), .clk ( clk ), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, new_AGEMA_signal_2004, n2727}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2803 ( .a ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, n2732}), .b ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, n2731}), .clk ( clk ), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2733}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2807 ( .a ({new_AGEMA_signal_9610, new_AGEMA_signal_9608, new_AGEMA_signal_9606, new_AGEMA_signal_9604}), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, n2738}), .clk ( clk ), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, n2740}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2812 ( .a ({new_AGEMA_signal_1382, new_AGEMA_signal_1381, new_AGEMA_signal_1380, n2748}), .b ({new_AGEMA_signal_9082, new_AGEMA_signal_9080, new_AGEMA_signal_9078, new_AGEMA_signal_9076}), .clk ( clk ), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, new_AGEMA_signal_2013, n2749}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2815 ( .a ({new_AGEMA_signal_1637, new_AGEMA_signal_1636, new_AGEMA_signal_1635, n2754}), .b ({new_AGEMA_signal_9242, new_AGEMA_signal_9240, new_AGEMA_signal_9238, new_AGEMA_signal_9236}), .clk ( clk ), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, n2757}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2816 ( .a ({new_AGEMA_signal_1208, new_AGEMA_signal_1207, new_AGEMA_signal_1206, n2755}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9616, new_AGEMA_signal_9614, new_AGEMA_signal_9612}), .clk ( clk ), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, n2756}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2819 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, n2761}), .b ({new_AGEMA_signal_9474, new_AGEMA_signal_9472, new_AGEMA_signal_9470, new_AGEMA_signal_9468}), .clk ( clk ), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2762}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2823 ( .a ({new_AGEMA_signal_9082, new_AGEMA_signal_9080, new_AGEMA_signal_9078, new_AGEMA_signal_9076}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, n2768}), .clk ( clk ), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, n2770}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2825 ( .a ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, n2773}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9616, new_AGEMA_signal_9614, new_AGEMA_signal_9612}), .clk ( clk ), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2776}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2826 ( .a ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, n2774}), .b ({new_AGEMA_signal_9090, new_AGEMA_signal_9088, new_AGEMA_signal_9086, new_AGEMA_signal_9084}), .clk ( clk ), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, n2775}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2830 ( .a ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, n2782}), .b ({new_AGEMA_signal_1493, new_AGEMA_signal_1492, new_AGEMA_signal_1491, n2781}), .clk ( clk ), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2783}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2836 ( .a ({new_AGEMA_signal_2030, new_AGEMA_signal_2029, new_AGEMA_signal_2028, n2794}), .b ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, n2793}), .clk ( clk ), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, n2795}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2845 ( .a ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, n2812}), .b ({new_AGEMA_signal_1700, new_AGEMA_signal_1699, new_AGEMA_signal_1698, n2811}), .clk ( clk ), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2814}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2848 ( .a ({new_AGEMA_signal_9178, new_AGEMA_signal_9176, new_AGEMA_signal_9174, new_AGEMA_signal_9172}), .b ({new_AGEMA_signal_1304, new_AGEMA_signal_1303, new_AGEMA_signal_1302, n2817}), .clk ( clk ), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, n2819}) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C ( clk ), .D ( new_AGEMA_signal_9619 ), .Q ( new_AGEMA_signal_9620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C ( clk ), .D ( new_AGEMA_signal_9621 ), .Q ( new_AGEMA_signal_9622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C ( clk ), .D ( new_AGEMA_signal_9623 ), .Q ( new_AGEMA_signal_9624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C ( clk ), .D ( new_AGEMA_signal_9625 ), .Q ( new_AGEMA_signal_9626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C ( clk ), .D ( new_AGEMA_signal_9627 ), .Q ( new_AGEMA_signal_9628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C ( clk ), .D ( new_AGEMA_signal_9629 ), .Q ( new_AGEMA_signal_9630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C ( clk ), .D ( new_AGEMA_signal_9631 ), .Q ( new_AGEMA_signal_9632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C ( clk ), .D ( new_AGEMA_signal_9633 ), .Q ( new_AGEMA_signal_9634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C ( clk ), .D ( new_AGEMA_signal_9637 ), .Q ( new_AGEMA_signal_9638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C ( clk ), .D ( new_AGEMA_signal_9641 ), .Q ( new_AGEMA_signal_9642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C ( clk ), .D ( new_AGEMA_signal_9645 ), .Q ( new_AGEMA_signal_9646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C ( clk ), .D ( new_AGEMA_signal_9649 ), .Q ( new_AGEMA_signal_9650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C ( clk ), .D ( new_AGEMA_signal_9651 ), .Q ( new_AGEMA_signal_9652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C ( clk ), .D ( new_AGEMA_signal_9653 ), .Q ( new_AGEMA_signal_9654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C ( clk ), .D ( new_AGEMA_signal_9655 ), .Q ( new_AGEMA_signal_9656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C ( clk ), .D ( new_AGEMA_signal_9657 ), .Q ( new_AGEMA_signal_9658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C ( clk ), .D ( new_AGEMA_signal_9659 ), .Q ( new_AGEMA_signal_9660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C ( clk ), .D ( new_AGEMA_signal_9661 ), .Q ( new_AGEMA_signal_9662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C ( clk ), .D ( new_AGEMA_signal_9663 ), .Q ( new_AGEMA_signal_9664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C ( clk ), .D ( new_AGEMA_signal_9665 ), .Q ( new_AGEMA_signal_9666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C ( clk ), .D ( new_AGEMA_signal_9667 ), .Q ( new_AGEMA_signal_9668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C ( clk ), .D ( new_AGEMA_signal_9669 ), .Q ( new_AGEMA_signal_9670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C ( clk ), .D ( new_AGEMA_signal_9671 ), .Q ( new_AGEMA_signal_9672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C ( clk ), .D ( new_AGEMA_signal_9673 ), .Q ( new_AGEMA_signal_9674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C ( clk ), .D ( new_AGEMA_signal_9675 ), .Q ( new_AGEMA_signal_9676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C ( clk ), .D ( new_AGEMA_signal_9677 ), .Q ( new_AGEMA_signal_9678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C ( clk ), .D ( new_AGEMA_signal_9679 ), .Q ( new_AGEMA_signal_9680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C ( clk ), .D ( new_AGEMA_signal_9681 ), .Q ( new_AGEMA_signal_9682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C ( clk ), .D ( new_AGEMA_signal_9683 ), .Q ( new_AGEMA_signal_9684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C ( clk ), .D ( new_AGEMA_signal_9685 ), .Q ( new_AGEMA_signal_9686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C ( clk ), .D ( new_AGEMA_signal_9687 ), .Q ( new_AGEMA_signal_9688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C ( clk ), .D ( new_AGEMA_signal_9689 ), .Q ( new_AGEMA_signal_9690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C ( clk ), .D ( new_AGEMA_signal_9691 ), .Q ( new_AGEMA_signal_9692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C ( clk ), .D ( new_AGEMA_signal_9693 ), .Q ( new_AGEMA_signal_9694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C ( clk ), .D ( new_AGEMA_signal_9695 ), .Q ( new_AGEMA_signal_9696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C ( clk ), .D ( new_AGEMA_signal_9697 ), .Q ( new_AGEMA_signal_9698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C ( clk ), .D ( new_AGEMA_signal_9699 ), .Q ( new_AGEMA_signal_9700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C ( clk ), .D ( new_AGEMA_signal_9701 ), .Q ( new_AGEMA_signal_9702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C ( clk ), .D ( new_AGEMA_signal_9703 ), .Q ( new_AGEMA_signal_9704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C ( clk ), .D ( new_AGEMA_signal_9705 ), .Q ( new_AGEMA_signal_9706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C ( clk ), .D ( new_AGEMA_signal_9707 ), .Q ( new_AGEMA_signal_9708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C ( clk ), .D ( new_AGEMA_signal_9709 ), .Q ( new_AGEMA_signal_9710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C ( clk ), .D ( new_AGEMA_signal_9711 ), .Q ( new_AGEMA_signal_9712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C ( clk ), .D ( new_AGEMA_signal_9713 ), .Q ( new_AGEMA_signal_9714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C ( clk ), .D ( new_AGEMA_signal_9715 ), .Q ( new_AGEMA_signal_9716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C ( clk ), .D ( new_AGEMA_signal_9717 ), .Q ( new_AGEMA_signal_9718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C ( clk ), .D ( new_AGEMA_signal_9719 ), .Q ( new_AGEMA_signal_9720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C ( clk ), .D ( new_AGEMA_signal_9721 ), .Q ( new_AGEMA_signal_9722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C ( clk ), .D ( new_AGEMA_signal_9723 ), .Q ( new_AGEMA_signal_9724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C ( clk ), .D ( new_AGEMA_signal_9725 ), .Q ( new_AGEMA_signal_9726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C ( clk ), .D ( new_AGEMA_signal_9727 ), .Q ( new_AGEMA_signal_9728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C ( clk ), .D ( new_AGEMA_signal_9729 ), .Q ( new_AGEMA_signal_9730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C ( clk ), .D ( new_AGEMA_signal_9731 ), .Q ( new_AGEMA_signal_9732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C ( clk ), .D ( new_AGEMA_signal_9733 ), .Q ( new_AGEMA_signal_9734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C ( clk ), .D ( new_AGEMA_signal_9735 ), .Q ( new_AGEMA_signal_9736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C ( clk ), .D ( new_AGEMA_signal_9737 ), .Q ( new_AGEMA_signal_9738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C ( clk ), .D ( new_AGEMA_signal_9741 ), .Q ( new_AGEMA_signal_9742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C ( clk ), .D ( new_AGEMA_signal_9745 ), .Q ( new_AGEMA_signal_9746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C ( clk ), .D ( new_AGEMA_signal_9749 ), .Q ( new_AGEMA_signal_9750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C ( clk ), .D ( new_AGEMA_signal_9753 ), .Q ( new_AGEMA_signal_9754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C ( clk ), .D ( new_AGEMA_signal_9755 ), .Q ( new_AGEMA_signal_9756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C ( clk ), .D ( new_AGEMA_signal_9757 ), .Q ( new_AGEMA_signal_9758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C ( clk ), .D ( new_AGEMA_signal_9759 ), .Q ( new_AGEMA_signal_9760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C ( clk ), .D ( new_AGEMA_signal_9761 ), .Q ( new_AGEMA_signal_9762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C ( clk ), .D ( new_AGEMA_signal_9763 ), .Q ( new_AGEMA_signal_9764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C ( clk ), .D ( new_AGEMA_signal_9765 ), .Q ( new_AGEMA_signal_9766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C ( clk ), .D ( new_AGEMA_signal_9767 ), .Q ( new_AGEMA_signal_9768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C ( clk ), .D ( new_AGEMA_signal_9769 ), .Q ( new_AGEMA_signal_9770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C ( clk ), .D ( new_AGEMA_signal_9771 ), .Q ( new_AGEMA_signal_9772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C ( clk ), .D ( new_AGEMA_signal_9773 ), .Q ( new_AGEMA_signal_9774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C ( clk ), .D ( new_AGEMA_signal_9775 ), .Q ( new_AGEMA_signal_9776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C ( clk ), .D ( new_AGEMA_signal_9777 ), .Q ( new_AGEMA_signal_9778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C ( clk ), .D ( new_AGEMA_signal_9779 ), .Q ( new_AGEMA_signal_9780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C ( clk ), .D ( new_AGEMA_signal_9781 ), .Q ( new_AGEMA_signal_9782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C ( clk ), .D ( new_AGEMA_signal_9783 ), .Q ( new_AGEMA_signal_9784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C ( clk ), .D ( new_AGEMA_signal_9785 ), .Q ( new_AGEMA_signal_9786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C ( clk ), .D ( new_AGEMA_signal_9787 ), .Q ( new_AGEMA_signal_9788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C ( clk ), .D ( new_AGEMA_signal_9789 ), .Q ( new_AGEMA_signal_9790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C ( clk ), .D ( new_AGEMA_signal_9791 ), .Q ( new_AGEMA_signal_9792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C ( clk ), .D ( new_AGEMA_signal_9793 ), .Q ( new_AGEMA_signal_9794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C ( clk ), .D ( new_AGEMA_signal_9795 ), .Q ( new_AGEMA_signal_9796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C ( clk ), .D ( new_AGEMA_signal_9797 ), .Q ( new_AGEMA_signal_9798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C ( clk ), .D ( new_AGEMA_signal_9799 ), .Q ( new_AGEMA_signal_9800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C ( clk ), .D ( new_AGEMA_signal_9801 ), .Q ( new_AGEMA_signal_9802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C ( clk ), .D ( new_AGEMA_signal_9803 ), .Q ( new_AGEMA_signal_9804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C ( clk ), .D ( new_AGEMA_signal_9805 ), .Q ( new_AGEMA_signal_9806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C ( clk ), .D ( new_AGEMA_signal_9807 ), .Q ( new_AGEMA_signal_9808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C ( clk ), .D ( new_AGEMA_signal_9809 ), .Q ( new_AGEMA_signal_9810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C ( clk ), .D ( new_AGEMA_signal_9813 ), .Q ( new_AGEMA_signal_9814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C ( clk ), .D ( new_AGEMA_signal_9817 ), .Q ( new_AGEMA_signal_9818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C ( clk ), .D ( new_AGEMA_signal_9821 ), .Q ( new_AGEMA_signal_9822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C ( clk ), .D ( new_AGEMA_signal_9825 ), .Q ( new_AGEMA_signal_9826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C ( clk ), .D ( new_AGEMA_signal_9827 ), .Q ( new_AGEMA_signal_9828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C ( clk ), .D ( new_AGEMA_signal_9829 ), .Q ( new_AGEMA_signal_9830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C ( clk ), .D ( new_AGEMA_signal_9831 ), .Q ( new_AGEMA_signal_9832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C ( clk ), .D ( new_AGEMA_signal_9833 ), .Q ( new_AGEMA_signal_9834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C ( clk ), .D ( new_AGEMA_signal_9835 ), .Q ( new_AGEMA_signal_9836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C ( clk ), .D ( new_AGEMA_signal_9837 ), .Q ( new_AGEMA_signal_9838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C ( clk ), .D ( new_AGEMA_signal_9839 ), .Q ( new_AGEMA_signal_9840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C ( clk ), .D ( new_AGEMA_signal_9841 ), .Q ( new_AGEMA_signal_9842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C ( clk ), .D ( new_AGEMA_signal_9843 ), .Q ( new_AGEMA_signal_9844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C ( clk ), .D ( new_AGEMA_signal_9845 ), .Q ( new_AGEMA_signal_9846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C ( clk ), .D ( new_AGEMA_signal_9847 ), .Q ( new_AGEMA_signal_9848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C ( clk ), .D ( new_AGEMA_signal_9849 ), .Q ( new_AGEMA_signal_9850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C ( clk ), .D ( new_AGEMA_signal_9851 ), .Q ( new_AGEMA_signal_9852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C ( clk ), .D ( new_AGEMA_signal_9853 ), .Q ( new_AGEMA_signal_9854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C ( clk ), .D ( new_AGEMA_signal_9855 ), .Q ( new_AGEMA_signal_9856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C ( clk ), .D ( new_AGEMA_signal_9857 ), .Q ( new_AGEMA_signal_9858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C ( clk ), .D ( new_AGEMA_signal_9859 ), .Q ( new_AGEMA_signal_9860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C ( clk ), .D ( new_AGEMA_signal_9861 ), .Q ( new_AGEMA_signal_9862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C ( clk ), .D ( new_AGEMA_signal_9863 ), .Q ( new_AGEMA_signal_9864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C ( clk ), .D ( new_AGEMA_signal_9865 ), .Q ( new_AGEMA_signal_9866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C ( clk ), .D ( new_AGEMA_signal_9869 ), .Q ( new_AGEMA_signal_9870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C ( clk ), .D ( new_AGEMA_signal_9873 ), .Q ( new_AGEMA_signal_9874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C ( clk ), .D ( new_AGEMA_signal_9877 ), .Q ( new_AGEMA_signal_9878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C ( clk ), .D ( new_AGEMA_signal_9881 ), .Q ( new_AGEMA_signal_9882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C ( clk ), .D ( new_AGEMA_signal_9883 ), .Q ( new_AGEMA_signal_9884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C ( clk ), .D ( new_AGEMA_signal_9885 ), .Q ( new_AGEMA_signal_9886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C ( clk ), .D ( new_AGEMA_signal_9887 ), .Q ( new_AGEMA_signal_9888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C ( clk ), .D ( new_AGEMA_signal_9889 ), .Q ( new_AGEMA_signal_9890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C ( clk ), .D ( new_AGEMA_signal_9891 ), .Q ( new_AGEMA_signal_9892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C ( clk ), .D ( new_AGEMA_signal_9893 ), .Q ( new_AGEMA_signal_9894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C ( clk ), .D ( new_AGEMA_signal_9895 ), .Q ( new_AGEMA_signal_9896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C ( clk ), .D ( new_AGEMA_signal_9897 ), .Q ( new_AGEMA_signal_9898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C ( clk ), .D ( new_AGEMA_signal_9899 ), .Q ( new_AGEMA_signal_9900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C ( clk ), .D ( new_AGEMA_signal_9901 ), .Q ( new_AGEMA_signal_9902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C ( clk ), .D ( new_AGEMA_signal_9903 ), .Q ( new_AGEMA_signal_9904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C ( clk ), .D ( new_AGEMA_signal_9905 ), .Q ( new_AGEMA_signal_9906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C ( clk ), .D ( new_AGEMA_signal_9909 ), .Q ( new_AGEMA_signal_9910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C ( clk ), .D ( new_AGEMA_signal_9913 ), .Q ( new_AGEMA_signal_9914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C ( clk ), .D ( new_AGEMA_signal_9917 ), .Q ( new_AGEMA_signal_9918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C ( clk ), .D ( new_AGEMA_signal_9921 ), .Q ( new_AGEMA_signal_9922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C ( clk ), .D ( new_AGEMA_signal_9923 ), .Q ( new_AGEMA_signal_9924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C ( clk ), .D ( new_AGEMA_signal_9925 ), .Q ( new_AGEMA_signal_9926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C ( clk ), .D ( new_AGEMA_signal_9927 ), .Q ( new_AGEMA_signal_9928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C ( clk ), .D ( new_AGEMA_signal_9929 ), .Q ( new_AGEMA_signal_9930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C ( clk ), .D ( new_AGEMA_signal_9931 ), .Q ( new_AGEMA_signal_9932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C ( clk ), .D ( new_AGEMA_signal_9933 ), .Q ( new_AGEMA_signal_9934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C ( clk ), .D ( new_AGEMA_signal_9935 ), .Q ( new_AGEMA_signal_9936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C ( clk ), .D ( new_AGEMA_signal_9937 ), .Q ( new_AGEMA_signal_9938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C ( clk ), .D ( new_AGEMA_signal_9939 ), .Q ( new_AGEMA_signal_9940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C ( clk ), .D ( new_AGEMA_signal_9941 ), .Q ( new_AGEMA_signal_9942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C ( clk ), .D ( new_AGEMA_signal_9943 ), .Q ( new_AGEMA_signal_9944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C ( clk ), .D ( new_AGEMA_signal_9945 ), .Q ( new_AGEMA_signal_9946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C ( clk ), .D ( new_AGEMA_signal_9949 ), .Q ( new_AGEMA_signal_9950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C ( clk ), .D ( new_AGEMA_signal_9953 ), .Q ( new_AGEMA_signal_9954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C ( clk ), .D ( new_AGEMA_signal_9957 ), .Q ( new_AGEMA_signal_9958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C ( clk ), .D ( new_AGEMA_signal_9961 ), .Q ( new_AGEMA_signal_9962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C ( clk ), .D ( new_AGEMA_signal_9963 ), .Q ( new_AGEMA_signal_9964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C ( clk ), .D ( new_AGEMA_signal_9965 ), .Q ( new_AGEMA_signal_9966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C ( clk ), .D ( new_AGEMA_signal_9967 ), .Q ( new_AGEMA_signal_9968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C ( clk ), .D ( new_AGEMA_signal_9969 ), .Q ( new_AGEMA_signal_9970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C ( clk ), .D ( new_AGEMA_signal_9971 ), .Q ( new_AGEMA_signal_9972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C ( clk ), .D ( new_AGEMA_signal_9973 ), .Q ( new_AGEMA_signal_9974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C ( clk ), .D ( new_AGEMA_signal_9975 ), .Q ( new_AGEMA_signal_9976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C ( clk ), .D ( new_AGEMA_signal_9977 ), .Q ( new_AGEMA_signal_9978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C ( clk ), .D ( new_AGEMA_signal_9979 ), .Q ( new_AGEMA_signal_9980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C ( clk ), .D ( new_AGEMA_signal_9981 ), .Q ( new_AGEMA_signal_9982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C ( clk ), .D ( new_AGEMA_signal_9983 ), .Q ( new_AGEMA_signal_9984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C ( clk ), .D ( new_AGEMA_signal_9985 ), .Q ( new_AGEMA_signal_9986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C ( clk ), .D ( new_AGEMA_signal_9987 ), .Q ( new_AGEMA_signal_9988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C ( clk ), .D ( new_AGEMA_signal_9989 ), .Q ( new_AGEMA_signal_9990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C ( clk ), .D ( new_AGEMA_signal_9991 ), .Q ( new_AGEMA_signal_9992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C ( clk ), .D ( new_AGEMA_signal_9993 ), .Q ( new_AGEMA_signal_9994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C ( clk ), .D ( new_AGEMA_signal_9995 ), .Q ( new_AGEMA_signal_9996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C ( clk ), .D ( new_AGEMA_signal_9997 ), .Q ( new_AGEMA_signal_9998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C ( clk ), .D ( new_AGEMA_signal_9999 ), .Q ( new_AGEMA_signal_10000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C ( clk ), .D ( new_AGEMA_signal_10001 ), .Q ( new_AGEMA_signal_10002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C ( clk ), .D ( new_AGEMA_signal_10003 ), .Q ( new_AGEMA_signal_10004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C ( clk ), .D ( new_AGEMA_signal_10005 ), .Q ( new_AGEMA_signal_10006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C ( clk ), .D ( new_AGEMA_signal_10007 ), .Q ( new_AGEMA_signal_10008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C ( clk ), .D ( new_AGEMA_signal_10009 ), .Q ( new_AGEMA_signal_10010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C ( clk ), .D ( new_AGEMA_signal_10011 ), .Q ( new_AGEMA_signal_10012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C ( clk ), .D ( new_AGEMA_signal_10013 ), .Q ( new_AGEMA_signal_10014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C ( clk ), .D ( new_AGEMA_signal_10015 ), .Q ( new_AGEMA_signal_10016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C ( clk ), .D ( new_AGEMA_signal_10017 ), .Q ( new_AGEMA_signal_10018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C ( clk ), .D ( new_AGEMA_signal_10019 ), .Q ( new_AGEMA_signal_10020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C ( clk ), .D ( new_AGEMA_signal_10021 ), .Q ( new_AGEMA_signal_10022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C ( clk ), .D ( new_AGEMA_signal_10023 ), .Q ( new_AGEMA_signal_10024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C ( clk ), .D ( new_AGEMA_signal_10025 ), .Q ( new_AGEMA_signal_10026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C ( clk ), .D ( new_AGEMA_signal_10027 ), .Q ( new_AGEMA_signal_10028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C ( clk ), .D ( new_AGEMA_signal_10029 ), .Q ( new_AGEMA_signal_10030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C ( clk ), .D ( new_AGEMA_signal_10031 ), .Q ( new_AGEMA_signal_10032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C ( clk ), .D ( new_AGEMA_signal_10033 ), .Q ( new_AGEMA_signal_10034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C ( clk ), .D ( new_AGEMA_signal_10035 ), .Q ( new_AGEMA_signal_10036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C ( clk ), .D ( new_AGEMA_signal_10037 ), .Q ( new_AGEMA_signal_10038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C ( clk ), .D ( new_AGEMA_signal_10039 ), .Q ( new_AGEMA_signal_10040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C ( clk ), .D ( new_AGEMA_signal_10041 ), .Q ( new_AGEMA_signal_10042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C ( clk ), .D ( new_AGEMA_signal_10043 ), .Q ( new_AGEMA_signal_10044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C ( clk ), .D ( new_AGEMA_signal_10045 ), .Q ( new_AGEMA_signal_10046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C ( clk ), .D ( new_AGEMA_signal_10047 ), .Q ( new_AGEMA_signal_10048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C ( clk ), .D ( new_AGEMA_signal_10049 ), .Q ( new_AGEMA_signal_10050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C ( clk ), .D ( new_AGEMA_signal_10051 ), .Q ( new_AGEMA_signal_10052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C ( clk ), .D ( new_AGEMA_signal_10053 ), .Q ( new_AGEMA_signal_10054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C ( clk ), .D ( new_AGEMA_signal_10055 ), .Q ( new_AGEMA_signal_10056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C ( clk ), .D ( new_AGEMA_signal_10057 ), .Q ( new_AGEMA_signal_10058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C ( clk ), .D ( new_AGEMA_signal_10059 ), .Q ( new_AGEMA_signal_10060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C ( clk ), .D ( new_AGEMA_signal_10061 ), .Q ( new_AGEMA_signal_10062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C ( clk ), .D ( new_AGEMA_signal_10063 ), .Q ( new_AGEMA_signal_10064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C ( clk ), .D ( new_AGEMA_signal_10065 ), .Q ( new_AGEMA_signal_10066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C ( clk ), .D ( new_AGEMA_signal_10067 ), .Q ( new_AGEMA_signal_10068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C ( clk ), .D ( new_AGEMA_signal_10069 ), .Q ( new_AGEMA_signal_10070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C ( clk ), .D ( new_AGEMA_signal_10071 ), .Q ( new_AGEMA_signal_10072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C ( clk ), .D ( new_AGEMA_signal_10073 ), .Q ( new_AGEMA_signal_10074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C ( clk ), .D ( new_AGEMA_signal_10075 ), .Q ( new_AGEMA_signal_10076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C ( clk ), .D ( new_AGEMA_signal_10077 ), .Q ( new_AGEMA_signal_10078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C ( clk ), .D ( new_AGEMA_signal_10079 ), .Q ( new_AGEMA_signal_10080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C ( clk ), .D ( new_AGEMA_signal_10081 ), .Q ( new_AGEMA_signal_10082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C ( clk ), .D ( new_AGEMA_signal_10083 ), .Q ( new_AGEMA_signal_10084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C ( clk ), .D ( new_AGEMA_signal_10085 ), .Q ( new_AGEMA_signal_10086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C ( clk ), .D ( new_AGEMA_signal_10087 ), .Q ( new_AGEMA_signal_10088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C ( clk ), .D ( new_AGEMA_signal_10089 ), .Q ( new_AGEMA_signal_10090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C ( clk ), .D ( new_AGEMA_signal_10091 ), .Q ( new_AGEMA_signal_10092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C ( clk ), .D ( new_AGEMA_signal_10093 ), .Q ( new_AGEMA_signal_10094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C ( clk ), .D ( new_AGEMA_signal_10095 ), .Q ( new_AGEMA_signal_10096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C ( clk ), .D ( new_AGEMA_signal_10097 ), .Q ( new_AGEMA_signal_10098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C ( clk ), .D ( new_AGEMA_signal_10103 ), .Q ( new_AGEMA_signal_10104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C ( clk ), .D ( new_AGEMA_signal_10109 ), .Q ( new_AGEMA_signal_10110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C ( clk ), .D ( new_AGEMA_signal_10115 ), .Q ( new_AGEMA_signal_10116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C ( clk ), .D ( new_AGEMA_signal_10121 ), .Q ( new_AGEMA_signal_10122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C ( clk ), .D ( new_AGEMA_signal_10123 ), .Q ( new_AGEMA_signal_10124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C ( clk ), .D ( new_AGEMA_signal_10125 ), .Q ( new_AGEMA_signal_10126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C ( clk ), .D ( new_AGEMA_signal_10127 ), .Q ( new_AGEMA_signal_10128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C ( clk ), .D ( new_AGEMA_signal_10129 ), .Q ( new_AGEMA_signal_10130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C ( clk ), .D ( new_AGEMA_signal_10131 ), .Q ( new_AGEMA_signal_10132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C ( clk ), .D ( new_AGEMA_signal_10133 ), .Q ( new_AGEMA_signal_10134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C ( clk ), .D ( new_AGEMA_signal_10135 ), .Q ( new_AGEMA_signal_10136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C ( clk ), .D ( new_AGEMA_signal_10137 ), .Q ( new_AGEMA_signal_10138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C ( clk ), .D ( new_AGEMA_signal_10139 ), .Q ( new_AGEMA_signal_10140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C ( clk ), .D ( new_AGEMA_signal_10141 ), .Q ( new_AGEMA_signal_10142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C ( clk ), .D ( new_AGEMA_signal_10143 ), .Q ( new_AGEMA_signal_10144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C ( clk ), .D ( new_AGEMA_signal_10145 ), .Q ( new_AGEMA_signal_10146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C ( clk ), .D ( new_AGEMA_signal_10149 ), .Q ( new_AGEMA_signal_10150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C ( clk ), .D ( new_AGEMA_signal_10153 ), .Q ( new_AGEMA_signal_10154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C ( clk ), .D ( new_AGEMA_signal_10157 ), .Q ( new_AGEMA_signal_10158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C ( clk ), .D ( new_AGEMA_signal_10161 ), .Q ( new_AGEMA_signal_10162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C ( clk ), .D ( new_AGEMA_signal_10163 ), .Q ( new_AGEMA_signal_10164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C ( clk ), .D ( new_AGEMA_signal_10165 ), .Q ( new_AGEMA_signal_10166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C ( clk ), .D ( new_AGEMA_signal_10167 ), .Q ( new_AGEMA_signal_10168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C ( clk ), .D ( new_AGEMA_signal_10169 ), .Q ( new_AGEMA_signal_10170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C ( clk ), .D ( new_AGEMA_signal_10171 ), .Q ( new_AGEMA_signal_10172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C ( clk ), .D ( new_AGEMA_signal_10173 ), .Q ( new_AGEMA_signal_10174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C ( clk ), .D ( new_AGEMA_signal_10175 ), .Q ( new_AGEMA_signal_10176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C ( clk ), .D ( new_AGEMA_signal_10177 ), .Q ( new_AGEMA_signal_10178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C ( clk ), .D ( new_AGEMA_signal_10179 ), .Q ( new_AGEMA_signal_10180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C ( clk ), .D ( new_AGEMA_signal_10181 ), .Q ( new_AGEMA_signal_10182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C ( clk ), .D ( new_AGEMA_signal_10183 ), .Q ( new_AGEMA_signal_10184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C ( clk ), .D ( new_AGEMA_signal_10185 ), .Q ( new_AGEMA_signal_10186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C ( clk ), .D ( new_AGEMA_signal_10189 ), .Q ( new_AGEMA_signal_10190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C ( clk ), .D ( new_AGEMA_signal_10193 ), .Q ( new_AGEMA_signal_10194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C ( clk ), .D ( new_AGEMA_signal_10197 ), .Q ( new_AGEMA_signal_10198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C ( clk ), .D ( new_AGEMA_signal_10201 ), .Q ( new_AGEMA_signal_10202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C ( clk ), .D ( new_AGEMA_signal_10203 ), .Q ( new_AGEMA_signal_10204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C ( clk ), .D ( new_AGEMA_signal_10205 ), .Q ( new_AGEMA_signal_10206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C ( clk ), .D ( new_AGEMA_signal_10207 ), .Q ( new_AGEMA_signal_10208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C ( clk ), .D ( new_AGEMA_signal_10209 ), .Q ( new_AGEMA_signal_10210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C ( clk ), .D ( new_AGEMA_signal_10211 ), .Q ( new_AGEMA_signal_10212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C ( clk ), .D ( new_AGEMA_signal_10213 ), .Q ( new_AGEMA_signal_10214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C ( clk ), .D ( new_AGEMA_signal_10215 ), .Q ( new_AGEMA_signal_10216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C ( clk ), .D ( new_AGEMA_signal_10217 ), .Q ( new_AGEMA_signal_10218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C ( clk ), .D ( new_AGEMA_signal_10219 ), .Q ( new_AGEMA_signal_10220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C ( clk ), .D ( new_AGEMA_signal_10221 ), .Q ( new_AGEMA_signal_10222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C ( clk ), .D ( new_AGEMA_signal_10223 ), .Q ( new_AGEMA_signal_10224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C ( clk ), .D ( new_AGEMA_signal_10225 ), .Q ( new_AGEMA_signal_10226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C ( clk ), .D ( new_AGEMA_signal_10227 ), .Q ( new_AGEMA_signal_10228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C ( clk ), .D ( new_AGEMA_signal_10229 ), .Q ( new_AGEMA_signal_10230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C ( clk ), .D ( new_AGEMA_signal_10231 ), .Q ( new_AGEMA_signal_10232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C ( clk ), .D ( new_AGEMA_signal_10233 ), .Q ( new_AGEMA_signal_10234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C ( clk ), .D ( new_AGEMA_signal_10235 ), .Q ( new_AGEMA_signal_10236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C ( clk ), .D ( new_AGEMA_signal_10237 ), .Q ( new_AGEMA_signal_10238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C ( clk ), .D ( new_AGEMA_signal_10239 ), .Q ( new_AGEMA_signal_10240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C ( clk ), .D ( new_AGEMA_signal_10241 ), .Q ( new_AGEMA_signal_10242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C ( clk ), .D ( new_AGEMA_signal_10243 ), .Q ( new_AGEMA_signal_10244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C ( clk ), .D ( new_AGEMA_signal_10245 ), .Q ( new_AGEMA_signal_10246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C ( clk ), .D ( new_AGEMA_signal_10247 ), .Q ( new_AGEMA_signal_10248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C ( clk ), .D ( new_AGEMA_signal_10249 ), .Q ( new_AGEMA_signal_10250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C ( clk ), .D ( new_AGEMA_signal_10251 ), .Q ( new_AGEMA_signal_10252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C ( clk ), .D ( new_AGEMA_signal_10253 ), .Q ( new_AGEMA_signal_10254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C ( clk ), .D ( new_AGEMA_signal_10255 ), .Q ( new_AGEMA_signal_10256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C ( clk ), .D ( new_AGEMA_signal_10257 ), .Q ( new_AGEMA_signal_10258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C ( clk ), .D ( new_AGEMA_signal_10261 ), .Q ( new_AGEMA_signal_10262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C ( clk ), .D ( new_AGEMA_signal_10265 ), .Q ( new_AGEMA_signal_10266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C ( clk ), .D ( new_AGEMA_signal_10269 ), .Q ( new_AGEMA_signal_10270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C ( clk ), .D ( new_AGEMA_signal_10273 ), .Q ( new_AGEMA_signal_10274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C ( clk ), .D ( new_AGEMA_signal_10275 ), .Q ( new_AGEMA_signal_10276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C ( clk ), .D ( new_AGEMA_signal_10277 ), .Q ( new_AGEMA_signal_10278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C ( clk ), .D ( new_AGEMA_signal_10279 ), .Q ( new_AGEMA_signal_10280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C ( clk ), .D ( new_AGEMA_signal_10281 ), .Q ( new_AGEMA_signal_10282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C ( clk ), .D ( new_AGEMA_signal_10283 ), .Q ( new_AGEMA_signal_10284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C ( clk ), .D ( new_AGEMA_signal_10285 ), .Q ( new_AGEMA_signal_10286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C ( clk ), .D ( new_AGEMA_signal_10287 ), .Q ( new_AGEMA_signal_10288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C ( clk ), .D ( new_AGEMA_signal_10289 ), .Q ( new_AGEMA_signal_10290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C ( clk ), .D ( new_AGEMA_signal_10293 ), .Q ( new_AGEMA_signal_10294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C ( clk ), .D ( new_AGEMA_signal_10297 ), .Q ( new_AGEMA_signal_10298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C ( clk ), .D ( new_AGEMA_signal_10301 ), .Q ( new_AGEMA_signal_10302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C ( clk ), .D ( new_AGEMA_signal_10305 ), .Q ( new_AGEMA_signal_10306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C ( clk ), .D ( new_AGEMA_signal_10307 ), .Q ( new_AGEMA_signal_10308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C ( clk ), .D ( new_AGEMA_signal_10309 ), .Q ( new_AGEMA_signal_10310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C ( clk ), .D ( new_AGEMA_signal_10311 ), .Q ( new_AGEMA_signal_10312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C ( clk ), .D ( new_AGEMA_signal_10313 ), .Q ( new_AGEMA_signal_10314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C ( clk ), .D ( new_AGEMA_signal_10315 ), .Q ( new_AGEMA_signal_10316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C ( clk ), .D ( new_AGEMA_signal_10319 ), .Q ( new_AGEMA_signal_10320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C ( clk ), .D ( new_AGEMA_signal_10323 ), .Q ( new_AGEMA_signal_10324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C ( clk ), .D ( new_AGEMA_signal_10327 ), .Q ( new_AGEMA_signal_10328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C ( clk ), .D ( new_AGEMA_signal_10331 ), .Q ( new_AGEMA_signal_10332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C ( clk ), .D ( new_AGEMA_signal_10335 ), .Q ( new_AGEMA_signal_10336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C ( clk ), .D ( new_AGEMA_signal_10339 ), .Q ( new_AGEMA_signal_10340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C ( clk ), .D ( new_AGEMA_signal_10343 ), .Q ( new_AGEMA_signal_10344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C ( clk ), .D ( new_AGEMA_signal_10363 ), .Q ( new_AGEMA_signal_10364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C ( clk ), .D ( new_AGEMA_signal_10367 ), .Q ( new_AGEMA_signal_10368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C ( clk ), .D ( new_AGEMA_signal_10371 ), .Q ( new_AGEMA_signal_10372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C ( clk ), .D ( new_AGEMA_signal_10375 ), .Q ( new_AGEMA_signal_10376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C ( clk ), .D ( new_AGEMA_signal_10387 ), .Q ( new_AGEMA_signal_10388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C ( clk ), .D ( new_AGEMA_signal_10391 ), .Q ( new_AGEMA_signal_10392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C ( clk ), .D ( new_AGEMA_signal_10395 ), .Q ( new_AGEMA_signal_10396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C ( clk ), .D ( new_AGEMA_signal_10399 ), .Q ( new_AGEMA_signal_10400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C ( clk ), .D ( new_AGEMA_signal_10411 ), .Q ( new_AGEMA_signal_10412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C ( clk ), .D ( new_AGEMA_signal_10415 ), .Q ( new_AGEMA_signal_10416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C ( clk ), .D ( new_AGEMA_signal_10419 ), .Q ( new_AGEMA_signal_10420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C ( clk ), .D ( new_AGEMA_signal_10423 ), .Q ( new_AGEMA_signal_10424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C ( clk ), .D ( new_AGEMA_signal_10427 ), .Q ( new_AGEMA_signal_10428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C ( clk ), .D ( new_AGEMA_signal_10431 ), .Q ( new_AGEMA_signal_10432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C ( clk ), .D ( new_AGEMA_signal_10435 ), .Q ( new_AGEMA_signal_10436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C ( clk ), .D ( new_AGEMA_signal_10439 ), .Q ( new_AGEMA_signal_10440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C ( clk ), .D ( new_AGEMA_signal_10475 ), .Q ( new_AGEMA_signal_10476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C ( clk ), .D ( new_AGEMA_signal_10479 ), .Q ( new_AGEMA_signal_10480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C ( clk ), .D ( new_AGEMA_signal_10483 ), .Q ( new_AGEMA_signal_10484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C ( clk ), .D ( new_AGEMA_signal_10487 ), .Q ( new_AGEMA_signal_10488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C ( clk ), .D ( new_AGEMA_signal_10491 ), .Q ( new_AGEMA_signal_10492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C ( clk ), .D ( new_AGEMA_signal_10495 ), .Q ( new_AGEMA_signal_10496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C ( clk ), .D ( new_AGEMA_signal_10499 ), .Q ( new_AGEMA_signal_10500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C ( clk ), .D ( new_AGEMA_signal_10503 ), .Q ( new_AGEMA_signal_10504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C ( clk ), .D ( new_AGEMA_signal_10507 ), .Q ( new_AGEMA_signal_10508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C ( clk ), .D ( new_AGEMA_signal_10511 ), .Q ( new_AGEMA_signal_10512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C ( clk ), .D ( new_AGEMA_signal_10515 ), .Q ( new_AGEMA_signal_10516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C ( clk ), .D ( new_AGEMA_signal_10519 ), .Q ( new_AGEMA_signal_10520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C ( clk ), .D ( new_AGEMA_signal_10547 ), .Q ( new_AGEMA_signal_10548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C ( clk ), .D ( new_AGEMA_signal_10551 ), .Q ( new_AGEMA_signal_10552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C ( clk ), .D ( new_AGEMA_signal_10555 ), .Q ( new_AGEMA_signal_10556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C ( clk ), .D ( new_AGEMA_signal_10559 ), .Q ( new_AGEMA_signal_10560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C ( clk ), .D ( new_AGEMA_signal_10571 ), .Q ( new_AGEMA_signal_10572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C ( clk ), .D ( new_AGEMA_signal_10575 ), .Q ( new_AGEMA_signal_10576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C ( clk ), .D ( new_AGEMA_signal_10579 ), .Q ( new_AGEMA_signal_10580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C ( clk ), .D ( new_AGEMA_signal_10583 ), .Q ( new_AGEMA_signal_10584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C ( clk ), .D ( new_AGEMA_signal_10589 ), .Q ( new_AGEMA_signal_10590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C ( clk ), .D ( new_AGEMA_signal_10595 ), .Q ( new_AGEMA_signal_10596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C ( clk ), .D ( new_AGEMA_signal_10601 ), .Q ( new_AGEMA_signal_10602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C ( clk ), .D ( new_AGEMA_signal_10607 ), .Q ( new_AGEMA_signal_10608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C ( clk ), .D ( new_AGEMA_signal_10611 ), .Q ( new_AGEMA_signal_10612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C ( clk ), .D ( new_AGEMA_signal_10615 ), .Q ( new_AGEMA_signal_10616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C ( clk ), .D ( new_AGEMA_signal_10619 ), .Q ( new_AGEMA_signal_10620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C ( clk ), .D ( new_AGEMA_signal_10623 ), .Q ( new_AGEMA_signal_10624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C ( clk ), .D ( new_AGEMA_signal_10627 ), .Q ( new_AGEMA_signal_10628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C ( clk ), .D ( new_AGEMA_signal_10631 ), .Q ( new_AGEMA_signal_10632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C ( clk ), .D ( new_AGEMA_signal_10635 ), .Q ( new_AGEMA_signal_10636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C ( clk ), .D ( new_AGEMA_signal_10639 ), .Q ( new_AGEMA_signal_10640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C ( clk ), .D ( new_AGEMA_signal_10675 ), .Q ( new_AGEMA_signal_10676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C ( clk ), .D ( new_AGEMA_signal_10679 ), .Q ( new_AGEMA_signal_10680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C ( clk ), .D ( new_AGEMA_signal_10683 ), .Q ( new_AGEMA_signal_10684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C ( clk ), .D ( new_AGEMA_signal_10687 ), .Q ( new_AGEMA_signal_10688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C ( clk ), .D ( new_AGEMA_signal_10693 ), .Q ( new_AGEMA_signal_10694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C ( clk ), .D ( new_AGEMA_signal_10699 ), .Q ( new_AGEMA_signal_10700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C ( clk ), .D ( new_AGEMA_signal_10705 ), .Q ( new_AGEMA_signal_10706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C ( clk ), .D ( new_AGEMA_signal_10711 ), .Q ( new_AGEMA_signal_10712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C ( clk ), .D ( new_AGEMA_signal_10715 ), .Q ( new_AGEMA_signal_10716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C ( clk ), .D ( new_AGEMA_signal_10719 ), .Q ( new_AGEMA_signal_10720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C ( clk ), .D ( new_AGEMA_signal_10723 ), .Q ( new_AGEMA_signal_10724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C ( clk ), .D ( new_AGEMA_signal_10727 ), .Q ( new_AGEMA_signal_10728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C ( clk ), .D ( new_AGEMA_signal_10755 ), .Q ( new_AGEMA_signal_10756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C ( clk ), .D ( new_AGEMA_signal_10759 ), .Q ( new_AGEMA_signal_10760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C ( clk ), .D ( new_AGEMA_signal_10763 ), .Q ( new_AGEMA_signal_10764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C ( clk ), .D ( new_AGEMA_signal_10767 ), .Q ( new_AGEMA_signal_10768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C ( clk ), .D ( new_AGEMA_signal_10787 ), .Q ( new_AGEMA_signal_10788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C ( clk ), .D ( new_AGEMA_signal_10791 ), .Q ( new_AGEMA_signal_10792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C ( clk ), .D ( new_AGEMA_signal_10795 ), .Q ( new_AGEMA_signal_10796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C ( clk ), .D ( new_AGEMA_signal_10799 ), .Q ( new_AGEMA_signal_10800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C ( clk ), .D ( new_AGEMA_signal_10803 ), .Q ( new_AGEMA_signal_10804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C ( clk ), .D ( new_AGEMA_signal_10807 ), .Q ( new_AGEMA_signal_10808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C ( clk ), .D ( new_AGEMA_signal_10811 ), .Q ( new_AGEMA_signal_10812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C ( clk ), .D ( new_AGEMA_signal_10815 ), .Q ( new_AGEMA_signal_10816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C ( clk ), .D ( new_AGEMA_signal_10819 ), .Q ( new_AGEMA_signal_10820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C ( clk ), .D ( new_AGEMA_signal_10823 ), .Q ( new_AGEMA_signal_10824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C ( clk ), .D ( new_AGEMA_signal_10827 ), .Q ( new_AGEMA_signal_10828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C ( clk ), .D ( new_AGEMA_signal_10831 ), .Q ( new_AGEMA_signal_10832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C ( clk ), .D ( new_AGEMA_signal_10835 ), .Q ( new_AGEMA_signal_10836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C ( clk ), .D ( new_AGEMA_signal_10839 ), .Q ( new_AGEMA_signal_10840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C ( clk ), .D ( new_AGEMA_signal_10843 ), .Q ( new_AGEMA_signal_10844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C ( clk ), .D ( new_AGEMA_signal_10847 ), .Q ( new_AGEMA_signal_10848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C ( clk ), .D ( new_AGEMA_signal_10851 ), .Q ( new_AGEMA_signal_10852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C ( clk ), .D ( new_AGEMA_signal_10855 ), .Q ( new_AGEMA_signal_10856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C ( clk ), .D ( new_AGEMA_signal_10859 ), .Q ( new_AGEMA_signal_10860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C ( clk ), .D ( new_AGEMA_signal_10863 ), .Q ( new_AGEMA_signal_10864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C ( clk ), .D ( new_AGEMA_signal_10899 ), .Q ( new_AGEMA_signal_10900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C ( clk ), .D ( new_AGEMA_signal_10903 ), .Q ( new_AGEMA_signal_10904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C ( clk ), .D ( new_AGEMA_signal_10907 ), .Q ( new_AGEMA_signal_10908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C ( clk ), .D ( new_AGEMA_signal_10911 ), .Q ( new_AGEMA_signal_10912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C ( clk ), .D ( new_AGEMA_signal_10915 ), .Q ( new_AGEMA_signal_10916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C ( clk ), .D ( new_AGEMA_signal_10919 ), .Q ( new_AGEMA_signal_10920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C ( clk ), .D ( new_AGEMA_signal_10923 ), .Q ( new_AGEMA_signal_10924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C ( clk ), .D ( new_AGEMA_signal_10927 ), .Q ( new_AGEMA_signal_10928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2976 ( .C ( clk ), .D ( new_AGEMA_signal_11003 ), .Q ( new_AGEMA_signal_11004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2980 ( .C ( clk ), .D ( new_AGEMA_signal_11007 ), .Q ( new_AGEMA_signal_11008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2984 ( .C ( clk ), .D ( new_AGEMA_signal_11011 ), .Q ( new_AGEMA_signal_11012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2988 ( .C ( clk ), .D ( new_AGEMA_signal_11015 ), .Q ( new_AGEMA_signal_11016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3032 ( .C ( clk ), .D ( new_AGEMA_signal_11059 ), .Q ( new_AGEMA_signal_11060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3036 ( .C ( clk ), .D ( new_AGEMA_signal_11063 ), .Q ( new_AGEMA_signal_11064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3040 ( .C ( clk ), .D ( new_AGEMA_signal_11067 ), .Q ( new_AGEMA_signal_11068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3044 ( .C ( clk ), .D ( new_AGEMA_signal_11071 ), .Q ( new_AGEMA_signal_11072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3048 ( .C ( clk ), .D ( new_AGEMA_signal_11075 ), .Q ( new_AGEMA_signal_11076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3052 ( .C ( clk ), .D ( new_AGEMA_signal_11079 ), .Q ( new_AGEMA_signal_11080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3056 ( .C ( clk ), .D ( new_AGEMA_signal_11083 ), .Q ( new_AGEMA_signal_11084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3060 ( .C ( clk ), .D ( new_AGEMA_signal_11087 ), .Q ( new_AGEMA_signal_11088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3064 ( .C ( clk ), .D ( new_AGEMA_signal_11091 ), .Q ( new_AGEMA_signal_11092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3068 ( .C ( clk ), .D ( new_AGEMA_signal_11095 ), .Q ( new_AGEMA_signal_11096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3072 ( .C ( clk ), .D ( new_AGEMA_signal_11099 ), .Q ( new_AGEMA_signal_11100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3076 ( .C ( clk ), .D ( new_AGEMA_signal_11103 ), .Q ( new_AGEMA_signal_11104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3080 ( .C ( clk ), .D ( new_AGEMA_signal_11107 ), .Q ( new_AGEMA_signal_11108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3084 ( .C ( clk ), .D ( new_AGEMA_signal_11111 ), .Q ( new_AGEMA_signal_11112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3088 ( .C ( clk ), .D ( new_AGEMA_signal_11115 ), .Q ( new_AGEMA_signal_11116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3092 ( .C ( clk ), .D ( new_AGEMA_signal_11119 ), .Q ( new_AGEMA_signal_11120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3130 ( .C ( clk ), .D ( new_AGEMA_signal_11157 ), .Q ( new_AGEMA_signal_11158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3138 ( .C ( clk ), .D ( new_AGEMA_signal_11165 ), .Q ( new_AGEMA_signal_11166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3146 ( .C ( clk ), .D ( new_AGEMA_signal_11173 ), .Q ( new_AGEMA_signal_11174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3154 ( .C ( clk ), .D ( new_AGEMA_signal_11181 ), .Q ( new_AGEMA_signal_11182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3170 ( .C ( clk ), .D ( new_AGEMA_signal_11197 ), .Q ( new_AGEMA_signal_11198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3178 ( .C ( clk ), .D ( new_AGEMA_signal_11205 ), .Q ( new_AGEMA_signal_11206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3186 ( .C ( clk ), .D ( new_AGEMA_signal_11213 ), .Q ( new_AGEMA_signal_11214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3194 ( .C ( clk ), .D ( new_AGEMA_signal_11221 ), .Q ( new_AGEMA_signal_11222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3200 ( .C ( clk ), .D ( new_AGEMA_signal_11227 ), .Q ( new_AGEMA_signal_11228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3206 ( .C ( clk ), .D ( new_AGEMA_signal_11233 ), .Q ( new_AGEMA_signal_11234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3212 ( .C ( clk ), .D ( new_AGEMA_signal_11239 ), .Q ( new_AGEMA_signal_11240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3218 ( .C ( clk ), .D ( new_AGEMA_signal_11245 ), .Q ( new_AGEMA_signal_11246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3240 ( .C ( clk ), .D ( new_AGEMA_signal_11267 ), .Q ( new_AGEMA_signal_11268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3246 ( .C ( clk ), .D ( new_AGEMA_signal_11273 ), .Q ( new_AGEMA_signal_11274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3252 ( .C ( clk ), .D ( new_AGEMA_signal_11279 ), .Q ( new_AGEMA_signal_11280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3258 ( .C ( clk ), .D ( new_AGEMA_signal_11285 ), .Q ( new_AGEMA_signal_11286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3272 ( .C ( clk ), .D ( new_AGEMA_signal_11299 ), .Q ( new_AGEMA_signal_11300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3278 ( .C ( clk ), .D ( new_AGEMA_signal_11305 ), .Q ( new_AGEMA_signal_11306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3284 ( .C ( clk ), .D ( new_AGEMA_signal_11311 ), .Q ( new_AGEMA_signal_11312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3290 ( .C ( clk ), .D ( new_AGEMA_signal_11317 ), .Q ( new_AGEMA_signal_11318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3296 ( .C ( clk ), .D ( new_AGEMA_signal_11323 ), .Q ( new_AGEMA_signal_11324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3302 ( .C ( clk ), .D ( new_AGEMA_signal_11329 ), .Q ( new_AGEMA_signal_11330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3308 ( .C ( clk ), .D ( new_AGEMA_signal_11335 ), .Q ( new_AGEMA_signal_11336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3314 ( .C ( clk ), .D ( new_AGEMA_signal_11341 ), .Q ( new_AGEMA_signal_11342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3344 ( .C ( clk ), .D ( new_AGEMA_signal_11371 ), .Q ( new_AGEMA_signal_11372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3350 ( .C ( clk ), .D ( new_AGEMA_signal_11377 ), .Q ( new_AGEMA_signal_11378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3356 ( .C ( clk ), .D ( new_AGEMA_signal_11383 ), .Q ( new_AGEMA_signal_11384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3362 ( .C ( clk ), .D ( new_AGEMA_signal_11389 ), .Q ( new_AGEMA_signal_11390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3368 ( .C ( clk ), .D ( new_AGEMA_signal_11395 ), .Q ( new_AGEMA_signal_11396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3374 ( .C ( clk ), .D ( new_AGEMA_signal_11401 ), .Q ( new_AGEMA_signal_11402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3380 ( .C ( clk ), .D ( new_AGEMA_signal_11407 ), .Q ( new_AGEMA_signal_11408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3386 ( .C ( clk ), .D ( new_AGEMA_signal_11413 ), .Q ( new_AGEMA_signal_11414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3400 ( .C ( clk ), .D ( new_AGEMA_signal_11427 ), .Q ( new_AGEMA_signal_11428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3406 ( .C ( clk ), .D ( new_AGEMA_signal_11433 ), .Q ( new_AGEMA_signal_11434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3412 ( .C ( clk ), .D ( new_AGEMA_signal_11439 ), .Q ( new_AGEMA_signal_11440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3418 ( .C ( clk ), .D ( new_AGEMA_signal_11445 ), .Q ( new_AGEMA_signal_11446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3474 ( .C ( clk ), .D ( new_AGEMA_signal_11501 ), .Q ( new_AGEMA_signal_11502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3482 ( .C ( clk ), .D ( new_AGEMA_signal_11509 ), .Q ( new_AGEMA_signal_11510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3490 ( .C ( clk ), .D ( new_AGEMA_signal_11517 ), .Q ( new_AGEMA_signal_11518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3498 ( .C ( clk ), .D ( new_AGEMA_signal_11525 ), .Q ( new_AGEMA_signal_11526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3504 ( .C ( clk ), .D ( new_AGEMA_signal_11531 ), .Q ( new_AGEMA_signal_11532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3510 ( .C ( clk ), .D ( new_AGEMA_signal_11537 ), .Q ( new_AGEMA_signal_11538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3516 ( .C ( clk ), .D ( new_AGEMA_signal_11543 ), .Q ( new_AGEMA_signal_11544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3522 ( .C ( clk ), .D ( new_AGEMA_signal_11549 ), .Q ( new_AGEMA_signal_11550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3616 ( .C ( clk ), .D ( new_AGEMA_signal_11643 ), .Q ( new_AGEMA_signal_11644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3622 ( .C ( clk ), .D ( new_AGEMA_signal_11649 ), .Q ( new_AGEMA_signal_11650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3628 ( .C ( clk ), .D ( new_AGEMA_signal_11655 ), .Q ( new_AGEMA_signal_11656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3634 ( .C ( clk ), .D ( new_AGEMA_signal_11661 ), .Q ( new_AGEMA_signal_11662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3744 ( .C ( clk ), .D ( new_AGEMA_signal_11771 ), .Q ( new_AGEMA_signal_11772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3750 ( .C ( clk ), .D ( new_AGEMA_signal_11777 ), .Q ( new_AGEMA_signal_11778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3756 ( .C ( clk ), .D ( new_AGEMA_signal_11783 ), .Q ( new_AGEMA_signal_11784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3762 ( .C ( clk ), .D ( new_AGEMA_signal_11789 ), .Q ( new_AGEMA_signal_11790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3768 ( .C ( clk ), .D ( new_AGEMA_signal_11795 ), .Q ( new_AGEMA_signal_11796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3774 ( .C ( clk ), .D ( new_AGEMA_signal_11801 ), .Q ( new_AGEMA_signal_11802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3780 ( .C ( clk ), .D ( new_AGEMA_signal_11807 ), .Q ( new_AGEMA_signal_11808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3786 ( .C ( clk ), .D ( new_AGEMA_signal_11813 ), .Q ( new_AGEMA_signal_11814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3818 ( .C ( clk ), .D ( new_AGEMA_signal_11845 ), .Q ( new_AGEMA_signal_11846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3826 ( .C ( clk ), .D ( new_AGEMA_signal_11853 ), .Q ( new_AGEMA_signal_11854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3834 ( .C ( clk ), .D ( new_AGEMA_signal_11861 ), .Q ( new_AGEMA_signal_11862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3842 ( .C ( clk ), .D ( new_AGEMA_signal_11869 ), .Q ( new_AGEMA_signal_11870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3938 ( .C ( clk ), .D ( new_AGEMA_signal_11965 ), .Q ( new_AGEMA_signal_11966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3946 ( .C ( clk ), .D ( new_AGEMA_signal_11973 ), .Q ( new_AGEMA_signal_11974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3954 ( .C ( clk ), .D ( new_AGEMA_signal_11981 ), .Q ( new_AGEMA_signal_11982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3962 ( .C ( clk ), .D ( new_AGEMA_signal_11989 ), .Q ( new_AGEMA_signal_11990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4000 ( .C ( clk ), .D ( new_AGEMA_signal_12027 ), .Q ( new_AGEMA_signal_12028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4006 ( .C ( clk ), .D ( new_AGEMA_signal_12033 ), .Q ( new_AGEMA_signal_12034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4012 ( .C ( clk ), .D ( new_AGEMA_signal_12039 ), .Q ( new_AGEMA_signal_12040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4018 ( .C ( clk ), .D ( new_AGEMA_signal_12045 ), .Q ( new_AGEMA_signal_12046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4032 ( .C ( clk ), .D ( new_AGEMA_signal_12059 ), .Q ( new_AGEMA_signal_12060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4040 ( .C ( clk ), .D ( new_AGEMA_signal_12067 ), .Q ( new_AGEMA_signal_12068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4048 ( .C ( clk ), .D ( new_AGEMA_signal_12075 ), .Q ( new_AGEMA_signal_12076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4056 ( .C ( clk ), .D ( new_AGEMA_signal_12083 ), .Q ( new_AGEMA_signal_12084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4088 ( .C ( clk ), .D ( new_AGEMA_signal_12115 ), .Q ( new_AGEMA_signal_12116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4096 ( .C ( clk ), .D ( new_AGEMA_signal_12123 ), .Q ( new_AGEMA_signal_12124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4104 ( .C ( clk ), .D ( new_AGEMA_signal_12131 ), .Q ( new_AGEMA_signal_12132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4112 ( .C ( clk ), .D ( new_AGEMA_signal_12139 ), .Q ( new_AGEMA_signal_12140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4168 ( .C ( clk ), .D ( new_AGEMA_signal_12195 ), .Q ( new_AGEMA_signal_12196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4176 ( .C ( clk ), .D ( new_AGEMA_signal_12203 ), .Q ( new_AGEMA_signal_12204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4184 ( .C ( clk ), .D ( new_AGEMA_signal_12211 ), .Q ( new_AGEMA_signal_12212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4192 ( .C ( clk ), .D ( new_AGEMA_signal_12219 ), .Q ( new_AGEMA_signal_12220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4352 ( .C ( clk ), .D ( new_AGEMA_signal_12379 ), .Q ( new_AGEMA_signal_12380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4360 ( .C ( clk ), .D ( new_AGEMA_signal_12387 ), .Q ( new_AGEMA_signal_12388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4368 ( .C ( clk ), .D ( new_AGEMA_signal_12395 ), .Q ( new_AGEMA_signal_12396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4376 ( .C ( clk ), .D ( new_AGEMA_signal_12403 ), .Q ( new_AGEMA_signal_12404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4424 ( .C ( clk ), .D ( new_AGEMA_signal_12451 ), .Q ( new_AGEMA_signal_12452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4432 ( .C ( clk ), .D ( new_AGEMA_signal_12459 ), .Q ( new_AGEMA_signal_12460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4440 ( .C ( clk ), .D ( new_AGEMA_signal_12467 ), .Q ( new_AGEMA_signal_12468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4448 ( .C ( clk ), .D ( new_AGEMA_signal_12475 ), .Q ( new_AGEMA_signal_12476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4552 ( .C ( clk ), .D ( new_AGEMA_signal_12579 ), .Q ( new_AGEMA_signal_12580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4560 ( .C ( clk ), .D ( new_AGEMA_signal_12587 ), .Q ( new_AGEMA_signal_12588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4568 ( .C ( clk ), .D ( new_AGEMA_signal_12595 ), .Q ( new_AGEMA_signal_12596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4576 ( .C ( clk ), .D ( new_AGEMA_signal_12603 ), .Q ( new_AGEMA_signal_12604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4584 ( .C ( clk ), .D ( new_AGEMA_signal_12611 ), .Q ( new_AGEMA_signal_12612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4592 ( .C ( clk ), .D ( new_AGEMA_signal_12619 ), .Q ( new_AGEMA_signal_12620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4600 ( .C ( clk ), .D ( new_AGEMA_signal_12627 ), .Q ( new_AGEMA_signal_12628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4608 ( .C ( clk ), .D ( new_AGEMA_signal_12635 ), .Q ( new_AGEMA_signal_12636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4928 ( .C ( clk ), .D ( new_AGEMA_signal_12955 ), .Q ( new_AGEMA_signal_12956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4938 ( .C ( clk ), .D ( new_AGEMA_signal_12965 ), .Q ( new_AGEMA_signal_12966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4948 ( .C ( clk ), .D ( new_AGEMA_signal_12975 ), .Q ( new_AGEMA_signal_12976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4958 ( .C ( clk ), .D ( new_AGEMA_signal_12985 ), .Q ( new_AGEMA_signal_12986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5128 ( .C ( clk ), .D ( new_AGEMA_signal_13155 ), .Q ( new_AGEMA_signal_13156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5138 ( .C ( clk ), .D ( new_AGEMA_signal_13165 ), .Q ( new_AGEMA_signal_13166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5148 ( .C ( clk ), .D ( new_AGEMA_signal_13175 ), .Q ( new_AGEMA_signal_13176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5158 ( .C ( clk ), .D ( new_AGEMA_signal_13185 ), .Q ( new_AGEMA_signal_13186 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_2289 ( .C ( clk ), .D ( new_AGEMA_signal_10316 ), .Q ( new_AGEMA_signal_10317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C ( clk ), .D ( new_AGEMA_signal_10320 ), .Q ( new_AGEMA_signal_10321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C ( clk ), .D ( new_AGEMA_signal_10324 ), .Q ( new_AGEMA_signal_10325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C ( clk ), .D ( new_AGEMA_signal_10328 ), .Q ( new_AGEMA_signal_10329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C ( clk ), .D ( new_AGEMA_signal_10332 ), .Q ( new_AGEMA_signal_10333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C ( clk ), .D ( new_AGEMA_signal_10336 ), .Q ( new_AGEMA_signal_10337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C ( clk ), .D ( new_AGEMA_signal_10340 ), .Q ( new_AGEMA_signal_10341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C ( clk ), .D ( new_AGEMA_signal_10344 ), .Q ( new_AGEMA_signal_10345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C ( clk ), .D ( new_AGEMA_signal_10164 ), .Q ( new_AGEMA_signal_10347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C ( clk ), .D ( new_AGEMA_signal_10166 ), .Q ( new_AGEMA_signal_10349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C ( clk ), .D ( new_AGEMA_signal_10168 ), .Q ( new_AGEMA_signal_10351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C ( clk ), .D ( new_AGEMA_signal_10170 ), .Q ( new_AGEMA_signal_10353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C ( clk ), .D ( n1966 ), .Q ( new_AGEMA_signal_10355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C ( clk ), .D ( new_AGEMA_signal_2079 ), .Q ( new_AGEMA_signal_10357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C ( clk ), .D ( new_AGEMA_signal_2080 ), .Q ( new_AGEMA_signal_10359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C ( clk ), .D ( new_AGEMA_signal_2081 ), .Q ( new_AGEMA_signal_10361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C ( clk ), .D ( new_AGEMA_signal_10364 ), .Q ( new_AGEMA_signal_10365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C ( clk ), .D ( new_AGEMA_signal_10368 ), .Q ( new_AGEMA_signal_10369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C ( clk ), .D ( new_AGEMA_signal_10372 ), .Q ( new_AGEMA_signal_10373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C ( clk ), .D ( new_AGEMA_signal_10376 ), .Q ( new_AGEMA_signal_10377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C ( clk ), .D ( new_AGEMA_signal_10020 ), .Q ( new_AGEMA_signal_10379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C ( clk ), .D ( new_AGEMA_signal_10022 ), .Q ( new_AGEMA_signal_10381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C ( clk ), .D ( new_AGEMA_signal_10024 ), .Q ( new_AGEMA_signal_10383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C ( clk ), .D ( new_AGEMA_signal_10026 ), .Q ( new_AGEMA_signal_10385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C ( clk ), .D ( new_AGEMA_signal_10388 ), .Q ( new_AGEMA_signal_10389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C ( clk ), .D ( new_AGEMA_signal_10392 ), .Q ( new_AGEMA_signal_10393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C ( clk ), .D ( new_AGEMA_signal_10396 ), .Q ( new_AGEMA_signal_10397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C ( clk ), .D ( new_AGEMA_signal_10400 ), .Q ( new_AGEMA_signal_10401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C ( clk ), .D ( n1996 ), .Q ( new_AGEMA_signal_10403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C ( clk ), .D ( new_AGEMA_signal_2109 ), .Q ( new_AGEMA_signal_10405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C ( clk ), .D ( new_AGEMA_signal_2110 ), .Q ( new_AGEMA_signal_10407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C ( clk ), .D ( new_AGEMA_signal_2111 ), .Q ( new_AGEMA_signal_10409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C ( clk ), .D ( new_AGEMA_signal_10412 ), .Q ( new_AGEMA_signal_10413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C ( clk ), .D ( new_AGEMA_signal_10416 ), .Q ( new_AGEMA_signal_10417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C ( clk ), .D ( new_AGEMA_signal_10420 ), .Q ( new_AGEMA_signal_10421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C ( clk ), .D ( new_AGEMA_signal_10424 ), .Q ( new_AGEMA_signal_10425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C ( clk ), .D ( new_AGEMA_signal_10428 ), .Q ( new_AGEMA_signal_10429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C ( clk ), .D ( new_AGEMA_signal_10432 ), .Q ( new_AGEMA_signal_10433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C ( clk ), .D ( new_AGEMA_signal_10436 ), .Q ( new_AGEMA_signal_10437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C ( clk ), .D ( new_AGEMA_signal_10440 ), .Q ( new_AGEMA_signal_10441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C ( clk ), .D ( n2033 ), .Q ( new_AGEMA_signal_10443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C ( clk ), .D ( new_AGEMA_signal_2127 ), .Q ( new_AGEMA_signal_10445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C ( clk ), .D ( new_AGEMA_signal_2128 ), .Q ( new_AGEMA_signal_10447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C ( clk ), .D ( new_AGEMA_signal_2129 ), .Q ( new_AGEMA_signal_10449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C ( clk ), .D ( new_AGEMA_signal_9844 ), .Q ( new_AGEMA_signal_10451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C ( clk ), .D ( new_AGEMA_signal_9846 ), .Q ( new_AGEMA_signal_10453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C ( clk ), .D ( new_AGEMA_signal_9848 ), .Q ( new_AGEMA_signal_10455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C ( clk ), .D ( new_AGEMA_signal_9850 ), .Q ( new_AGEMA_signal_10457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C ( clk ), .D ( new_AGEMA_signal_9884 ), .Q ( new_AGEMA_signal_10459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C ( clk ), .D ( new_AGEMA_signal_9886 ), .Q ( new_AGEMA_signal_10461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C ( clk ), .D ( new_AGEMA_signal_9888 ), .Q ( new_AGEMA_signal_10463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C ( clk ), .D ( new_AGEMA_signal_9890 ), .Q ( new_AGEMA_signal_10465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C ( clk ), .D ( new_AGEMA_signal_9996 ), .Q ( new_AGEMA_signal_10467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C ( clk ), .D ( new_AGEMA_signal_9998 ), .Q ( new_AGEMA_signal_10469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C ( clk ), .D ( new_AGEMA_signal_10000 ), .Q ( new_AGEMA_signal_10471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C ( clk ), .D ( new_AGEMA_signal_10002 ), .Q ( new_AGEMA_signal_10473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C ( clk ), .D ( new_AGEMA_signal_10476 ), .Q ( new_AGEMA_signal_10477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C ( clk ), .D ( new_AGEMA_signal_10480 ), .Q ( new_AGEMA_signal_10481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C ( clk ), .D ( new_AGEMA_signal_10484 ), .Q ( new_AGEMA_signal_10485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C ( clk ), .D ( new_AGEMA_signal_10488 ), .Q ( new_AGEMA_signal_10489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C ( clk ), .D ( new_AGEMA_signal_10492 ), .Q ( new_AGEMA_signal_10493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C ( clk ), .D ( new_AGEMA_signal_10496 ), .Q ( new_AGEMA_signal_10497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C ( clk ), .D ( new_AGEMA_signal_10500 ), .Q ( new_AGEMA_signal_10501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C ( clk ), .D ( new_AGEMA_signal_10504 ), .Q ( new_AGEMA_signal_10505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C ( clk ), .D ( new_AGEMA_signal_10508 ), .Q ( new_AGEMA_signal_10509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C ( clk ), .D ( new_AGEMA_signal_10512 ), .Q ( new_AGEMA_signal_10513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C ( clk ), .D ( new_AGEMA_signal_10516 ), .Q ( new_AGEMA_signal_10517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C ( clk ), .D ( new_AGEMA_signal_10520 ), .Q ( new_AGEMA_signal_10521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C ( clk ), .D ( n2089 ), .Q ( new_AGEMA_signal_10523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C ( clk ), .D ( new_AGEMA_signal_2172 ), .Q ( new_AGEMA_signal_10525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C ( clk ), .D ( new_AGEMA_signal_2173 ), .Q ( new_AGEMA_signal_10527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C ( clk ), .D ( new_AGEMA_signal_2174 ), .Q ( new_AGEMA_signal_10529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C ( clk ), .D ( n2092 ), .Q ( new_AGEMA_signal_10531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C ( clk ), .D ( new_AGEMA_signal_2178 ), .Q ( new_AGEMA_signal_10533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C ( clk ), .D ( new_AGEMA_signal_2179 ), .Q ( new_AGEMA_signal_10535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C ( clk ), .D ( new_AGEMA_signal_2180 ), .Q ( new_AGEMA_signal_10537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C ( clk ), .D ( n2115 ), .Q ( new_AGEMA_signal_10539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C ( clk ), .D ( new_AGEMA_signal_1686 ), .Q ( new_AGEMA_signal_10541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C ( clk ), .D ( new_AGEMA_signal_1687 ), .Q ( new_AGEMA_signal_10543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C ( clk ), .D ( new_AGEMA_signal_1688 ), .Q ( new_AGEMA_signal_10545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C ( clk ), .D ( new_AGEMA_signal_10548 ), .Q ( new_AGEMA_signal_10549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C ( clk ), .D ( new_AGEMA_signal_10552 ), .Q ( new_AGEMA_signal_10553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C ( clk ), .D ( new_AGEMA_signal_10556 ), .Q ( new_AGEMA_signal_10557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C ( clk ), .D ( new_AGEMA_signal_10560 ), .Q ( new_AGEMA_signal_10561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C ( clk ), .D ( n2687 ), .Q ( new_AGEMA_signal_10563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C ( clk ), .D ( new_AGEMA_signal_2076 ), .Q ( new_AGEMA_signal_10565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C ( clk ), .D ( new_AGEMA_signal_2077 ), .Q ( new_AGEMA_signal_10567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C ( clk ), .D ( new_AGEMA_signal_2078 ), .Q ( new_AGEMA_signal_10569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C ( clk ), .D ( new_AGEMA_signal_10572 ), .Q ( new_AGEMA_signal_10573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C ( clk ), .D ( new_AGEMA_signal_10576 ), .Q ( new_AGEMA_signal_10577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C ( clk ), .D ( new_AGEMA_signal_10580 ), .Q ( new_AGEMA_signal_10581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C ( clk ), .D ( new_AGEMA_signal_10584 ), .Q ( new_AGEMA_signal_10585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C ( clk ), .D ( new_AGEMA_signal_10590 ), .Q ( new_AGEMA_signal_10591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C ( clk ), .D ( new_AGEMA_signal_10596 ), .Q ( new_AGEMA_signal_10597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C ( clk ), .D ( new_AGEMA_signal_10602 ), .Q ( new_AGEMA_signal_10603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C ( clk ), .D ( new_AGEMA_signal_10608 ), .Q ( new_AGEMA_signal_10609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C ( clk ), .D ( new_AGEMA_signal_10612 ), .Q ( new_AGEMA_signal_10613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C ( clk ), .D ( new_AGEMA_signal_10616 ), .Q ( new_AGEMA_signal_10617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C ( clk ), .D ( new_AGEMA_signal_10620 ), .Q ( new_AGEMA_signal_10621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C ( clk ), .D ( new_AGEMA_signal_10624 ), .Q ( new_AGEMA_signal_10625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C ( clk ), .D ( new_AGEMA_signal_10628 ), .Q ( new_AGEMA_signal_10629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C ( clk ), .D ( new_AGEMA_signal_10632 ), .Q ( new_AGEMA_signal_10633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C ( clk ), .D ( new_AGEMA_signal_10636 ), .Q ( new_AGEMA_signal_10637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C ( clk ), .D ( new_AGEMA_signal_10640 ), .Q ( new_AGEMA_signal_10641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C ( clk ), .D ( n2193 ), .Q ( new_AGEMA_signal_10643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C ( clk ), .D ( new_AGEMA_signal_2232 ), .Q ( new_AGEMA_signal_10645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C ( clk ), .D ( new_AGEMA_signal_2233 ), .Q ( new_AGEMA_signal_10647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C ( clk ), .D ( new_AGEMA_signal_2234 ), .Q ( new_AGEMA_signal_10649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C ( clk ), .D ( n2202 ), .Q ( new_AGEMA_signal_10651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C ( clk ), .D ( new_AGEMA_signal_2664 ), .Q ( new_AGEMA_signal_10653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C ( clk ), .D ( new_AGEMA_signal_2665 ), .Q ( new_AGEMA_signal_10655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C ( clk ), .D ( new_AGEMA_signal_2666 ), .Q ( new_AGEMA_signal_10657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C ( clk ), .D ( n2228 ), .Q ( new_AGEMA_signal_10659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C ( clk ), .D ( new_AGEMA_signal_1758 ), .Q ( new_AGEMA_signal_10661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C ( clk ), .D ( new_AGEMA_signal_1759 ), .Q ( new_AGEMA_signal_10663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C ( clk ), .D ( new_AGEMA_signal_1760 ), .Q ( new_AGEMA_signal_10665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C ( clk ), .D ( n2235 ), .Q ( new_AGEMA_signal_10667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C ( clk ), .D ( new_AGEMA_signal_2061 ), .Q ( new_AGEMA_signal_10669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C ( clk ), .D ( new_AGEMA_signal_2062 ), .Q ( new_AGEMA_signal_10671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C ( clk ), .D ( new_AGEMA_signal_2063 ), .Q ( new_AGEMA_signal_10673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C ( clk ), .D ( new_AGEMA_signal_10676 ), .Q ( new_AGEMA_signal_10677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C ( clk ), .D ( new_AGEMA_signal_10680 ), .Q ( new_AGEMA_signal_10681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C ( clk ), .D ( new_AGEMA_signal_10684 ), .Q ( new_AGEMA_signal_10685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C ( clk ), .D ( new_AGEMA_signal_10688 ), .Q ( new_AGEMA_signal_10689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C ( clk ), .D ( new_AGEMA_signal_10694 ), .Q ( new_AGEMA_signal_10695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C ( clk ), .D ( new_AGEMA_signal_10700 ), .Q ( new_AGEMA_signal_10701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C ( clk ), .D ( new_AGEMA_signal_10706 ), .Q ( new_AGEMA_signal_10707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C ( clk ), .D ( new_AGEMA_signal_10712 ), .Q ( new_AGEMA_signal_10713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C ( clk ), .D ( new_AGEMA_signal_10716 ), .Q ( new_AGEMA_signal_10717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C ( clk ), .D ( new_AGEMA_signal_10720 ), .Q ( new_AGEMA_signal_10721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C ( clk ), .D ( new_AGEMA_signal_10724 ), .Q ( new_AGEMA_signal_10725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C ( clk ), .D ( new_AGEMA_signal_10728 ), .Q ( new_AGEMA_signal_10729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C ( clk ), .D ( n2752 ), .Q ( new_AGEMA_signal_10731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C ( clk ), .D ( new_AGEMA_signal_2691 ), .Q ( new_AGEMA_signal_10733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C ( clk ), .D ( new_AGEMA_signal_2692 ), .Q ( new_AGEMA_signal_10735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C ( clk ), .D ( new_AGEMA_signal_2693 ), .Q ( new_AGEMA_signal_10737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C ( clk ), .D ( new_AGEMA_signal_10104 ), .Q ( new_AGEMA_signal_10739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C ( clk ), .D ( new_AGEMA_signal_10110 ), .Q ( new_AGEMA_signal_10741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C ( clk ), .D ( new_AGEMA_signal_10116 ), .Q ( new_AGEMA_signal_10743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C ( clk ), .D ( new_AGEMA_signal_10122 ), .Q ( new_AGEMA_signal_10745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C ( clk ), .D ( n2293 ), .Q ( new_AGEMA_signal_10747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C ( clk ), .D ( new_AGEMA_signal_2295 ), .Q ( new_AGEMA_signal_10749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C ( clk ), .D ( new_AGEMA_signal_2296 ), .Q ( new_AGEMA_signal_10751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C ( clk ), .D ( new_AGEMA_signal_2297 ), .Q ( new_AGEMA_signal_10753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C ( clk ), .D ( new_AGEMA_signal_10756 ), .Q ( new_AGEMA_signal_10757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C ( clk ), .D ( new_AGEMA_signal_10760 ), .Q ( new_AGEMA_signal_10761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C ( clk ), .D ( new_AGEMA_signal_10764 ), .Q ( new_AGEMA_signal_10765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C ( clk ), .D ( new_AGEMA_signal_10768 ), .Q ( new_AGEMA_signal_10769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C ( clk ), .D ( n2357 ), .Q ( new_AGEMA_signal_10771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C ( clk ), .D ( new_AGEMA_signal_2322 ), .Q ( new_AGEMA_signal_10773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C ( clk ), .D ( new_AGEMA_signal_2323 ), .Q ( new_AGEMA_signal_10775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C ( clk ), .D ( new_AGEMA_signal_2324 ), .Q ( new_AGEMA_signal_10777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C ( clk ), .D ( n2386 ), .Q ( new_AGEMA_signal_10779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C ( clk ), .D ( new_AGEMA_signal_2337 ), .Q ( new_AGEMA_signal_10781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C ( clk ), .D ( new_AGEMA_signal_2338 ), .Q ( new_AGEMA_signal_10783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C ( clk ), .D ( new_AGEMA_signal_2339 ), .Q ( new_AGEMA_signal_10785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C ( clk ), .D ( new_AGEMA_signal_10788 ), .Q ( new_AGEMA_signal_10789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C ( clk ), .D ( new_AGEMA_signal_10792 ), .Q ( new_AGEMA_signal_10793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C ( clk ), .D ( new_AGEMA_signal_10796 ), .Q ( new_AGEMA_signal_10797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C ( clk ), .D ( new_AGEMA_signal_10800 ), .Q ( new_AGEMA_signal_10801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C ( clk ), .D ( new_AGEMA_signal_10804 ), .Q ( new_AGEMA_signal_10805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C ( clk ), .D ( new_AGEMA_signal_10808 ), .Q ( new_AGEMA_signal_10809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C ( clk ), .D ( new_AGEMA_signal_10812 ), .Q ( new_AGEMA_signal_10813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C ( clk ), .D ( new_AGEMA_signal_10816 ), .Q ( new_AGEMA_signal_10817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C ( clk ), .D ( new_AGEMA_signal_10820 ), .Q ( new_AGEMA_signal_10821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C ( clk ), .D ( new_AGEMA_signal_10824 ), .Q ( new_AGEMA_signal_10825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C ( clk ), .D ( new_AGEMA_signal_10828 ), .Q ( new_AGEMA_signal_10829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C ( clk ), .D ( new_AGEMA_signal_10832 ), .Q ( new_AGEMA_signal_10833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C ( clk ), .D ( new_AGEMA_signal_10836 ), .Q ( new_AGEMA_signal_10837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C ( clk ), .D ( new_AGEMA_signal_10840 ), .Q ( new_AGEMA_signal_10841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C ( clk ), .D ( new_AGEMA_signal_10844 ), .Q ( new_AGEMA_signal_10845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C ( clk ), .D ( new_AGEMA_signal_10848 ), .Q ( new_AGEMA_signal_10849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C ( clk ), .D ( new_AGEMA_signal_10852 ), .Q ( new_AGEMA_signal_10853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C ( clk ), .D ( new_AGEMA_signal_10856 ), .Q ( new_AGEMA_signal_10857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C ( clk ), .D ( new_AGEMA_signal_10860 ), .Q ( new_AGEMA_signal_10861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C ( clk ), .D ( new_AGEMA_signal_10864 ), .Q ( new_AGEMA_signal_10865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C ( clk ), .D ( n2433 ), .Q ( new_AGEMA_signal_10867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C ( clk ), .D ( new_AGEMA_signal_2358 ), .Q ( new_AGEMA_signal_10869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C ( clk ), .D ( new_AGEMA_signal_2359 ), .Q ( new_AGEMA_signal_10871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C ( clk ), .D ( new_AGEMA_signal_2360 ), .Q ( new_AGEMA_signal_10873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C ( clk ), .D ( new_AGEMA_signal_9870 ), .Q ( new_AGEMA_signal_10875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C ( clk ), .D ( new_AGEMA_signal_9874 ), .Q ( new_AGEMA_signal_10877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C ( clk ), .D ( new_AGEMA_signal_9878 ), .Q ( new_AGEMA_signal_10879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C ( clk ), .D ( new_AGEMA_signal_9882 ), .Q ( new_AGEMA_signal_10881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C ( clk ), .D ( n2459 ), .Q ( new_AGEMA_signal_10883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C ( clk ), .D ( new_AGEMA_signal_2286 ), .Q ( new_AGEMA_signal_10885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C ( clk ), .D ( new_AGEMA_signal_2287 ), .Q ( new_AGEMA_signal_10887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C ( clk ), .D ( new_AGEMA_signal_2288 ), .Q ( new_AGEMA_signal_10889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C ( clk ), .D ( n2467 ), .Q ( new_AGEMA_signal_10891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C ( clk ), .D ( new_AGEMA_signal_1854 ), .Q ( new_AGEMA_signal_10893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C ( clk ), .D ( new_AGEMA_signal_1855 ), .Q ( new_AGEMA_signal_10895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C ( clk ), .D ( new_AGEMA_signal_1856 ), .Q ( new_AGEMA_signal_10897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C ( clk ), .D ( new_AGEMA_signal_10900 ), .Q ( new_AGEMA_signal_10901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C ( clk ), .D ( new_AGEMA_signal_10904 ), .Q ( new_AGEMA_signal_10905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C ( clk ), .D ( new_AGEMA_signal_10908 ), .Q ( new_AGEMA_signal_10909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C ( clk ), .D ( new_AGEMA_signal_10912 ), .Q ( new_AGEMA_signal_10913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C ( clk ), .D ( new_AGEMA_signal_10916 ), .Q ( new_AGEMA_signal_10917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C ( clk ), .D ( new_AGEMA_signal_10920 ), .Q ( new_AGEMA_signal_10921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C ( clk ), .D ( new_AGEMA_signal_10924 ), .Q ( new_AGEMA_signal_10925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C ( clk ), .D ( new_AGEMA_signal_10928 ), .Q ( new_AGEMA_signal_10929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C ( clk ), .D ( n2489 ), .Q ( new_AGEMA_signal_10931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C ( clk ), .D ( new_AGEMA_signal_1914 ), .Q ( new_AGEMA_signal_10933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C ( clk ), .D ( new_AGEMA_signal_1915 ), .Q ( new_AGEMA_signal_10935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C ( clk ), .D ( new_AGEMA_signal_1916 ), .Q ( new_AGEMA_signal_10937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C ( clk ), .D ( n2497 ), .Q ( new_AGEMA_signal_10939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C ( clk ), .D ( new_AGEMA_signal_1917 ), .Q ( new_AGEMA_signal_10941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C ( clk ), .D ( new_AGEMA_signal_1918 ), .Q ( new_AGEMA_signal_10943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C ( clk ), .D ( new_AGEMA_signal_1919 ), .Q ( new_AGEMA_signal_10945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C ( clk ), .D ( n2506 ), .Q ( new_AGEMA_signal_10947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C ( clk ), .D ( new_AGEMA_signal_2397 ), .Q ( new_AGEMA_signal_10949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C ( clk ), .D ( new_AGEMA_signal_2398 ), .Q ( new_AGEMA_signal_10951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2925 ( .C ( clk ), .D ( new_AGEMA_signal_2399 ), .Q ( new_AGEMA_signal_10953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2927 ( .C ( clk ), .D ( n2542 ), .Q ( new_AGEMA_signal_10955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2929 ( .C ( clk ), .D ( new_AGEMA_signal_2415 ), .Q ( new_AGEMA_signal_10957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2931 ( .C ( clk ), .D ( new_AGEMA_signal_2416 ), .Q ( new_AGEMA_signal_10959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C ( clk ), .D ( new_AGEMA_signal_2417 ), .Q ( new_AGEMA_signal_10961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C ( clk ), .D ( n2558 ), .Q ( new_AGEMA_signal_10963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2937 ( .C ( clk ), .D ( new_AGEMA_signal_2424 ), .Q ( new_AGEMA_signal_10965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2939 ( .C ( clk ), .D ( new_AGEMA_signal_2425 ), .Q ( new_AGEMA_signal_10967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2941 ( .C ( clk ), .D ( new_AGEMA_signal_2426 ), .Q ( new_AGEMA_signal_10969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2943 ( .C ( clk ), .D ( n2566 ), .Q ( new_AGEMA_signal_10971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2945 ( .C ( clk ), .D ( new_AGEMA_signal_2430 ), .Q ( new_AGEMA_signal_10973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2947 ( .C ( clk ), .D ( new_AGEMA_signal_2431 ), .Q ( new_AGEMA_signal_10975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2949 ( .C ( clk ), .D ( new_AGEMA_signal_2432 ), .Q ( new_AGEMA_signal_10977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2951 ( .C ( clk ), .D ( n2581 ), .Q ( new_AGEMA_signal_10979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2953 ( .C ( clk ), .D ( new_AGEMA_signal_1944 ), .Q ( new_AGEMA_signal_10981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2955 ( .C ( clk ), .D ( new_AGEMA_signal_1945 ), .Q ( new_AGEMA_signal_10983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2957 ( .C ( clk ), .D ( new_AGEMA_signal_1946 ), .Q ( new_AGEMA_signal_10985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2959 ( .C ( clk ), .D ( n2603 ), .Q ( new_AGEMA_signal_10987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2961 ( .C ( clk ), .D ( new_AGEMA_signal_2454 ), .Q ( new_AGEMA_signal_10989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2963 ( .C ( clk ), .D ( new_AGEMA_signal_2455 ), .Q ( new_AGEMA_signal_10991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2965 ( .C ( clk ), .D ( new_AGEMA_signal_2456 ), .Q ( new_AGEMA_signal_10993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2967 ( .C ( clk ), .D ( n2620 ), .Q ( new_AGEMA_signal_10995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2969 ( .C ( clk ), .D ( new_AGEMA_signal_2457 ), .Q ( new_AGEMA_signal_10997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2971 ( .C ( clk ), .D ( new_AGEMA_signal_2458 ), .Q ( new_AGEMA_signal_10999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2973 ( .C ( clk ), .D ( new_AGEMA_signal_2459 ), .Q ( new_AGEMA_signal_11001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2977 ( .C ( clk ), .D ( new_AGEMA_signal_11004 ), .Q ( new_AGEMA_signal_11005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2981 ( .C ( clk ), .D ( new_AGEMA_signal_11008 ), .Q ( new_AGEMA_signal_11009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2985 ( .C ( clk ), .D ( new_AGEMA_signal_11012 ), .Q ( new_AGEMA_signal_11013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2989 ( .C ( clk ), .D ( new_AGEMA_signal_11016 ), .Q ( new_AGEMA_signal_11017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2991 ( .C ( clk ), .D ( n2653 ), .Q ( new_AGEMA_signal_11019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2993 ( .C ( clk ), .D ( new_AGEMA_signal_1983 ), .Q ( new_AGEMA_signal_11021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2995 ( .C ( clk ), .D ( new_AGEMA_signal_1984 ), .Q ( new_AGEMA_signal_11023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2997 ( .C ( clk ), .D ( new_AGEMA_signal_1985 ), .Q ( new_AGEMA_signal_11025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2999 ( .C ( clk ), .D ( n2665 ), .Q ( new_AGEMA_signal_11027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3001 ( .C ( clk ), .D ( new_AGEMA_signal_2055 ), .Q ( new_AGEMA_signal_11029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3003 ( .C ( clk ), .D ( new_AGEMA_signal_2056 ), .Q ( new_AGEMA_signal_11031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3005 ( .C ( clk ), .D ( new_AGEMA_signal_2057 ), .Q ( new_AGEMA_signal_11033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3007 ( .C ( clk ), .D ( n2691 ), .Q ( new_AGEMA_signal_11035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3009 ( .C ( clk ), .D ( new_AGEMA_signal_1992 ), .Q ( new_AGEMA_signal_11037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3011 ( .C ( clk ), .D ( new_AGEMA_signal_1993 ), .Q ( new_AGEMA_signal_11039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3013 ( .C ( clk ), .D ( new_AGEMA_signal_1994 ), .Q ( new_AGEMA_signal_11041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3015 ( .C ( clk ), .D ( n2717 ), .Q ( new_AGEMA_signal_11043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3017 ( .C ( clk ), .D ( new_AGEMA_signal_2484 ), .Q ( new_AGEMA_signal_11045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3019 ( .C ( clk ), .D ( new_AGEMA_signal_2485 ), .Q ( new_AGEMA_signal_11047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3021 ( .C ( clk ), .D ( new_AGEMA_signal_2486 ), .Q ( new_AGEMA_signal_11049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3023 ( .C ( clk ), .D ( n2729 ), .Q ( new_AGEMA_signal_11051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3025 ( .C ( clk ), .D ( new_AGEMA_signal_2844 ), .Q ( new_AGEMA_signal_11053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3027 ( .C ( clk ), .D ( new_AGEMA_signal_2845 ), .Q ( new_AGEMA_signal_11055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3029 ( .C ( clk ), .D ( new_AGEMA_signal_2846 ), .Q ( new_AGEMA_signal_11057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3033 ( .C ( clk ), .D ( new_AGEMA_signal_11060 ), .Q ( new_AGEMA_signal_11061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3037 ( .C ( clk ), .D ( new_AGEMA_signal_11064 ), .Q ( new_AGEMA_signal_11065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3041 ( .C ( clk ), .D ( new_AGEMA_signal_11068 ), .Q ( new_AGEMA_signal_11069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3045 ( .C ( clk ), .D ( new_AGEMA_signal_11072 ), .Q ( new_AGEMA_signal_11073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3049 ( .C ( clk ), .D ( new_AGEMA_signal_11076 ), .Q ( new_AGEMA_signal_11077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3053 ( .C ( clk ), .D ( new_AGEMA_signal_11080 ), .Q ( new_AGEMA_signal_11081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3057 ( .C ( clk ), .D ( new_AGEMA_signal_11084 ), .Q ( new_AGEMA_signal_11085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3061 ( .C ( clk ), .D ( new_AGEMA_signal_11088 ), .Q ( new_AGEMA_signal_11089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3065 ( .C ( clk ), .D ( new_AGEMA_signal_11092 ), .Q ( new_AGEMA_signal_11093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3069 ( .C ( clk ), .D ( new_AGEMA_signal_11096 ), .Q ( new_AGEMA_signal_11097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3073 ( .C ( clk ), .D ( new_AGEMA_signal_11100 ), .Q ( new_AGEMA_signal_11101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3077 ( .C ( clk ), .D ( new_AGEMA_signal_11104 ), .Q ( new_AGEMA_signal_11105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3081 ( .C ( clk ), .D ( new_AGEMA_signal_11108 ), .Q ( new_AGEMA_signal_11109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3085 ( .C ( clk ), .D ( new_AGEMA_signal_11112 ), .Q ( new_AGEMA_signal_11113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3089 ( .C ( clk ), .D ( new_AGEMA_signal_11116 ), .Q ( new_AGEMA_signal_11117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3093 ( .C ( clk ), .D ( new_AGEMA_signal_11120 ), .Q ( new_AGEMA_signal_11121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3095 ( .C ( clk ), .D ( new_AGEMA_signal_10052 ), .Q ( new_AGEMA_signal_11123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3099 ( .C ( clk ), .D ( new_AGEMA_signal_10054 ), .Q ( new_AGEMA_signal_11127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3103 ( .C ( clk ), .D ( new_AGEMA_signal_10056 ), .Q ( new_AGEMA_signal_11131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3107 ( .C ( clk ), .D ( new_AGEMA_signal_10058 ), .Q ( new_AGEMA_signal_11135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3111 ( .C ( clk ), .D ( n1956 ), .Q ( new_AGEMA_signal_11139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3115 ( .C ( clk ), .D ( new_AGEMA_signal_2067 ), .Q ( new_AGEMA_signal_11143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3119 ( .C ( clk ), .D ( new_AGEMA_signal_2068 ), .Q ( new_AGEMA_signal_11147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3123 ( .C ( clk ), .D ( new_AGEMA_signal_2069 ), .Q ( new_AGEMA_signal_11151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3131 ( .C ( clk ), .D ( new_AGEMA_signal_11158 ), .Q ( new_AGEMA_signal_11159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3139 ( .C ( clk ), .D ( new_AGEMA_signal_11166 ), .Q ( new_AGEMA_signal_11167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3147 ( .C ( clk ), .D ( new_AGEMA_signal_11174 ), .Q ( new_AGEMA_signal_11175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3155 ( .C ( clk ), .D ( new_AGEMA_signal_11182 ), .Q ( new_AGEMA_signal_11183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3171 ( .C ( clk ), .D ( new_AGEMA_signal_11198 ), .Q ( new_AGEMA_signal_11199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3179 ( .C ( clk ), .D ( new_AGEMA_signal_11206 ), .Q ( new_AGEMA_signal_11207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3187 ( .C ( clk ), .D ( new_AGEMA_signal_11214 ), .Q ( new_AGEMA_signal_11215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3195 ( .C ( clk ), .D ( new_AGEMA_signal_11222 ), .Q ( new_AGEMA_signal_11223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3201 ( .C ( clk ), .D ( new_AGEMA_signal_11228 ), .Q ( new_AGEMA_signal_11229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3207 ( .C ( clk ), .D ( new_AGEMA_signal_11234 ), .Q ( new_AGEMA_signal_11235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3213 ( .C ( clk ), .D ( new_AGEMA_signal_11240 ), .Q ( new_AGEMA_signal_11241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3219 ( .C ( clk ), .D ( new_AGEMA_signal_11246 ), .Q ( new_AGEMA_signal_11247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3223 ( .C ( clk ), .D ( n2023 ), .Q ( new_AGEMA_signal_11251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3227 ( .C ( clk ), .D ( new_AGEMA_signal_1614 ), .Q ( new_AGEMA_signal_11255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3231 ( .C ( clk ), .D ( new_AGEMA_signal_1615 ), .Q ( new_AGEMA_signal_11259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3235 ( .C ( clk ), .D ( new_AGEMA_signal_1616 ), .Q ( new_AGEMA_signal_11263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3241 ( .C ( clk ), .D ( new_AGEMA_signal_11268 ), .Q ( new_AGEMA_signal_11269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3247 ( .C ( clk ), .D ( new_AGEMA_signal_11274 ), .Q ( new_AGEMA_signal_11275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3253 ( .C ( clk ), .D ( new_AGEMA_signal_11280 ), .Q ( new_AGEMA_signal_11281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3259 ( .C ( clk ), .D ( new_AGEMA_signal_11286 ), .Q ( new_AGEMA_signal_11287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3273 ( .C ( clk ), .D ( new_AGEMA_signal_11300 ), .Q ( new_AGEMA_signal_11301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3279 ( .C ( clk ), .D ( new_AGEMA_signal_11306 ), .Q ( new_AGEMA_signal_11307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3285 ( .C ( clk ), .D ( new_AGEMA_signal_11312 ), .Q ( new_AGEMA_signal_11313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3291 ( .C ( clk ), .D ( new_AGEMA_signal_11318 ), .Q ( new_AGEMA_signal_11319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3297 ( .C ( clk ), .D ( new_AGEMA_signal_11324 ), .Q ( new_AGEMA_signal_11325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3303 ( .C ( clk ), .D ( new_AGEMA_signal_11330 ), .Q ( new_AGEMA_signal_11331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3309 ( .C ( clk ), .D ( new_AGEMA_signal_11336 ), .Q ( new_AGEMA_signal_11337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3315 ( .C ( clk ), .D ( new_AGEMA_signal_11342 ), .Q ( new_AGEMA_signal_11343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3327 ( .C ( clk ), .D ( n2094 ), .Q ( new_AGEMA_signal_11355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3331 ( .C ( clk ), .D ( new_AGEMA_signal_2181 ), .Q ( new_AGEMA_signal_11359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3335 ( .C ( clk ), .D ( new_AGEMA_signal_2182 ), .Q ( new_AGEMA_signal_11363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3339 ( .C ( clk ), .D ( new_AGEMA_signal_2183 ), .Q ( new_AGEMA_signal_11367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3345 ( .C ( clk ), .D ( new_AGEMA_signal_11372 ), .Q ( new_AGEMA_signal_11373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3351 ( .C ( clk ), .D ( new_AGEMA_signal_11378 ), .Q ( new_AGEMA_signal_11379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3357 ( .C ( clk ), .D ( new_AGEMA_signal_11384 ), .Q ( new_AGEMA_signal_11385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3363 ( .C ( clk ), .D ( new_AGEMA_signal_11390 ), .Q ( new_AGEMA_signal_11391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3369 ( .C ( clk ), .D ( new_AGEMA_signal_11396 ), .Q ( new_AGEMA_signal_11397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3375 ( .C ( clk ), .D ( new_AGEMA_signal_11402 ), .Q ( new_AGEMA_signal_11403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3381 ( .C ( clk ), .D ( new_AGEMA_signal_11408 ), .Q ( new_AGEMA_signal_11409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3387 ( .C ( clk ), .D ( new_AGEMA_signal_11414 ), .Q ( new_AGEMA_signal_11415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3401 ( .C ( clk ), .D ( new_AGEMA_signal_11428 ), .Q ( new_AGEMA_signal_11429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3407 ( .C ( clk ), .D ( new_AGEMA_signal_11434 ), .Q ( new_AGEMA_signal_11435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3413 ( .C ( clk ), .D ( new_AGEMA_signal_11440 ), .Q ( new_AGEMA_signal_11441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3419 ( .C ( clk ), .D ( new_AGEMA_signal_11446 ), .Q ( new_AGEMA_signal_11447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3431 ( .C ( clk ), .D ( n2181 ), .Q ( new_AGEMA_signal_11459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3435 ( .C ( clk ), .D ( new_AGEMA_signal_2223 ), .Q ( new_AGEMA_signal_11463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3439 ( .C ( clk ), .D ( new_AGEMA_signal_2224 ), .Q ( new_AGEMA_signal_11467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3443 ( .C ( clk ), .D ( new_AGEMA_signal_2225 ), .Q ( new_AGEMA_signal_11471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3447 ( .C ( clk ), .D ( n2195 ), .Q ( new_AGEMA_signal_11475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3451 ( .C ( clk ), .D ( new_AGEMA_signal_2229 ), .Q ( new_AGEMA_signal_11479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3455 ( .C ( clk ), .D ( new_AGEMA_signal_2230 ), .Q ( new_AGEMA_signal_11483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3459 ( .C ( clk ), .D ( new_AGEMA_signal_2231 ), .Q ( new_AGEMA_signal_11487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3475 ( .C ( clk ), .D ( new_AGEMA_signal_11502 ), .Q ( new_AGEMA_signal_11503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3483 ( .C ( clk ), .D ( new_AGEMA_signal_11510 ), .Q ( new_AGEMA_signal_11511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3491 ( .C ( clk ), .D ( new_AGEMA_signal_11518 ), .Q ( new_AGEMA_signal_11519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3499 ( .C ( clk ), .D ( new_AGEMA_signal_11526 ), .Q ( new_AGEMA_signal_11527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3505 ( .C ( clk ), .D ( new_AGEMA_signal_11532 ), .Q ( new_AGEMA_signal_11533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3511 ( .C ( clk ), .D ( new_AGEMA_signal_11538 ), .Q ( new_AGEMA_signal_11539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3517 ( .C ( clk ), .D ( new_AGEMA_signal_11544 ), .Q ( new_AGEMA_signal_11545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3523 ( .C ( clk ), .D ( new_AGEMA_signal_11550 ), .Q ( new_AGEMA_signal_11551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3527 ( .C ( clk ), .D ( n2237 ), .Q ( new_AGEMA_signal_11555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3531 ( .C ( clk ), .D ( new_AGEMA_signal_1761 ), .Q ( new_AGEMA_signal_11559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3535 ( .C ( clk ), .D ( new_AGEMA_signal_1762 ), .Q ( new_AGEMA_signal_11563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3539 ( .C ( clk ), .D ( new_AGEMA_signal_1763 ), .Q ( new_AGEMA_signal_11567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3543 ( .C ( clk ), .D ( n2248 ), .Q ( new_AGEMA_signal_11571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3547 ( .C ( clk ), .D ( new_AGEMA_signal_2256 ), .Q ( new_AGEMA_signal_11575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3551 ( .C ( clk ), .D ( new_AGEMA_signal_2257 ), .Q ( new_AGEMA_signal_11579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3555 ( .C ( clk ), .D ( new_AGEMA_signal_2258 ), .Q ( new_AGEMA_signal_11583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3575 ( .C ( clk ), .D ( n2294 ), .Q ( new_AGEMA_signal_11603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3579 ( .C ( clk ), .D ( new_AGEMA_signal_1806 ), .Q ( new_AGEMA_signal_11607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3583 ( .C ( clk ), .D ( new_AGEMA_signal_1807 ), .Q ( new_AGEMA_signal_11611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3587 ( .C ( clk ), .D ( new_AGEMA_signal_1808 ), .Q ( new_AGEMA_signal_11615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3591 ( .C ( clk ), .D ( n2323 ), .Q ( new_AGEMA_signal_11619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3595 ( .C ( clk ), .D ( new_AGEMA_signal_2301 ), .Q ( new_AGEMA_signal_11623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3599 ( .C ( clk ), .D ( new_AGEMA_signal_2302 ), .Q ( new_AGEMA_signal_11627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3603 ( .C ( clk ), .D ( new_AGEMA_signal_2303 ), .Q ( new_AGEMA_signal_11631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3617 ( .C ( clk ), .D ( new_AGEMA_signal_11644 ), .Q ( new_AGEMA_signal_11645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3623 ( .C ( clk ), .D ( new_AGEMA_signal_11650 ), .Q ( new_AGEMA_signal_11651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3629 ( .C ( clk ), .D ( new_AGEMA_signal_11656 ), .Q ( new_AGEMA_signal_11657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3635 ( .C ( clk ), .D ( new_AGEMA_signal_11662 ), .Q ( new_AGEMA_signal_11663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3639 ( .C ( clk ), .D ( n2360 ), .Q ( new_AGEMA_signal_11667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3643 ( .C ( clk ), .D ( new_AGEMA_signal_2325 ), .Q ( new_AGEMA_signal_11671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3647 ( .C ( clk ), .D ( new_AGEMA_signal_2326 ), .Q ( new_AGEMA_signal_11675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3651 ( .C ( clk ), .D ( new_AGEMA_signal_2327 ), .Q ( new_AGEMA_signal_11679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3663 ( .C ( clk ), .D ( n2394 ), .Q ( new_AGEMA_signal_11691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3667 ( .C ( clk ), .D ( new_AGEMA_signal_1863 ), .Q ( new_AGEMA_signal_11695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3671 ( .C ( clk ), .D ( new_AGEMA_signal_1864 ), .Q ( new_AGEMA_signal_11699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3675 ( .C ( clk ), .D ( new_AGEMA_signal_1865 ), .Q ( new_AGEMA_signal_11703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3679 ( .C ( clk ), .D ( n2406 ), .Q ( new_AGEMA_signal_11707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3683 ( .C ( clk ), .D ( new_AGEMA_signal_2343 ), .Q ( new_AGEMA_signal_11711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3687 ( .C ( clk ), .D ( new_AGEMA_signal_2344 ), .Q ( new_AGEMA_signal_11715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3691 ( .C ( clk ), .D ( new_AGEMA_signal_2345 ), .Q ( new_AGEMA_signal_11719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3695 ( .C ( clk ), .D ( new_AGEMA_signal_9652 ), .Q ( new_AGEMA_signal_11723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3699 ( .C ( clk ), .D ( new_AGEMA_signal_9654 ), .Q ( new_AGEMA_signal_11727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3703 ( .C ( clk ), .D ( new_AGEMA_signal_9656 ), .Q ( new_AGEMA_signal_11731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3707 ( .C ( clk ), .D ( new_AGEMA_signal_9658 ), .Q ( new_AGEMA_signal_11735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3719 ( .C ( clk ), .D ( new_AGEMA_signal_9660 ), .Q ( new_AGEMA_signal_11747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3723 ( .C ( clk ), .D ( new_AGEMA_signal_9662 ), .Q ( new_AGEMA_signal_11751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3727 ( .C ( clk ), .D ( new_AGEMA_signal_9664 ), .Q ( new_AGEMA_signal_11755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3731 ( .C ( clk ), .D ( new_AGEMA_signal_9666 ), .Q ( new_AGEMA_signal_11759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3745 ( .C ( clk ), .D ( new_AGEMA_signal_11772 ), .Q ( new_AGEMA_signal_11773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3751 ( .C ( clk ), .D ( new_AGEMA_signal_11778 ), .Q ( new_AGEMA_signal_11779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3757 ( .C ( clk ), .D ( new_AGEMA_signal_11784 ), .Q ( new_AGEMA_signal_11785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3763 ( .C ( clk ), .D ( new_AGEMA_signal_11790 ), .Q ( new_AGEMA_signal_11791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3769 ( .C ( clk ), .D ( new_AGEMA_signal_11796 ), .Q ( new_AGEMA_signal_11797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3775 ( .C ( clk ), .D ( new_AGEMA_signal_11802 ), .Q ( new_AGEMA_signal_11803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3781 ( .C ( clk ), .D ( new_AGEMA_signal_11808 ), .Q ( new_AGEMA_signal_11809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3787 ( .C ( clk ), .D ( new_AGEMA_signal_11814 ), .Q ( new_AGEMA_signal_11815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3791 ( .C ( clk ), .D ( n2499 ), .Q ( new_AGEMA_signal_11819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3795 ( .C ( clk ), .D ( new_AGEMA_signal_1923 ), .Q ( new_AGEMA_signal_11823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3799 ( .C ( clk ), .D ( new_AGEMA_signal_1924 ), .Q ( new_AGEMA_signal_11827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3803 ( .C ( clk ), .D ( new_AGEMA_signal_1925 ), .Q ( new_AGEMA_signal_11831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3819 ( .C ( clk ), .D ( new_AGEMA_signal_11846 ), .Q ( new_AGEMA_signal_11847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3827 ( .C ( clk ), .D ( new_AGEMA_signal_11854 ), .Q ( new_AGEMA_signal_11855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3835 ( .C ( clk ), .D ( new_AGEMA_signal_11862 ), .Q ( new_AGEMA_signal_11863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3843 ( .C ( clk ), .D ( new_AGEMA_signal_11870 ), .Q ( new_AGEMA_signal_11871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3855 ( .C ( clk ), .D ( n2582 ), .Q ( new_AGEMA_signal_11883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3859 ( .C ( clk ), .D ( new_AGEMA_signal_2445 ), .Q ( new_AGEMA_signal_11887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3863 ( .C ( clk ), .D ( new_AGEMA_signal_2446 ), .Q ( new_AGEMA_signal_11891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3867 ( .C ( clk ), .D ( new_AGEMA_signal_2447 ), .Q ( new_AGEMA_signal_11895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3871 ( .C ( clk ), .D ( n2605 ), .Q ( new_AGEMA_signal_11899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3875 ( .C ( clk ), .D ( new_AGEMA_signal_2451 ), .Q ( new_AGEMA_signal_11903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3879 ( .C ( clk ), .D ( new_AGEMA_signal_2452 ), .Q ( new_AGEMA_signal_11907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3883 ( .C ( clk ), .D ( new_AGEMA_signal_2453 ), .Q ( new_AGEMA_signal_11911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3887 ( .C ( clk ), .D ( n2632 ), .Q ( new_AGEMA_signal_11915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3891 ( .C ( clk ), .D ( new_AGEMA_signal_1974 ), .Q ( new_AGEMA_signal_11919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3895 ( .C ( clk ), .D ( new_AGEMA_signal_1975 ), .Q ( new_AGEMA_signal_11923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3899 ( .C ( clk ), .D ( new_AGEMA_signal_1976 ), .Q ( new_AGEMA_signal_11927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3903 ( .C ( clk ), .D ( n2655 ), .Q ( new_AGEMA_signal_11931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3907 ( .C ( clk ), .D ( new_AGEMA_signal_2472 ), .Q ( new_AGEMA_signal_11935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3911 ( .C ( clk ), .D ( new_AGEMA_signal_2473 ), .Q ( new_AGEMA_signal_11939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3915 ( .C ( clk ), .D ( new_AGEMA_signal_2474 ), .Q ( new_AGEMA_signal_11943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3919 ( .C ( clk ), .D ( n2695 ), .Q ( new_AGEMA_signal_11947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3923 ( .C ( clk ), .D ( new_AGEMA_signal_2481 ), .Q ( new_AGEMA_signal_11951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3927 ( .C ( clk ), .D ( new_AGEMA_signal_2482 ), .Q ( new_AGEMA_signal_11955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3931 ( .C ( clk ), .D ( new_AGEMA_signal_2483 ), .Q ( new_AGEMA_signal_11959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3939 ( .C ( clk ), .D ( new_AGEMA_signal_11966 ), .Q ( new_AGEMA_signal_11967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3947 ( .C ( clk ), .D ( new_AGEMA_signal_11974 ), .Q ( new_AGEMA_signal_11975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3955 ( .C ( clk ), .D ( new_AGEMA_signal_11982 ), .Q ( new_AGEMA_signal_11983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3963 ( .C ( clk ), .D ( new_AGEMA_signal_11990 ), .Q ( new_AGEMA_signal_11991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3975 ( .C ( clk ), .D ( n2770 ), .Q ( new_AGEMA_signal_12003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3979 ( .C ( clk ), .D ( new_AGEMA_signal_2505 ), .Q ( new_AGEMA_signal_12007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3983 ( .C ( clk ), .D ( new_AGEMA_signal_2506 ), .Q ( new_AGEMA_signal_12011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3987 ( .C ( clk ), .D ( new_AGEMA_signal_2507 ), .Q ( new_AGEMA_signal_12015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4001 ( .C ( clk ), .D ( new_AGEMA_signal_12028 ), .Q ( new_AGEMA_signal_12029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4007 ( .C ( clk ), .D ( new_AGEMA_signal_12034 ), .Q ( new_AGEMA_signal_12035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4013 ( .C ( clk ), .D ( new_AGEMA_signal_12040 ), .Q ( new_AGEMA_signal_12041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4019 ( .C ( clk ), .D ( new_AGEMA_signal_12046 ), .Q ( new_AGEMA_signal_12047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4033 ( .C ( clk ), .D ( new_AGEMA_signal_12060 ), .Q ( new_AGEMA_signal_12061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4041 ( .C ( clk ), .D ( new_AGEMA_signal_12068 ), .Q ( new_AGEMA_signal_12069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4049 ( .C ( clk ), .D ( new_AGEMA_signal_12076 ), .Q ( new_AGEMA_signal_12077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4057 ( .C ( clk ), .D ( new_AGEMA_signal_12084 ), .Q ( new_AGEMA_signal_12085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4089 ( .C ( clk ), .D ( new_AGEMA_signal_12116 ), .Q ( new_AGEMA_signal_12117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4097 ( .C ( clk ), .D ( new_AGEMA_signal_12124 ), .Q ( new_AGEMA_signal_12125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4105 ( .C ( clk ), .D ( new_AGEMA_signal_12132 ), .Q ( new_AGEMA_signal_12133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4113 ( .C ( clk ), .D ( new_AGEMA_signal_12140 ), .Q ( new_AGEMA_signal_12141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4127 ( .C ( clk ), .D ( n2050 ), .Q ( new_AGEMA_signal_12155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4133 ( .C ( clk ), .D ( new_AGEMA_signal_1629 ), .Q ( new_AGEMA_signal_12161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4139 ( .C ( clk ), .D ( new_AGEMA_signal_1630 ), .Q ( new_AGEMA_signal_12167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4145 ( .C ( clk ), .D ( new_AGEMA_signal_1631 ), .Q ( new_AGEMA_signal_12173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4169 ( .C ( clk ), .D ( new_AGEMA_signal_12196 ), .Q ( new_AGEMA_signal_12197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4177 ( .C ( clk ), .D ( new_AGEMA_signal_12204 ), .Q ( new_AGEMA_signal_12205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4185 ( .C ( clk ), .D ( new_AGEMA_signal_12212 ), .Q ( new_AGEMA_signal_12213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4193 ( .C ( clk ), .D ( new_AGEMA_signal_12220 ), .Q ( new_AGEMA_signal_12221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4215 ( .C ( clk ), .D ( n2183 ), .Q ( new_AGEMA_signal_12243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4221 ( .C ( clk ), .D ( new_AGEMA_signal_1374 ), .Q ( new_AGEMA_signal_12249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4227 ( .C ( clk ), .D ( new_AGEMA_signal_1375 ), .Q ( new_AGEMA_signal_12255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4233 ( .C ( clk ), .D ( new_AGEMA_signal_1376 ), .Q ( new_AGEMA_signal_12261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4239 ( .C ( clk ), .D ( n2196 ), .Q ( new_AGEMA_signal_12267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4245 ( .C ( clk ), .D ( new_AGEMA_signal_1743 ), .Q ( new_AGEMA_signal_12273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4251 ( .C ( clk ), .D ( new_AGEMA_signal_1744 ), .Q ( new_AGEMA_signal_12279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4257 ( .C ( clk ), .D ( new_AGEMA_signal_1745 ), .Q ( new_AGEMA_signal_12285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4263 ( .C ( clk ), .D ( n2238 ), .Q ( new_AGEMA_signal_12291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4269 ( .C ( clk ), .D ( new_AGEMA_signal_1764 ), .Q ( new_AGEMA_signal_12297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4275 ( .C ( clk ), .D ( new_AGEMA_signal_1765 ), .Q ( new_AGEMA_signal_12303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4281 ( .C ( clk ), .D ( new_AGEMA_signal_1766 ), .Q ( new_AGEMA_signal_12309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4287 ( .C ( clk ), .D ( n2249 ), .Q ( new_AGEMA_signal_12315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4293 ( .C ( clk ), .D ( new_AGEMA_signal_2262 ), .Q ( new_AGEMA_signal_12321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4299 ( .C ( clk ), .D ( new_AGEMA_signal_2263 ), .Q ( new_AGEMA_signal_12327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4305 ( .C ( clk ), .D ( new_AGEMA_signal_2264 ), .Q ( new_AGEMA_signal_12333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4311 ( .C ( clk ), .D ( n2273 ), .Q ( new_AGEMA_signal_12339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4317 ( .C ( clk ), .D ( new_AGEMA_signal_2688 ), .Q ( new_AGEMA_signal_12345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4323 ( .C ( clk ), .D ( new_AGEMA_signal_2689 ), .Q ( new_AGEMA_signal_12351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4329 ( .C ( clk ), .D ( new_AGEMA_signal_2690 ), .Q ( new_AGEMA_signal_12357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4353 ( .C ( clk ), .D ( new_AGEMA_signal_12380 ), .Q ( new_AGEMA_signal_12381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4361 ( .C ( clk ), .D ( new_AGEMA_signal_12388 ), .Q ( new_AGEMA_signal_12389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4369 ( .C ( clk ), .D ( new_AGEMA_signal_12396 ), .Q ( new_AGEMA_signal_12397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4377 ( .C ( clk ), .D ( new_AGEMA_signal_12404 ), .Q ( new_AGEMA_signal_12405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4399 ( .C ( clk ), .D ( n2349 ), .Q ( new_AGEMA_signal_12427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4405 ( .C ( clk ), .D ( new_AGEMA_signal_1836 ), .Q ( new_AGEMA_signal_12433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4411 ( .C ( clk ), .D ( new_AGEMA_signal_1837 ), .Q ( new_AGEMA_signal_12439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4417 ( .C ( clk ), .D ( new_AGEMA_signal_1838 ), .Q ( new_AGEMA_signal_12445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4425 ( .C ( clk ), .D ( new_AGEMA_signal_12452 ), .Q ( new_AGEMA_signal_12453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4433 ( .C ( clk ), .D ( new_AGEMA_signal_12460 ), .Q ( new_AGEMA_signal_12461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4441 ( .C ( clk ), .D ( new_AGEMA_signal_12468 ), .Q ( new_AGEMA_signal_12469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4449 ( .C ( clk ), .D ( new_AGEMA_signal_12476 ), .Q ( new_AGEMA_signal_12477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4463 ( .C ( clk ), .D ( n2396 ), .Q ( new_AGEMA_signal_12491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4469 ( .C ( clk ), .D ( new_AGEMA_signal_1869 ), .Q ( new_AGEMA_signal_12497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4475 ( .C ( clk ), .D ( new_AGEMA_signal_1870 ), .Q ( new_AGEMA_signal_12503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4481 ( .C ( clk ), .D ( new_AGEMA_signal_1871 ), .Q ( new_AGEMA_signal_12509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4503 ( .C ( clk ), .D ( n2439 ), .Q ( new_AGEMA_signal_12531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4509 ( .C ( clk ), .D ( new_AGEMA_signal_2367 ), .Q ( new_AGEMA_signal_12537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4515 ( .C ( clk ), .D ( new_AGEMA_signal_2368 ), .Q ( new_AGEMA_signal_12543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4521 ( .C ( clk ), .D ( new_AGEMA_signal_2369 ), .Q ( new_AGEMA_signal_12549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4527 ( .C ( clk ), .D ( n2470 ), .Q ( new_AGEMA_signal_12555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4533 ( .C ( clk ), .D ( new_AGEMA_signal_1899 ), .Q ( new_AGEMA_signal_12561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4539 ( .C ( clk ), .D ( new_AGEMA_signal_1900 ), .Q ( new_AGEMA_signal_12567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4545 ( .C ( clk ), .D ( new_AGEMA_signal_1901 ), .Q ( new_AGEMA_signal_12573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4553 ( .C ( clk ), .D ( new_AGEMA_signal_12580 ), .Q ( new_AGEMA_signal_12581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4561 ( .C ( clk ), .D ( new_AGEMA_signal_12588 ), .Q ( new_AGEMA_signal_12589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4569 ( .C ( clk ), .D ( new_AGEMA_signal_12596 ), .Q ( new_AGEMA_signal_12597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4577 ( .C ( clk ), .D ( new_AGEMA_signal_12604 ), .Q ( new_AGEMA_signal_12605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4585 ( .C ( clk ), .D ( new_AGEMA_signal_12612 ), .Q ( new_AGEMA_signal_12613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4593 ( .C ( clk ), .D ( new_AGEMA_signal_12620 ), .Q ( new_AGEMA_signal_12621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4601 ( .C ( clk ), .D ( new_AGEMA_signal_12628 ), .Q ( new_AGEMA_signal_12629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4609 ( .C ( clk ), .D ( new_AGEMA_signal_12636 ), .Q ( new_AGEMA_signal_12637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4615 ( .C ( clk ), .D ( n2585 ), .Q ( new_AGEMA_signal_12643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4621 ( .C ( clk ), .D ( new_AGEMA_signal_2439 ), .Q ( new_AGEMA_signal_12649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4627 ( .C ( clk ), .D ( new_AGEMA_signal_2440 ), .Q ( new_AGEMA_signal_12655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4633 ( .C ( clk ), .D ( new_AGEMA_signal_2441 ), .Q ( new_AGEMA_signal_12661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4639 ( .C ( clk ), .D ( n2607 ), .Q ( new_AGEMA_signal_12667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4645 ( .C ( clk ), .D ( new_AGEMA_signal_1953 ), .Q ( new_AGEMA_signal_12673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4651 ( .C ( clk ), .D ( new_AGEMA_signal_1954 ), .Q ( new_AGEMA_signal_12679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4657 ( .C ( clk ), .D ( new_AGEMA_signal_1955 ), .Q ( new_AGEMA_signal_12685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4775 ( .C ( clk ), .D ( n2013 ), .Q ( new_AGEMA_signal_12803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4783 ( .C ( clk ), .D ( new_AGEMA_signal_2121 ), .Q ( new_AGEMA_signal_12811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4791 ( .C ( clk ), .D ( new_AGEMA_signal_2122 ), .Q ( new_AGEMA_signal_12819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4799 ( .C ( clk ), .D ( new_AGEMA_signal_2123 ), .Q ( new_AGEMA_signal_12827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4807 ( .C ( clk ), .D ( n2028 ), .Q ( new_AGEMA_signal_12835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4815 ( .C ( clk ), .D ( new_AGEMA_signal_1329 ), .Q ( new_AGEMA_signal_12843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4823 ( .C ( clk ), .D ( new_AGEMA_signal_1330 ), .Q ( new_AGEMA_signal_12851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4831 ( .C ( clk ), .D ( new_AGEMA_signal_1331 ), .Q ( new_AGEMA_signal_12859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4839 ( .C ( clk ), .D ( n2051 ), .Q ( new_AGEMA_signal_12867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4847 ( .C ( clk ), .D ( new_AGEMA_signal_2139 ), .Q ( new_AGEMA_signal_12875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4855 ( .C ( clk ), .D ( new_AGEMA_signal_2140 ), .Q ( new_AGEMA_signal_12883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4863 ( .C ( clk ), .D ( new_AGEMA_signal_2141 ), .Q ( new_AGEMA_signal_12891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4871 ( .C ( clk ), .D ( n2069 ), .Q ( new_AGEMA_signal_12899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4879 ( .C ( clk ), .D ( new_AGEMA_signal_2154 ), .Q ( new_AGEMA_signal_12907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4887 ( .C ( clk ), .D ( new_AGEMA_signal_2155 ), .Q ( new_AGEMA_signal_12915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4895 ( .C ( clk ), .D ( new_AGEMA_signal_2156 ), .Q ( new_AGEMA_signal_12923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4929 ( .C ( clk ), .D ( new_AGEMA_signal_12956 ), .Q ( new_AGEMA_signal_12957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4939 ( .C ( clk ), .D ( new_AGEMA_signal_12966 ), .Q ( new_AGEMA_signal_12967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4949 ( .C ( clk ), .D ( new_AGEMA_signal_12976 ), .Q ( new_AGEMA_signal_12977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4959 ( .C ( clk ), .D ( new_AGEMA_signal_12986 ), .Q ( new_AGEMA_signal_12987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4967 ( .C ( clk ), .D ( n2144 ), .Q ( new_AGEMA_signal_12995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4975 ( .C ( clk ), .D ( new_AGEMA_signal_2205 ), .Q ( new_AGEMA_signal_13003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4983 ( .C ( clk ), .D ( new_AGEMA_signal_2206 ), .Q ( new_AGEMA_signal_13011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4991 ( .C ( clk ), .D ( new_AGEMA_signal_2207 ), .Q ( new_AGEMA_signal_13019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4999 ( .C ( clk ), .D ( n2170 ), .Q ( new_AGEMA_signal_13027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5007 ( .C ( clk ), .D ( new_AGEMA_signal_2211 ), .Q ( new_AGEMA_signal_13035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5015 ( .C ( clk ), .D ( new_AGEMA_signal_2212 ), .Q ( new_AGEMA_signal_13043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5023 ( .C ( clk ), .D ( new_AGEMA_signal_2213 ), .Q ( new_AGEMA_signal_13051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5031 ( .C ( clk ), .D ( n2186 ), .Q ( new_AGEMA_signal_13059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5039 ( .C ( clk ), .D ( new_AGEMA_signal_1368 ), .Q ( new_AGEMA_signal_13067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5047 ( .C ( clk ), .D ( new_AGEMA_signal_1369 ), .Q ( new_AGEMA_signal_13075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5055 ( .C ( clk ), .D ( new_AGEMA_signal_1370 ), .Q ( new_AGEMA_signal_13083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5129 ( .C ( clk ), .D ( new_AGEMA_signal_13156 ), .Q ( new_AGEMA_signal_13157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5139 ( .C ( clk ), .D ( new_AGEMA_signal_13166 ), .Q ( new_AGEMA_signal_13167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5149 ( .C ( clk ), .D ( new_AGEMA_signal_13176 ), .Q ( new_AGEMA_signal_13177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5159 ( .C ( clk ), .D ( new_AGEMA_signal_13186 ), .Q ( new_AGEMA_signal_13187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5167 ( .C ( clk ), .D ( new_AGEMA_signal_10172 ), .Q ( new_AGEMA_signal_13195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5175 ( .C ( clk ), .D ( new_AGEMA_signal_10174 ), .Q ( new_AGEMA_signal_13203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5183 ( .C ( clk ), .D ( new_AGEMA_signal_10176 ), .Q ( new_AGEMA_signal_13211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5191 ( .C ( clk ), .D ( new_AGEMA_signal_10178 ), .Q ( new_AGEMA_signal_13219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C ( clk ), .D ( n2551 ), .Q ( new_AGEMA_signal_13251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C ( clk ), .D ( new_AGEMA_signal_2421 ), .Q ( new_AGEMA_signal_13259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C ( clk ), .D ( new_AGEMA_signal_2422 ), .Q ( new_AGEMA_signal_13267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C ( clk ), .D ( new_AGEMA_signal_2423 ), .Q ( new_AGEMA_signal_13275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5255 ( .C ( clk ), .D ( n2588 ), .Q ( new_AGEMA_signal_13283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5263 ( .C ( clk ), .D ( new_AGEMA_signal_2448 ), .Q ( new_AGEMA_signal_13291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5271 ( .C ( clk ), .D ( new_AGEMA_signal_2449 ), .Q ( new_AGEMA_signal_13299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5279 ( .C ( clk ), .D ( new_AGEMA_signal_2450 ), .Q ( new_AGEMA_signal_13307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5327 ( .C ( clk ), .D ( n2701 ), .Q ( new_AGEMA_signal_13355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5335 ( .C ( clk ), .D ( new_AGEMA_signal_1995 ), .Q ( new_AGEMA_signal_13363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5343 ( .C ( clk ), .D ( new_AGEMA_signal_1996 ), .Q ( new_AGEMA_signal_13371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5351 ( .C ( clk ), .D ( new_AGEMA_signal_1997 ), .Q ( new_AGEMA_signal_13379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5591 ( .C ( clk ), .D ( n2172 ), .Q ( new_AGEMA_signal_13619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5601 ( .C ( clk ), .D ( new_AGEMA_signal_2220 ), .Q ( new_AGEMA_signal_13629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5611 ( .C ( clk ), .D ( new_AGEMA_signal_2221 ), .Q ( new_AGEMA_signal_13639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5621 ( .C ( clk ), .D ( new_AGEMA_signal_2222 ), .Q ( new_AGEMA_signal_13649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6375 ( .C ( clk ), .D ( n2150 ), .Q ( new_AGEMA_signal_14403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6389 ( .C ( clk ), .D ( new_AGEMA_signal_1707 ), .Q ( new_AGEMA_signal_14417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6403 ( .C ( clk ), .D ( new_AGEMA_signal_1708 ), .Q ( new_AGEMA_signal_14431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6417 ( .C ( clk ), .D ( new_AGEMA_signal_1709 ), .Q ( new_AGEMA_signal_14445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6463 ( .C ( clk ), .D ( n2369 ), .Q ( new_AGEMA_signal_14491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6477 ( .C ( clk ), .D ( new_AGEMA_signal_2736 ), .Q ( new_AGEMA_signal_14505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6491 ( .C ( clk ), .D ( new_AGEMA_signal_2737 ), .Q ( new_AGEMA_signal_14519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6505 ( .C ( clk ), .D ( new_AGEMA_signal_2738 ), .Q ( new_AGEMA_signal_14533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6607 ( .C ( clk ), .D ( n2152 ), .Q ( new_AGEMA_signal_14635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6623 ( .C ( clk ), .D ( new_AGEMA_signal_2208 ), .Q ( new_AGEMA_signal_14651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6639 ( .C ( clk ), .D ( new_AGEMA_signal_2209 ), .Q ( new_AGEMA_signal_14667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6655 ( .C ( clk ), .D ( new_AGEMA_signal_2210 ), .Q ( new_AGEMA_signal_14683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6695 ( .C ( clk ), .D ( n2372 ), .Q ( new_AGEMA_signal_14723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6711 ( .C ( clk ), .D ( new_AGEMA_signal_2328 ), .Q ( new_AGEMA_signal_14739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6727 ( .C ( clk ), .D ( new_AGEMA_signal_2329 ), .Q ( new_AGEMA_signal_14755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6743 ( .C ( clk ), .D ( new_AGEMA_signal_2330 ), .Q ( new_AGEMA_signal_14771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6999 ( .C ( clk ), .D ( n2375 ), .Q ( new_AGEMA_signal_15027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7017 ( .C ( clk ), .D ( new_AGEMA_signal_1839 ), .Q ( new_AGEMA_signal_15045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7035 ( .C ( clk ), .D ( new_AGEMA_signal_1840 ), .Q ( new_AGEMA_signal_15063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7053 ( .C ( clk ), .D ( new_AGEMA_signal_1841 ), .Q ( new_AGEMA_signal_15081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7199 ( .C ( clk ), .D ( n2377 ), .Q ( new_AGEMA_signal_15227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7219 ( .C ( clk ), .D ( new_AGEMA_signal_2331 ), .Q ( new_AGEMA_signal_15247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7239 ( .C ( clk ), .D ( new_AGEMA_signal_2332 ), .Q ( new_AGEMA_signal_15267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7259 ( .C ( clk ), .D ( new_AGEMA_signal_2333 ), .Q ( new_AGEMA_signal_15287 ) ) ;

    /* cells in depth 8 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1968 ( .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, n1924}), .b ({new_AGEMA_signal_2048, new_AGEMA_signal_2047, new_AGEMA_signal_2046, n1923}), .clk ( clk ), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, n1936}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1982 ( .a ({new_AGEMA_signal_9626, new_AGEMA_signal_9624, new_AGEMA_signal_9622, new_AGEMA_signal_9620}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, n1927}), .clk ( clk ), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, n1928}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U1994 ( .a ({new_AGEMA_signal_9634, new_AGEMA_signal_9632, new_AGEMA_signal_9630, new_AGEMA_signal_9628}), .b ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, n1929}), .clk ( clk ), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, n1931}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2012 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .b ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, n1938}), .clk ( clk ), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, n1939}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2024 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, n2235}), .b ({new_AGEMA_signal_1529, new_AGEMA_signal_1528, new_AGEMA_signal_1527, n1943}), .clk ( clk ), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n1948}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2032 ( .a ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, n1946}), .b ({new_AGEMA_signal_2066, new_AGEMA_signal_2065, new_AGEMA_signal_2064, n1945}), .clk ( clk ), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, n1947}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2041 ( .a ({new_AGEMA_signal_9650, new_AGEMA_signal_9646, new_AGEMA_signal_9642, new_AGEMA_signal_9638}), .b ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, n1951}), .clk ( clk ), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, n1954}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2049 ( .a ({new_AGEMA_signal_9658, new_AGEMA_signal_9656, new_AGEMA_signal_9654, new_AGEMA_signal_9652}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, n1952}), .clk ( clk ), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, n1953}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2058 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9664, new_AGEMA_signal_9662, new_AGEMA_signal_9660}), .b ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .clk ( clk ), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, n2658}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2065 ( .a ({new_AGEMA_signal_9674, new_AGEMA_signal_9672, new_AGEMA_signal_9670, new_AGEMA_signal_9668}), .b ({new_AGEMA_signal_1547, new_AGEMA_signal_1546, new_AGEMA_signal_1545, n1963}), .clk ( clk ), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n1965}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2078 ( .a ({new_AGEMA_signal_9682, new_AGEMA_signal_9680, new_AGEMA_signal_9678, new_AGEMA_signal_9676}), .b ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, n1968}), .clk ( clk ), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, n1970}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2084 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9688, new_AGEMA_signal_9686, new_AGEMA_signal_9684}), .clk ( clk ), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, n1969}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2093 ( .a ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, n1972}), .b ({new_AGEMA_signal_1565, new_AGEMA_signal_1564, new_AGEMA_signal_1563, n1971}), .clk ( clk ), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, n1978}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2102 ( .a ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, n1974}), .b ({new_AGEMA_signal_9698, new_AGEMA_signal_9696, new_AGEMA_signal_9694, new_AGEMA_signal_9692}), .clk ( clk ), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, n1975}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2107 ( .a ({new_AGEMA_signal_9706, new_AGEMA_signal_9704, new_AGEMA_signal_9702, new_AGEMA_signal_9700}), .b ({new_AGEMA_signal_2102, new_AGEMA_signal_2101, new_AGEMA_signal_2100, n1979}), .clk ( clk ), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, n1980}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2114 ( .a ({new_AGEMA_signal_1574, new_AGEMA_signal_1573, new_AGEMA_signal_1572, n1985}), .b ({new_AGEMA_signal_9714, new_AGEMA_signal_9712, new_AGEMA_signal_9710, new_AGEMA_signal_9708}), .clk ( clk ), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, n1986}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2124 ( .a ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, n1994}), .b ({new_AGEMA_signal_9722, new_AGEMA_signal_9720, new_AGEMA_signal_9718, new_AGEMA_signal_9716}), .clk ( clk ), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n1997}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2137 ( .a ({new_AGEMA_signal_9730, new_AGEMA_signal_9728, new_AGEMA_signal_9726, new_AGEMA_signal_9724}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}), .clk ( clk ), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, n2012}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2145 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, n2006}), .b ({new_AGEMA_signal_2120, new_AGEMA_signal_2119, new_AGEMA_signal_2118, n2005}), .clk ( clk ), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2007}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2161 ( .s ({new_AGEMA_signal_9738, new_AGEMA_signal_9736, new_AGEMA_signal_9734, new_AGEMA_signal_9732}), .b ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, n2020}), .a ({new_AGEMA_signal_9754, new_AGEMA_signal_9750, new_AGEMA_signal_9746, new_AGEMA_signal_9742}), .clk ( clk ), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2021}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2176 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9760, new_AGEMA_signal_9758, new_AGEMA_signal_9756}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, n2031}), .clk ( clk ), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2032}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2185 ( .a ({new_AGEMA_signal_9770, new_AGEMA_signal_9768, new_AGEMA_signal_9766, new_AGEMA_signal_9764}), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, n2040}), .clk ( clk ), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, n2041}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2189 ( .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, n2665}), .b ({new_AGEMA_signal_9778, new_AGEMA_signal_9776, new_AGEMA_signal_9774, new_AGEMA_signal_9772}), .clk ( clk ), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2043}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2194 ( .a ({new_AGEMA_signal_9786, new_AGEMA_signal_9784, new_AGEMA_signal_9782, new_AGEMA_signal_9780}), .b ({new_AGEMA_signal_2138, new_AGEMA_signal_2137, new_AGEMA_signal_2136, n2045}), .clk ( clk ), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, n2046}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2204 ( .s ({new_AGEMA_signal_9738, new_AGEMA_signal_9736, new_AGEMA_signal_9734, new_AGEMA_signal_9732}), .b ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, n2056}), .a ({new_AGEMA_signal_9794, new_AGEMA_signal_9792, new_AGEMA_signal_9790, new_AGEMA_signal_9788}), .clk ( clk ), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2058}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2210 ( .a ({new_AGEMA_signal_9802, new_AGEMA_signal_9800, new_AGEMA_signal_9798, new_AGEMA_signal_9796}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, n2060}), .clk ( clk ), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, n2063}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2218 ( .a ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, n2066}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, n2065}), .clk ( clk ), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2227 ( .a ({new_AGEMA_signal_9810, new_AGEMA_signal_9808, new_AGEMA_signal_9806, new_AGEMA_signal_9804}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, n2074}), .clk ( clk ), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, n2076}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2236 ( .a ({new_AGEMA_signal_9826, new_AGEMA_signal_9822, new_AGEMA_signal_9818, new_AGEMA_signal_9814}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, n2082}), .clk ( clk ), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, n2105}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2241 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9832, new_AGEMA_signal_9830, new_AGEMA_signal_9828}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, n2084}), .clk ( clk ), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, n2099}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2243 ( .a ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, n2085}), .b ({new_AGEMA_signal_9842, new_AGEMA_signal_9840, new_AGEMA_signal_9838, new_AGEMA_signal_9836}), .clk ( clk ), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, n2091}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) U2246 ( .a ({new_AGEMA_signal_9850, new_AGEMA_signal_9848, new_AGEMA_signal_9846, new_AGEMA_signal_9844}), .b ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}), .clk ( clk ), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, n2090}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2253 ( .a ({new_AGEMA_signal_9858, new_AGEMA_signal_9856, new_AGEMA_signal_9854, new_AGEMA_signal_9852}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}), .clk ( clk ), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2093}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2262 ( .a ({new_AGEMA_signal_9866, new_AGEMA_signal_9864, new_AGEMA_signal_9862, new_AGEMA_signal_9860}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}), .clk ( clk ), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, n2102}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2266 ( .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .b ({new_AGEMA_signal_9882, new_AGEMA_signal_9878, new_AGEMA_signal_9874, new_AGEMA_signal_9870}), .clk ( clk ), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, n2106}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2272 ( .a ({new_AGEMA_signal_9890, new_AGEMA_signal_9888, new_AGEMA_signal_9886, new_AGEMA_signal_9884}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, n2114}), .clk ( clk ), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2116}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2282 ( .a ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}), .b ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, n2119}), .clk ( clk ), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, n2120}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2293 ( .a ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, n2130}), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, n2129}), .clk ( clk ), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, n2155}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2296 ( .a ({new_AGEMA_signal_9898, new_AGEMA_signal_9896, new_AGEMA_signal_9894, new_AGEMA_signal_9892}), .b ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, n2131}), .clk ( clk ), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2299 ( .a ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, n2133}), .b ({new_AGEMA_signal_9906, new_AGEMA_signal_9904, new_AGEMA_signal_9902, new_AGEMA_signal_9900}), .clk ( clk ), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2134}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2303 ( .a ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, n2137}), .b ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, n2136}), .clk ( clk ), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, n2143}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2308 ( .a ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, n2139}), .b ({new_AGEMA_signal_9922, new_AGEMA_signal_9918, new_AGEMA_signal_9914, new_AGEMA_signal_9910}), .clk ( clk ), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, n2140}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2324 ( .a ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, n2157}), .b ({new_AGEMA_signal_9930, new_AGEMA_signal_9928, new_AGEMA_signal_9926, new_AGEMA_signal_9924}), .clk ( clk ), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, n2159}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2326 ( .a ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, n2160}), .b ({new_AGEMA_signal_9938, new_AGEMA_signal_9936, new_AGEMA_signal_9934, new_AGEMA_signal_9932}), .clk ( clk ), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, n2161}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2330 ( .a ({new_AGEMA_signal_9650, new_AGEMA_signal_9646, new_AGEMA_signal_9642, new_AGEMA_signal_9638}), .b ({new_AGEMA_signal_1727, new_AGEMA_signal_1726, new_AGEMA_signal_1725, n2163}), .clk ( clk ), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, n2164}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2345 ( .a ({new_AGEMA_signal_9946, new_AGEMA_signal_9944, new_AGEMA_signal_9942, new_AGEMA_signal_9940}), .b ({new_AGEMA_signal_2228, new_AGEMA_signal_2227, new_AGEMA_signal_2226, n2177}), .clk ( clk ), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, n2179}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2359 ( .a ({new_AGEMA_signal_9962, new_AGEMA_signal_9958, new_AGEMA_signal_9954, new_AGEMA_signal_9950}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, n2191}), .clk ( clk ), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2192}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2370 ( .a ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, n2201}), .b ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, n2200}), .clk ( clk ), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, n2203}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2382 ( .a ({new_AGEMA_signal_2246, new_AGEMA_signal_2245, new_AGEMA_signal_2244, n2217}), .b ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, n2216}), .clk ( clk ), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, n2224}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2388 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, n2222}), .b ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, n2221}), .clk ( clk ), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2223}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2392 ( .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .b ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, n2226}), .clk ( clk ), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, n2229}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2399 ( .a ({new_AGEMA_signal_9658, new_AGEMA_signal_9656, new_AGEMA_signal_9654, new_AGEMA_signal_9652}), .b ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, n2233}), .clk ( clk ), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, n2234}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2410 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9664, new_AGEMA_signal_9662, new_AGEMA_signal_9660}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, n2244}), .clk ( clk ), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, n2246}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2418 ( .a ({new_AGEMA_signal_9970, new_AGEMA_signal_9968, new_AGEMA_signal_9966, new_AGEMA_signal_9964}), .b ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, n2253}), .clk ( clk ), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2254}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2425 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9976, new_AGEMA_signal_9974, new_AGEMA_signal_9972}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, n2260}), .clk ( clk ), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, n2263}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2434 ( .a ({new_AGEMA_signal_9986, new_AGEMA_signal_9984, new_AGEMA_signal_9982, new_AGEMA_signal_9980}), .b ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, n2265}), .clk ( clk ), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, n2267}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2438 ( .a ({new_AGEMA_signal_9658, new_AGEMA_signal_9656, new_AGEMA_signal_9654, new_AGEMA_signal_9652}), .b ({new_AGEMA_signal_1790, new_AGEMA_signal_1789, new_AGEMA_signal_1788, n2269}), .clk ( clk ), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, n2270}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2445 ( .a ({new_AGEMA_signal_9994, new_AGEMA_signal_9992, new_AGEMA_signal_9990, new_AGEMA_signal_9988}), .b ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, n2277}), .clk ( clk ), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, n2279}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2450 ( .a ({new_AGEMA_signal_9754, new_AGEMA_signal_9750, new_AGEMA_signal_9746, new_AGEMA_signal_9742}), .b ({new_AGEMA_signal_1799, new_AGEMA_signal_1798, new_AGEMA_signal_1797, n2282}), .clk ( clk ), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2283}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2453 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9832, new_AGEMA_signal_9830, new_AGEMA_signal_9828}), .b ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, n2284}), .clk ( clk ), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, n2285}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2457 ( .a ({new_AGEMA_signal_9650, new_AGEMA_signal_9646, new_AGEMA_signal_9642, new_AGEMA_signal_9638}), .b ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, n2459}), .clk ( clk ), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2460 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9664, new_AGEMA_signal_9662, new_AGEMA_signal_9660}), .b ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, n2288}), .clk ( clk ), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2289}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2463 ( .a ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}), .b ({new_AGEMA_signal_10002, new_AGEMA_signal_10000, new_AGEMA_signal_9998, new_AGEMA_signal_9996}), .clk ( clk ), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, n2297}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2465 ( .a ({new_AGEMA_signal_10010, new_AGEMA_signal_10008, new_AGEMA_signal_10006, new_AGEMA_signal_10004}), .b ({new_AGEMA_signal_2192, new_AGEMA_signal_2191, new_AGEMA_signal_2190, n2291}), .clk ( clk ), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2292}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2473 ( .a ({new_AGEMA_signal_10018, new_AGEMA_signal_10016, new_AGEMA_signal_10014, new_AGEMA_signal_10012}), .b ({new_AGEMA_signal_2300, new_AGEMA_signal_2299, new_AGEMA_signal_2298, n2300}), .clk ( clk ), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, n2301}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2483 ( .a ({new_AGEMA_signal_10026, new_AGEMA_signal_10024, new_AGEMA_signal_10022, new_AGEMA_signal_10020}), .b ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, n2314}), .clk ( clk ), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2321}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2487 ( .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, n2319}), .b ({new_AGEMA_signal_10034, new_AGEMA_signal_10032, new_AGEMA_signal_10030, new_AGEMA_signal_10028}), .clk ( clk ), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, n2320}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2493 ( .a ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, n2326}), .b ({new_AGEMA_signal_10042, new_AGEMA_signal_10040, new_AGEMA_signal_10038, new_AGEMA_signal_10036}), .clk ( clk ), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, n2334}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2497 ( .a ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, n2329}), .b ({new_AGEMA_signal_9754, new_AGEMA_signal_9750, new_AGEMA_signal_9746, new_AGEMA_signal_9742}), .clk ( clk ), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, n2332}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2498 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10048, new_AGEMA_signal_10046, new_AGEMA_signal_10044}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, n2330}), .clk ( clk ), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2331}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2502 ( .a ({new_AGEMA_signal_10058, new_AGEMA_signal_10056, new_AGEMA_signal_10054, new_AGEMA_signal_10052}), .b ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, n2335}), .clk ( clk ), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, n2336}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2508 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, n2341}), .b ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, n2340}), .clk ( clk ), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2342}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2519 ( .a ({new_AGEMA_signal_1844, new_AGEMA_signal_1843, new_AGEMA_signal_1842, n2352}), .b ({new_AGEMA_signal_10066, new_AGEMA_signal_10064, new_AGEMA_signal_10062, new_AGEMA_signal_10060}), .clk ( clk ), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, n2367}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2523 ( .a ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, n2354}), .b ({new_AGEMA_signal_10074, new_AGEMA_signal_10072, new_AGEMA_signal_10070, new_AGEMA_signal_10068}), .clk ( clk ), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, n2358}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2547 ( .a ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, n2385}), .b ({new_AGEMA_signal_1862, new_AGEMA_signal_1861, new_AGEMA_signal_1860, n2384}), .clk ( clk ), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2387}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2555 ( .a ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, n2391}), .b ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, n2390}), .clk ( clk ), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2392}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2566 ( .a ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, n2403}), .b ({new_AGEMA_signal_10082, new_AGEMA_signal_10080, new_AGEMA_signal_10078, new_AGEMA_signal_10076}), .clk ( clk ), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2404}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2570 ( .a ({new_AGEMA_signal_9802, new_AGEMA_signal_9800, new_AGEMA_signal_9798, new_AGEMA_signal_9796}), .b ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, n2408}), .clk ( clk ), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2409}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2575 ( .a ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, n2413}), .clk ( clk ), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, n2414}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2578 ( .a ({new_AGEMA_signal_10090, new_AGEMA_signal_10088, new_AGEMA_signal_10086, new_AGEMA_signal_10084}), .b ({new_AGEMA_signal_1880, new_AGEMA_signal_1879, new_AGEMA_signal_1878, n2416}), .clk ( clk ), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, n2418}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2589 ( .a ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}), .b ({new_AGEMA_signal_10098, new_AGEMA_signal_10096, new_AGEMA_signal_10094, new_AGEMA_signal_10092}), .clk ( clk ), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, n2432}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2592 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10116, new_AGEMA_signal_10110, new_AGEMA_signal_10104}), .b ({new_AGEMA_signal_1889, new_AGEMA_signal_1888, new_AGEMA_signal_1887, n2434}), .clk ( clk ), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, n2435}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2601 ( .a ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, n2445}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, n2444}), .clk ( clk ), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2449}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2603 ( .a ({new_AGEMA_signal_10026, new_AGEMA_signal_10024, new_AGEMA_signal_10022, new_AGEMA_signal_10020}), .b ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, n2447}), .clk ( clk ), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, n2448}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2609 ( .a ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, n2454}), .b ({new_AGEMA_signal_10130, new_AGEMA_signal_10128, new_AGEMA_signal_10126, new_AGEMA_signal_10124}), .clk ( clk ), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2455}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2612 ( .a ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, n2458}), .clk ( clk ), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, n2460}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2618 ( .a ({new_AGEMA_signal_10010, new_AGEMA_signal_10008, new_AGEMA_signal_10006, new_AGEMA_signal_10004}), .b ({new_AGEMA_signal_1898, new_AGEMA_signal_1897, new_AGEMA_signal_1896, n2465}), .clk ( clk ), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2466}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2629 ( .a ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, n2476}), .b ({new_AGEMA_signal_10138, new_AGEMA_signal_10136, new_AGEMA_signal_10134, new_AGEMA_signal_10132}), .clk ( clk ), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, n2477}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2634 ( .a ({new_AGEMA_signal_9794, new_AGEMA_signal_9792, new_AGEMA_signal_9790, new_AGEMA_signal_9788}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, n2481}), .clk ( clk ), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2482}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2640 ( .a ({new_AGEMA_signal_10146, new_AGEMA_signal_10144, new_AGEMA_signal_10142, new_AGEMA_signal_10140}), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, n2486}), .clk ( clk ), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, n2490}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2648 ( .a ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, n2495}), .b ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, n2494}), .clk ( clk ), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2496}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2654 ( .a ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, n2504}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, n2503}), .clk ( clk ), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, n2507}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2664 ( .a ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, n2518}), .b ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, n2517}), .clk ( clk ), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, n2525}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2669 ( .a ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, n2523}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, n2522}), .clk ( clk ), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, n2524}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2676 ( .a ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, n2532}), .b ({new_AGEMA_signal_10162, new_AGEMA_signal_10158, new_AGEMA_signal_10154, new_AGEMA_signal_10150}), .clk ( clk ), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, n2537}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2678 ( .a ({new_AGEMA_signal_9802, new_AGEMA_signal_9800, new_AGEMA_signal_9798, new_AGEMA_signal_9796}), .b ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, n2534}), .clk ( clk ), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, n2536}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2684 ( .a ({new_AGEMA_signal_10170, new_AGEMA_signal_10168, new_AGEMA_signal_10166, new_AGEMA_signal_10164}), .b ({new_AGEMA_signal_1934, new_AGEMA_signal_1933, new_AGEMA_signal_1932, n2546}), .clk ( clk ), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, n2547}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2693 ( .a ({new_AGEMA_signal_10178, new_AGEMA_signal_10176, new_AGEMA_signal_10174, new_AGEMA_signal_10172}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, n2556}), .clk ( clk ), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2557}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2699 ( .a ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}), .b ({new_AGEMA_signal_10186, new_AGEMA_signal_10184, new_AGEMA_signal_10182, new_AGEMA_signal_10180}), .clk ( clk ), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, n2565}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2704 ( .a ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, n2574}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, n2573}), .clk ( clk ), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, n2591}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2709 ( .a ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, n2579}), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, n2578}), .clk ( clk ), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, n2580}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2727 ( .a ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, n2601}), .b ({new_AGEMA_signal_10202, new_AGEMA_signal_10198, new_AGEMA_signal_10194, new_AGEMA_signal_10190}), .clk ( clk ), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2602}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2738 ( .a ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, n2618}), .b ({new_AGEMA_signal_10210, new_AGEMA_signal_10208, new_AGEMA_signal_10206, new_AGEMA_signal_10204}), .clk ( clk ), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, n2619}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2744 ( .a ({new_AGEMA_signal_9842, new_AGEMA_signal_9840, new_AGEMA_signal_9838, new_AGEMA_signal_9836}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, n2626}), .clk ( clk ), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, n2628}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2753 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, n2644}), .b ({new_AGEMA_signal_9898, new_AGEMA_signal_9896, new_AGEMA_signal_9894, new_AGEMA_signal_9892}), .clk ( clk ), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, n2649}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2755 ( .a ({new_AGEMA_signal_10218, new_AGEMA_signal_10216, new_AGEMA_signal_10214, new_AGEMA_signal_10212}), .b ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, n2646}), .clk ( clk ), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, n2648}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2765 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9664, new_AGEMA_signal_9662, new_AGEMA_signal_9660}), .b ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, n2663}), .clk ( clk ), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2664}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2771 ( .a ({new_AGEMA_signal_1988, new_AGEMA_signal_1987, new_AGEMA_signal_1986, n2675}), .b ({new_AGEMA_signal_10226, new_AGEMA_signal_10224, new_AGEMA_signal_10222, new_AGEMA_signal_10220}), .clk ( clk ), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, n2681}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2773 ( .a ({new_AGEMA_signal_9930, new_AGEMA_signal_9928, new_AGEMA_signal_9926, new_AGEMA_signal_9924}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, n2678}), .clk ( clk ), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2680}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2776 ( .a ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, n2684}), .b ({new_AGEMA_signal_10234, new_AGEMA_signal_10232, new_AGEMA_signal_10230, new_AGEMA_signal_10228}), .clk ( clk ), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, n2685}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2778 ( .a ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, n2687}), .b ({new_AGEMA_signal_10170, new_AGEMA_signal_10168, new_AGEMA_signal_10166, new_AGEMA_signal_10164}), .clk ( clk ), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, n2698}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2779 ( .a ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, n2689}), .b ({new_AGEMA_signal_10178, new_AGEMA_signal_10176, new_AGEMA_signal_10174, new_AGEMA_signal_10172}), .clk ( clk ), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2692}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2793 ( .a ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, n2715}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10240, new_AGEMA_signal_10238, new_AGEMA_signal_10236}), .clk ( clk ), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, n2716}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2800 ( .a ({new_AGEMA_signal_2006, new_AGEMA_signal_2005, new_AGEMA_signal_2004, n2727}), .b ({new_AGEMA_signal_10250, new_AGEMA_signal_10248, new_AGEMA_signal_10246, new_AGEMA_signal_10244}), .clk ( clk ), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, n2728}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2804 ( .a ({new_AGEMA_signal_10258, new_AGEMA_signal_10256, new_AGEMA_signal_10254, new_AGEMA_signal_10252}), .b ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, n2733}), .clk ( clk ), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, n2735}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2808 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9712, new_AGEMA_signal_9710, new_AGEMA_signal_9708}), .b ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, n2740}), .clk ( clk ), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2743}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2813 ( .a ({new_AGEMA_signal_10274, new_AGEMA_signal_10270, new_AGEMA_signal_10266, new_AGEMA_signal_10262}), .b ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, new_AGEMA_signal_2013, n2749}), .clk ( clk ), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2751}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2817 ( .a ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, n2757}), .b ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, n2756}), .clk ( clk ), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, n2758}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2820 ( .a ({new_AGEMA_signal_10282, new_AGEMA_signal_10280, new_AGEMA_signal_10278, new_AGEMA_signal_10276}), .b ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, n2762}), .clk ( clk ), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, n2764}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2827 ( .a ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, n2776}), .b ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, n2775}), .clk ( clk ), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, n2800}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2831 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10288, new_AGEMA_signal_10286, new_AGEMA_signal_10284}), .b ({new_AGEMA_signal_2024, new_AGEMA_signal_2023, new_AGEMA_signal_2022, n2783}), .clk ( clk ), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2788}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2837 ( .a ({new_AGEMA_signal_10306, new_AGEMA_signal_10302, new_AGEMA_signal_10298, new_AGEMA_signal_10294}), .b ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, n2795}), .clk ( clk ), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, n2797}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2846 ( .a ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, n2814}), .b ({new_AGEMA_signal_9738, new_AGEMA_signal_9736, new_AGEMA_signal_9734, new_AGEMA_signal_9732}), .clk ( clk ), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, n2822}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2849 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10312, new_AGEMA_signal_10310, new_AGEMA_signal_10308}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, n2819}), .clk ( clk ), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, n2821}) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C ( clk ), .D ( new_AGEMA_signal_10317 ), .Q ( new_AGEMA_signal_10318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C ( clk ), .D ( new_AGEMA_signal_10321 ), .Q ( new_AGEMA_signal_10322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C ( clk ), .D ( new_AGEMA_signal_10325 ), .Q ( new_AGEMA_signal_10326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C ( clk ), .D ( new_AGEMA_signal_10329 ), .Q ( new_AGEMA_signal_10330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C ( clk ), .D ( new_AGEMA_signal_10333 ), .Q ( new_AGEMA_signal_10334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C ( clk ), .D ( new_AGEMA_signal_10337 ), .Q ( new_AGEMA_signal_10338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C ( clk ), .D ( new_AGEMA_signal_10341 ), .Q ( new_AGEMA_signal_10342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C ( clk ), .D ( new_AGEMA_signal_10345 ), .Q ( new_AGEMA_signal_10346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C ( clk ), .D ( new_AGEMA_signal_10347 ), .Q ( new_AGEMA_signal_10348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C ( clk ), .D ( new_AGEMA_signal_10349 ), .Q ( new_AGEMA_signal_10350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C ( clk ), .D ( new_AGEMA_signal_10351 ), .Q ( new_AGEMA_signal_10352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C ( clk ), .D ( new_AGEMA_signal_10353 ), .Q ( new_AGEMA_signal_10354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C ( clk ), .D ( new_AGEMA_signal_10355 ), .Q ( new_AGEMA_signal_10356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C ( clk ), .D ( new_AGEMA_signal_10357 ), .Q ( new_AGEMA_signal_10358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C ( clk ), .D ( new_AGEMA_signal_10359 ), .Q ( new_AGEMA_signal_10360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C ( clk ), .D ( new_AGEMA_signal_10361 ), .Q ( new_AGEMA_signal_10362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C ( clk ), .D ( new_AGEMA_signal_10365 ), .Q ( new_AGEMA_signal_10366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C ( clk ), .D ( new_AGEMA_signal_10369 ), .Q ( new_AGEMA_signal_10370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C ( clk ), .D ( new_AGEMA_signal_10373 ), .Q ( new_AGEMA_signal_10374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C ( clk ), .D ( new_AGEMA_signal_10377 ), .Q ( new_AGEMA_signal_10378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C ( clk ), .D ( new_AGEMA_signal_10379 ), .Q ( new_AGEMA_signal_10380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C ( clk ), .D ( new_AGEMA_signal_10381 ), .Q ( new_AGEMA_signal_10382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C ( clk ), .D ( new_AGEMA_signal_10383 ), .Q ( new_AGEMA_signal_10384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C ( clk ), .D ( new_AGEMA_signal_10385 ), .Q ( new_AGEMA_signal_10386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C ( clk ), .D ( new_AGEMA_signal_10389 ), .Q ( new_AGEMA_signal_10390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C ( clk ), .D ( new_AGEMA_signal_10393 ), .Q ( new_AGEMA_signal_10394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C ( clk ), .D ( new_AGEMA_signal_10397 ), .Q ( new_AGEMA_signal_10398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C ( clk ), .D ( new_AGEMA_signal_10401 ), .Q ( new_AGEMA_signal_10402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C ( clk ), .D ( new_AGEMA_signal_10403 ), .Q ( new_AGEMA_signal_10404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C ( clk ), .D ( new_AGEMA_signal_10405 ), .Q ( new_AGEMA_signal_10406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C ( clk ), .D ( new_AGEMA_signal_10407 ), .Q ( new_AGEMA_signal_10408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C ( clk ), .D ( new_AGEMA_signal_10409 ), .Q ( new_AGEMA_signal_10410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C ( clk ), .D ( new_AGEMA_signal_10413 ), .Q ( new_AGEMA_signal_10414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C ( clk ), .D ( new_AGEMA_signal_10417 ), .Q ( new_AGEMA_signal_10418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C ( clk ), .D ( new_AGEMA_signal_10421 ), .Q ( new_AGEMA_signal_10422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C ( clk ), .D ( new_AGEMA_signal_10425 ), .Q ( new_AGEMA_signal_10426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C ( clk ), .D ( new_AGEMA_signal_10429 ), .Q ( new_AGEMA_signal_10430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C ( clk ), .D ( new_AGEMA_signal_10433 ), .Q ( new_AGEMA_signal_10434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C ( clk ), .D ( new_AGEMA_signal_10437 ), .Q ( new_AGEMA_signal_10438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C ( clk ), .D ( new_AGEMA_signal_10441 ), .Q ( new_AGEMA_signal_10442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C ( clk ), .D ( new_AGEMA_signal_10443 ), .Q ( new_AGEMA_signal_10444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C ( clk ), .D ( new_AGEMA_signal_10445 ), .Q ( new_AGEMA_signal_10446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C ( clk ), .D ( new_AGEMA_signal_10447 ), .Q ( new_AGEMA_signal_10448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C ( clk ), .D ( new_AGEMA_signal_10449 ), .Q ( new_AGEMA_signal_10450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C ( clk ), .D ( new_AGEMA_signal_10451 ), .Q ( new_AGEMA_signal_10452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C ( clk ), .D ( new_AGEMA_signal_10453 ), .Q ( new_AGEMA_signal_10454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C ( clk ), .D ( new_AGEMA_signal_10455 ), .Q ( new_AGEMA_signal_10456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C ( clk ), .D ( new_AGEMA_signal_10457 ), .Q ( new_AGEMA_signal_10458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C ( clk ), .D ( new_AGEMA_signal_10459 ), .Q ( new_AGEMA_signal_10460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C ( clk ), .D ( new_AGEMA_signal_10461 ), .Q ( new_AGEMA_signal_10462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C ( clk ), .D ( new_AGEMA_signal_10463 ), .Q ( new_AGEMA_signal_10464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C ( clk ), .D ( new_AGEMA_signal_10465 ), .Q ( new_AGEMA_signal_10466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C ( clk ), .D ( new_AGEMA_signal_10467 ), .Q ( new_AGEMA_signal_10468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C ( clk ), .D ( new_AGEMA_signal_10469 ), .Q ( new_AGEMA_signal_10470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C ( clk ), .D ( new_AGEMA_signal_10471 ), .Q ( new_AGEMA_signal_10472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C ( clk ), .D ( new_AGEMA_signal_10473 ), .Q ( new_AGEMA_signal_10474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C ( clk ), .D ( new_AGEMA_signal_10477 ), .Q ( new_AGEMA_signal_10478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C ( clk ), .D ( new_AGEMA_signal_10481 ), .Q ( new_AGEMA_signal_10482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C ( clk ), .D ( new_AGEMA_signal_10485 ), .Q ( new_AGEMA_signal_10486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C ( clk ), .D ( new_AGEMA_signal_10489 ), .Q ( new_AGEMA_signal_10490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C ( clk ), .D ( new_AGEMA_signal_10493 ), .Q ( new_AGEMA_signal_10494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C ( clk ), .D ( new_AGEMA_signal_10497 ), .Q ( new_AGEMA_signal_10498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C ( clk ), .D ( new_AGEMA_signal_10501 ), .Q ( new_AGEMA_signal_10502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C ( clk ), .D ( new_AGEMA_signal_10505 ), .Q ( new_AGEMA_signal_10506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C ( clk ), .D ( new_AGEMA_signal_10509 ), .Q ( new_AGEMA_signal_10510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C ( clk ), .D ( new_AGEMA_signal_10513 ), .Q ( new_AGEMA_signal_10514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C ( clk ), .D ( new_AGEMA_signal_10517 ), .Q ( new_AGEMA_signal_10518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C ( clk ), .D ( new_AGEMA_signal_10521 ), .Q ( new_AGEMA_signal_10522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C ( clk ), .D ( new_AGEMA_signal_10523 ), .Q ( new_AGEMA_signal_10524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C ( clk ), .D ( new_AGEMA_signal_10525 ), .Q ( new_AGEMA_signal_10526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C ( clk ), .D ( new_AGEMA_signal_10527 ), .Q ( new_AGEMA_signal_10528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C ( clk ), .D ( new_AGEMA_signal_10529 ), .Q ( new_AGEMA_signal_10530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C ( clk ), .D ( new_AGEMA_signal_10531 ), .Q ( new_AGEMA_signal_10532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C ( clk ), .D ( new_AGEMA_signal_10533 ), .Q ( new_AGEMA_signal_10534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C ( clk ), .D ( new_AGEMA_signal_10535 ), .Q ( new_AGEMA_signal_10536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C ( clk ), .D ( new_AGEMA_signal_10537 ), .Q ( new_AGEMA_signal_10538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C ( clk ), .D ( new_AGEMA_signal_10539 ), .Q ( new_AGEMA_signal_10540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C ( clk ), .D ( new_AGEMA_signal_10541 ), .Q ( new_AGEMA_signal_10542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C ( clk ), .D ( new_AGEMA_signal_10543 ), .Q ( new_AGEMA_signal_10544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C ( clk ), .D ( new_AGEMA_signal_10545 ), .Q ( new_AGEMA_signal_10546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C ( clk ), .D ( new_AGEMA_signal_10549 ), .Q ( new_AGEMA_signal_10550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C ( clk ), .D ( new_AGEMA_signal_10553 ), .Q ( new_AGEMA_signal_10554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C ( clk ), .D ( new_AGEMA_signal_10557 ), .Q ( new_AGEMA_signal_10558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C ( clk ), .D ( new_AGEMA_signal_10561 ), .Q ( new_AGEMA_signal_10562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C ( clk ), .D ( new_AGEMA_signal_10563 ), .Q ( new_AGEMA_signal_10564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C ( clk ), .D ( new_AGEMA_signal_10565 ), .Q ( new_AGEMA_signal_10566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C ( clk ), .D ( new_AGEMA_signal_10567 ), .Q ( new_AGEMA_signal_10568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C ( clk ), .D ( new_AGEMA_signal_10569 ), .Q ( new_AGEMA_signal_10570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C ( clk ), .D ( new_AGEMA_signal_10573 ), .Q ( new_AGEMA_signal_10574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C ( clk ), .D ( new_AGEMA_signal_10577 ), .Q ( new_AGEMA_signal_10578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C ( clk ), .D ( new_AGEMA_signal_10581 ), .Q ( new_AGEMA_signal_10582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C ( clk ), .D ( new_AGEMA_signal_10585 ), .Q ( new_AGEMA_signal_10586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C ( clk ), .D ( new_AGEMA_signal_10591 ), .Q ( new_AGEMA_signal_10592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C ( clk ), .D ( new_AGEMA_signal_10597 ), .Q ( new_AGEMA_signal_10598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C ( clk ), .D ( new_AGEMA_signal_10603 ), .Q ( new_AGEMA_signal_10604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C ( clk ), .D ( new_AGEMA_signal_10609 ), .Q ( new_AGEMA_signal_10610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C ( clk ), .D ( new_AGEMA_signal_10613 ), .Q ( new_AGEMA_signal_10614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C ( clk ), .D ( new_AGEMA_signal_10617 ), .Q ( new_AGEMA_signal_10618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C ( clk ), .D ( new_AGEMA_signal_10621 ), .Q ( new_AGEMA_signal_10622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C ( clk ), .D ( new_AGEMA_signal_10625 ), .Q ( new_AGEMA_signal_10626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C ( clk ), .D ( new_AGEMA_signal_10629 ), .Q ( new_AGEMA_signal_10630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C ( clk ), .D ( new_AGEMA_signal_10633 ), .Q ( new_AGEMA_signal_10634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C ( clk ), .D ( new_AGEMA_signal_10637 ), .Q ( new_AGEMA_signal_10638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C ( clk ), .D ( new_AGEMA_signal_10641 ), .Q ( new_AGEMA_signal_10642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C ( clk ), .D ( new_AGEMA_signal_10643 ), .Q ( new_AGEMA_signal_10644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C ( clk ), .D ( new_AGEMA_signal_10645 ), .Q ( new_AGEMA_signal_10646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C ( clk ), .D ( new_AGEMA_signal_10647 ), .Q ( new_AGEMA_signal_10648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C ( clk ), .D ( new_AGEMA_signal_10649 ), .Q ( new_AGEMA_signal_10650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C ( clk ), .D ( new_AGEMA_signal_10651 ), .Q ( new_AGEMA_signal_10652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C ( clk ), .D ( new_AGEMA_signal_10653 ), .Q ( new_AGEMA_signal_10654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C ( clk ), .D ( new_AGEMA_signal_10655 ), .Q ( new_AGEMA_signal_10656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C ( clk ), .D ( new_AGEMA_signal_10657 ), .Q ( new_AGEMA_signal_10658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C ( clk ), .D ( new_AGEMA_signal_10659 ), .Q ( new_AGEMA_signal_10660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C ( clk ), .D ( new_AGEMA_signal_10661 ), .Q ( new_AGEMA_signal_10662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C ( clk ), .D ( new_AGEMA_signal_10663 ), .Q ( new_AGEMA_signal_10664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C ( clk ), .D ( new_AGEMA_signal_10665 ), .Q ( new_AGEMA_signal_10666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C ( clk ), .D ( new_AGEMA_signal_10667 ), .Q ( new_AGEMA_signal_10668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C ( clk ), .D ( new_AGEMA_signal_10669 ), .Q ( new_AGEMA_signal_10670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C ( clk ), .D ( new_AGEMA_signal_10671 ), .Q ( new_AGEMA_signal_10672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C ( clk ), .D ( new_AGEMA_signal_10673 ), .Q ( new_AGEMA_signal_10674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C ( clk ), .D ( new_AGEMA_signal_10677 ), .Q ( new_AGEMA_signal_10678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C ( clk ), .D ( new_AGEMA_signal_10681 ), .Q ( new_AGEMA_signal_10682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C ( clk ), .D ( new_AGEMA_signal_10685 ), .Q ( new_AGEMA_signal_10686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C ( clk ), .D ( new_AGEMA_signal_10689 ), .Q ( new_AGEMA_signal_10690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C ( clk ), .D ( new_AGEMA_signal_10695 ), .Q ( new_AGEMA_signal_10696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C ( clk ), .D ( new_AGEMA_signal_10701 ), .Q ( new_AGEMA_signal_10702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C ( clk ), .D ( new_AGEMA_signal_10707 ), .Q ( new_AGEMA_signal_10708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C ( clk ), .D ( new_AGEMA_signal_10713 ), .Q ( new_AGEMA_signal_10714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C ( clk ), .D ( new_AGEMA_signal_10717 ), .Q ( new_AGEMA_signal_10718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C ( clk ), .D ( new_AGEMA_signal_10721 ), .Q ( new_AGEMA_signal_10722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C ( clk ), .D ( new_AGEMA_signal_10725 ), .Q ( new_AGEMA_signal_10726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C ( clk ), .D ( new_AGEMA_signal_10729 ), .Q ( new_AGEMA_signal_10730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C ( clk ), .D ( new_AGEMA_signal_10731 ), .Q ( new_AGEMA_signal_10732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C ( clk ), .D ( new_AGEMA_signal_10733 ), .Q ( new_AGEMA_signal_10734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C ( clk ), .D ( new_AGEMA_signal_10735 ), .Q ( new_AGEMA_signal_10736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C ( clk ), .D ( new_AGEMA_signal_10737 ), .Q ( new_AGEMA_signal_10738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C ( clk ), .D ( new_AGEMA_signal_10739 ), .Q ( new_AGEMA_signal_10740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C ( clk ), .D ( new_AGEMA_signal_10741 ), .Q ( new_AGEMA_signal_10742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C ( clk ), .D ( new_AGEMA_signal_10743 ), .Q ( new_AGEMA_signal_10744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C ( clk ), .D ( new_AGEMA_signal_10745 ), .Q ( new_AGEMA_signal_10746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C ( clk ), .D ( new_AGEMA_signal_10747 ), .Q ( new_AGEMA_signal_10748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C ( clk ), .D ( new_AGEMA_signal_10749 ), .Q ( new_AGEMA_signal_10750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C ( clk ), .D ( new_AGEMA_signal_10751 ), .Q ( new_AGEMA_signal_10752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C ( clk ), .D ( new_AGEMA_signal_10753 ), .Q ( new_AGEMA_signal_10754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C ( clk ), .D ( new_AGEMA_signal_10757 ), .Q ( new_AGEMA_signal_10758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C ( clk ), .D ( new_AGEMA_signal_10761 ), .Q ( new_AGEMA_signal_10762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C ( clk ), .D ( new_AGEMA_signal_10765 ), .Q ( new_AGEMA_signal_10766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C ( clk ), .D ( new_AGEMA_signal_10769 ), .Q ( new_AGEMA_signal_10770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C ( clk ), .D ( new_AGEMA_signal_10771 ), .Q ( new_AGEMA_signal_10772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C ( clk ), .D ( new_AGEMA_signal_10773 ), .Q ( new_AGEMA_signal_10774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C ( clk ), .D ( new_AGEMA_signal_10775 ), .Q ( new_AGEMA_signal_10776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C ( clk ), .D ( new_AGEMA_signal_10777 ), .Q ( new_AGEMA_signal_10778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C ( clk ), .D ( new_AGEMA_signal_10779 ), .Q ( new_AGEMA_signal_10780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C ( clk ), .D ( new_AGEMA_signal_10781 ), .Q ( new_AGEMA_signal_10782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C ( clk ), .D ( new_AGEMA_signal_10783 ), .Q ( new_AGEMA_signal_10784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C ( clk ), .D ( new_AGEMA_signal_10785 ), .Q ( new_AGEMA_signal_10786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C ( clk ), .D ( new_AGEMA_signal_10789 ), .Q ( new_AGEMA_signal_10790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C ( clk ), .D ( new_AGEMA_signal_10793 ), .Q ( new_AGEMA_signal_10794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C ( clk ), .D ( new_AGEMA_signal_10797 ), .Q ( new_AGEMA_signal_10798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C ( clk ), .D ( new_AGEMA_signal_10801 ), .Q ( new_AGEMA_signal_10802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C ( clk ), .D ( new_AGEMA_signal_10805 ), .Q ( new_AGEMA_signal_10806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C ( clk ), .D ( new_AGEMA_signal_10809 ), .Q ( new_AGEMA_signal_10810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C ( clk ), .D ( new_AGEMA_signal_10813 ), .Q ( new_AGEMA_signal_10814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C ( clk ), .D ( new_AGEMA_signal_10817 ), .Q ( new_AGEMA_signal_10818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C ( clk ), .D ( new_AGEMA_signal_10821 ), .Q ( new_AGEMA_signal_10822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C ( clk ), .D ( new_AGEMA_signal_10825 ), .Q ( new_AGEMA_signal_10826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C ( clk ), .D ( new_AGEMA_signal_10829 ), .Q ( new_AGEMA_signal_10830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C ( clk ), .D ( new_AGEMA_signal_10833 ), .Q ( new_AGEMA_signal_10834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C ( clk ), .D ( new_AGEMA_signal_10837 ), .Q ( new_AGEMA_signal_10838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C ( clk ), .D ( new_AGEMA_signal_10841 ), .Q ( new_AGEMA_signal_10842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C ( clk ), .D ( new_AGEMA_signal_10845 ), .Q ( new_AGEMA_signal_10846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C ( clk ), .D ( new_AGEMA_signal_10849 ), .Q ( new_AGEMA_signal_10850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C ( clk ), .D ( new_AGEMA_signal_10853 ), .Q ( new_AGEMA_signal_10854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C ( clk ), .D ( new_AGEMA_signal_10857 ), .Q ( new_AGEMA_signal_10858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C ( clk ), .D ( new_AGEMA_signal_10861 ), .Q ( new_AGEMA_signal_10862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C ( clk ), .D ( new_AGEMA_signal_10865 ), .Q ( new_AGEMA_signal_10866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C ( clk ), .D ( new_AGEMA_signal_10867 ), .Q ( new_AGEMA_signal_10868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C ( clk ), .D ( new_AGEMA_signal_10869 ), .Q ( new_AGEMA_signal_10870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C ( clk ), .D ( new_AGEMA_signal_10871 ), .Q ( new_AGEMA_signal_10872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C ( clk ), .D ( new_AGEMA_signal_10873 ), .Q ( new_AGEMA_signal_10874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C ( clk ), .D ( new_AGEMA_signal_10875 ), .Q ( new_AGEMA_signal_10876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C ( clk ), .D ( new_AGEMA_signal_10877 ), .Q ( new_AGEMA_signal_10878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C ( clk ), .D ( new_AGEMA_signal_10879 ), .Q ( new_AGEMA_signal_10880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C ( clk ), .D ( new_AGEMA_signal_10881 ), .Q ( new_AGEMA_signal_10882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C ( clk ), .D ( new_AGEMA_signal_10883 ), .Q ( new_AGEMA_signal_10884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C ( clk ), .D ( new_AGEMA_signal_10885 ), .Q ( new_AGEMA_signal_10886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C ( clk ), .D ( new_AGEMA_signal_10887 ), .Q ( new_AGEMA_signal_10888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C ( clk ), .D ( new_AGEMA_signal_10889 ), .Q ( new_AGEMA_signal_10890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C ( clk ), .D ( new_AGEMA_signal_10891 ), .Q ( new_AGEMA_signal_10892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C ( clk ), .D ( new_AGEMA_signal_10893 ), .Q ( new_AGEMA_signal_10894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C ( clk ), .D ( new_AGEMA_signal_10895 ), .Q ( new_AGEMA_signal_10896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C ( clk ), .D ( new_AGEMA_signal_10897 ), .Q ( new_AGEMA_signal_10898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C ( clk ), .D ( new_AGEMA_signal_10901 ), .Q ( new_AGEMA_signal_10902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C ( clk ), .D ( new_AGEMA_signal_10905 ), .Q ( new_AGEMA_signal_10906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C ( clk ), .D ( new_AGEMA_signal_10909 ), .Q ( new_AGEMA_signal_10910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C ( clk ), .D ( new_AGEMA_signal_10913 ), .Q ( new_AGEMA_signal_10914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C ( clk ), .D ( new_AGEMA_signal_10917 ), .Q ( new_AGEMA_signal_10918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C ( clk ), .D ( new_AGEMA_signal_10921 ), .Q ( new_AGEMA_signal_10922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C ( clk ), .D ( new_AGEMA_signal_10925 ), .Q ( new_AGEMA_signal_10926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C ( clk ), .D ( new_AGEMA_signal_10929 ), .Q ( new_AGEMA_signal_10930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C ( clk ), .D ( new_AGEMA_signal_10931 ), .Q ( new_AGEMA_signal_10932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C ( clk ), .D ( new_AGEMA_signal_10933 ), .Q ( new_AGEMA_signal_10934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C ( clk ), .D ( new_AGEMA_signal_10935 ), .Q ( new_AGEMA_signal_10936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C ( clk ), .D ( new_AGEMA_signal_10937 ), .Q ( new_AGEMA_signal_10938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C ( clk ), .D ( new_AGEMA_signal_10939 ), .Q ( new_AGEMA_signal_10940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C ( clk ), .D ( new_AGEMA_signal_10941 ), .Q ( new_AGEMA_signal_10942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C ( clk ), .D ( new_AGEMA_signal_10943 ), .Q ( new_AGEMA_signal_10944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C ( clk ), .D ( new_AGEMA_signal_10945 ), .Q ( new_AGEMA_signal_10946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2920 ( .C ( clk ), .D ( new_AGEMA_signal_10947 ), .Q ( new_AGEMA_signal_10948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C ( clk ), .D ( new_AGEMA_signal_10949 ), .Q ( new_AGEMA_signal_10950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C ( clk ), .D ( new_AGEMA_signal_10951 ), .Q ( new_AGEMA_signal_10952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2926 ( .C ( clk ), .D ( new_AGEMA_signal_10953 ), .Q ( new_AGEMA_signal_10954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2928 ( .C ( clk ), .D ( new_AGEMA_signal_10955 ), .Q ( new_AGEMA_signal_10956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2930 ( .C ( clk ), .D ( new_AGEMA_signal_10957 ), .Q ( new_AGEMA_signal_10958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2932 ( .C ( clk ), .D ( new_AGEMA_signal_10959 ), .Q ( new_AGEMA_signal_10960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C ( clk ), .D ( new_AGEMA_signal_10961 ), .Q ( new_AGEMA_signal_10962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C ( clk ), .D ( new_AGEMA_signal_10963 ), .Q ( new_AGEMA_signal_10964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2938 ( .C ( clk ), .D ( new_AGEMA_signal_10965 ), .Q ( new_AGEMA_signal_10966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2940 ( .C ( clk ), .D ( new_AGEMA_signal_10967 ), .Q ( new_AGEMA_signal_10968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2942 ( .C ( clk ), .D ( new_AGEMA_signal_10969 ), .Q ( new_AGEMA_signal_10970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2944 ( .C ( clk ), .D ( new_AGEMA_signal_10971 ), .Q ( new_AGEMA_signal_10972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2946 ( .C ( clk ), .D ( new_AGEMA_signal_10973 ), .Q ( new_AGEMA_signal_10974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2948 ( .C ( clk ), .D ( new_AGEMA_signal_10975 ), .Q ( new_AGEMA_signal_10976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2950 ( .C ( clk ), .D ( new_AGEMA_signal_10977 ), .Q ( new_AGEMA_signal_10978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2952 ( .C ( clk ), .D ( new_AGEMA_signal_10979 ), .Q ( new_AGEMA_signal_10980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2954 ( .C ( clk ), .D ( new_AGEMA_signal_10981 ), .Q ( new_AGEMA_signal_10982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2956 ( .C ( clk ), .D ( new_AGEMA_signal_10983 ), .Q ( new_AGEMA_signal_10984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2958 ( .C ( clk ), .D ( new_AGEMA_signal_10985 ), .Q ( new_AGEMA_signal_10986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2960 ( .C ( clk ), .D ( new_AGEMA_signal_10987 ), .Q ( new_AGEMA_signal_10988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2962 ( .C ( clk ), .D ( new_AGEMA_signal_10989 ), .Q ( new_AGEMA_signal_10990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2964 ( .C ( clk ), .D ( new_AGEMA_signal_10991 ), .Q ( new_AGEMA_signal_10992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2966 ( .C ( clk ), .D ( new_AGEMA_signal_10993 ), .Q ( new_AGEMA_signal_10994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2968 ( .C ( clk ), .D ( new_AGEMA_signal_10995 ), .Q ( new_AGEMA_signal_10996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2970 ( .C ( clk ), .D ( new_AGEMA_signal_10997 ), .Q ( new_AGEMA_signal_10998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2972 ( .C ( clk ), .D ( new_AGEMA_signal_10999 ), .Q ( new_AGEMA_signal_11000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2974 ( .C ( clk ), .D ( new_AGEMA_signal_11001 ), .Q ( new_AGEMA_signal_11002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2978 ( .C ( clk ), .D ( new_AGEMA_signal_11005 ), .Q ( new_AGEMA_signal_11006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2982 ( .C ( clk ), .D ( new_AGEMA_signal_11009 ), .Q ( new_AGEMA_signal_11010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2986 ( .C ( clk ), .D ( new_AGEMA_signal_11013 ), .Q ( new_AGEMA_signal_11014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2990 ( .C ( clk ), .D ( new_AGEMA_signal_11017 ), .Q ( new_AGEMA_signal_11018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2992 ( .C ( clk ), .D ( new_AGEMA_signal_11019 ), .Q ( new_AGEMA_signal_11020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2994 ( .C ( clk ), .D ( new_AGEMA_signal_11021 ), .Q ( new_AGEMA_signal_11022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2996 ( .C ( clk ), .D ( new_AGEMA_signal_11023 ), .Q ( new_AGEMA_signal_11024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_2998 ( .C ( clk ), .D ( new_AGEMA_signal_11025 ), .Q ( new_AGEMA_signal_11026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3000 ( .C ( clk ), .D ( new_AGEMA_signal_11027 ), .Q ( new_AGEMA_signal_11028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3002 ( .C ( clk ), .D ( new_AGEMA_signal_11029 ), .Q ( new_AGEMA_signal_11030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3004 ( .C ( clk ), .D ( new_AGEMA_signal_11031 ), .Q ( new_AGEMA_signal_11032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3006 ( .C ( clk ), .D ( new_AGEMA_signal_11033 ), .Q ( new_AGEMA_signal_11034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3008 ( .C ( clk ), .D ( new_AGEMA_signal_11035 ), .Q ( new_AGEMA_signal_11036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3010 ( .C ( clk ), .D ( new_AGEMA_signal_11037 ), .Q ( new_AGEMA_signal_11038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3012 ( .C ( clk ), .D ( new_AGEMA_signal_11039 ), .Q ( new_AGEMA_signal_11040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3014 ( .C ( clk ), .D ( new_AGEMA_signal_11041 ), .Q ( new_AGEMA_signal_11042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3016 ( .C ( clk ), .D ( new_AGEMA_signal_11043 ), .Q ( new_AGEMA_signal_11044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3018 ( .C ( clk ), .D ( new_AGEMA_signal_11045 ), .Q ( new_AGEMA_signal_11046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3020 ( .C ( clk ), .D ( new_AGEMA_signal_11047 ), .Q ( new_AGEMA_signal_11048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3022 ( .C ( clk ), .D ( new_AGEMA_signal_11049 ), .Q ( new_AGEMA_signal_11050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3024 ( .C ( clk ), .D ( new_AGEMA_signal_11051 ), .Q ( new_AGEMA_signal_11052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3026 ( .C ( clk ), .D ( new_AGEMA_signal_11053 ), .Q ( new_AGEMA_signal_11054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3028 ( .C ( clk ), .D ( new_AGEMA_signal_11055 ), .Q ( new_AGEMA_signal_11056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3030 ( .C ( clk ), .D ( new_AGEMA_signal_11057 ), .Q ( new_AGEMA_signal_11058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3034 ( .C ( clk ), .D ( new_AGEMA_signal_11061 ), .Q ( new_AGEMA_signal_11062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3038 ( .C ( clk ), .D ( new_AGEMA_signal_11065 ), .Q ( new_AGEMA_signal_11066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3042 ( .C ( clk ), .D ( new_AGEMA_signal_11069 ), .Q ( new_AGEMA_signal_11070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3046 ( .C ( clk ), .D ( new_AGEMA_signal_11073 ), .Q ( new_AGEMA_signal_11074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3050 ( .C ( clk ), .D ( new_AGEMA_signal_11077 ), .Q ( new_AGEMA_signal_11078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3054 ( .C ( clk ), .D ( new_AGEMA_signal_11081 ), .Q ( new_AGEMA_signal_11082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3058 ( .C ( clk ), .D ( new_AGEMA_signal_11085 ), .Q ( new_AGEMA_signal_11086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3062 ( .C ( clk ), .D ( new_AGEMA_signal_11089 ), .Q ( new_AGEMA_signal_11090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3066 ( .C ( clk ), .D ( new_AGEMA_signal_11093 ), .Q ( new_AGEMA_signal_11094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3070 ( .C ( clk ), .D ( new_AGEMA_signal_11097 ), .Q ( new_AGEMA_signal_11098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3074 ( .C ( clk ), .D ( new_AGEMA_signal_11101 ), .Q ( new_AGEMA_signal_11102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3078 ( .C ( clk ), .D ( new_AGEMA_signal_11105 ), .Q ( new_AGEMA_signal_11106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3082 ( .C ( clk ), .D ( new_AGEMA_signal_11109 ), .Q ( new_AGEMA_signal_11110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3086 ( .C ( clk ), .D ( new_AGEMA_signal_11113 ), .Q ( new_AGEMA_signal_11114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3090 ( .C ( clk ), .D ( new_AGEMA_signal_11117 ), .Q ( new_AGEMA_signal_11118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3094 ( .C ( clk ), .D ( new_AGEMA_signal_11121 ), .Q ( new_AGEMA_signal_11122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3096 ( .C ( clk ), .D ( new_AGEMA_signal_11123 ), .Q ( new_AGEMA_signal_11124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3100 ( .C ( clk ), .D ( new_AGEMA_signal_11127 ), .Q ( new_AGEMA_signal_11128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3104 ( .C ( clk ), .D ( new_AGEMA_signal_11131 ), .Q ( new_AGEMA_signal_11132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3108 ( .C ( clk ), .D ( new_AGEMA_signal_11135 ), .Q ( new_AGEMA_signal_11136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3112 ( .C ( clk ), .D ( new_AGEMA_signal_11139 ), .Q ( new_AGEMA_signal_11140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3116 ( .C ( clk ), .D ( new_AGEMA_signal_11143 ), .Q ( new_AGEMA_signal_11144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3120 ( .C ( clk ), .D ( new_AGEMA_signal_11147 ), .Q ( new_AGEMA_signal_11148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3124 ( .C ( clk ), .D ( new_AGEMA_signal_11151 ), .Q ( new_AGEMA_signal_11152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3132 ( .C ( clk ), .D ( new_AGEMA_signal_11159 ), .Q ( new_AGEMA_signal_11160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3140 ( .C ( clk ), .D ( new_AGEMA_signal_11167 ), .Q ( new_AGEMA_signal_11168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3148 ( .C ( clk ), .D ( new_AGEMA_signal_11175 ), .Q ( new_AGEMA_signal_11176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3156 ( .C ( clk ), .D ( new_AGEMA_signal_11183 ), .Q ( new_AGEMA_signal_11184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3172 ( .C ( clk ), .D ( new_AGEMA_signal_11199 ), .Q ( new_AGEMA_signal_11200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3180 ( .C ( clk ), .D ( new_AGEMA_signal_11207 ), .Q ( new_AGEMA_signal_11208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3188 ( .C ( clk ), .D ( new_AGEMA_signal_11215 ), .Q ( new_AGEMA_signal_11216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3196 ( .C ( clk ), .D ( new_AGEMA_signal_11223 ), .Q ( new_AGEMA_signal_11224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3202 ( .C ( clk ), .D ( new_AGEMA_signal_11229 ), .Q ( new_AGEMA_signal_11230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3208 ( .C ( clk ), .D ( new_AGEMA_signal_11235 ), .Q ( new_AGEMA_signal_11236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3214 ( .C ( clk ), .D ( new_AGEMA_signal_11241 ), .Q ( new_AGEMA_signal_11242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3220 ( .C ( clk ), .D ( new_AGEMA_signal_11247 ), .Q ( new_AGEMA_signal_11248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3224 ( .C ( clk ), .D ( new_AGEMA_signal_11251 ), .Q ( new_AGEMA_signal_11252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3228 ( .C ( clk ), .D ( new_AGEMA_signal_11255 ), .Q ( new_AGEMA_signal_11256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3232 ( .C ( clk ), .D ( new_AGEMA_signal_11259 ), .Q ( new_AGEMA_signal_11260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3236 ( .C ( clk ), .D ( new_AGEMA_signal_11263 ), .Q ( new_AGEMA_signal_11264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3242 ( .C ( clk ), .D ( new_AGEMA_signal_11269 ), .Q ( new_AGEMA_signal_11270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3248 ( .C ( clk ), .D ( new_AGEMA_signal_11275 ), .Q ( new_AGEMA_signal_11276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3254 ( .C ( clk ), .D ( new_AGEMA_signal_11281 ), .Q ( new_AGEMA_signal_11282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3260 ( .C ( clk ), .D ( new_AGEMA_signal_11287 ), .Q ( new_AGEMA_signal_11288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3274 ( .C ( clk ), .D ( new_AGEMA_signal_11301 ), .Q ( new_AGEMA_signal_11302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3280 ( .C ( clk ), .D ( new_AGEMA_signal_11307 ), .Q ( new_AGEMA_signal_11308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3286 ( .C ( clk ), .D ( new_AGEMA_signal_11313 ), .Q ( new_AGEMA_signal_11314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3292 ( .C ( clk ), .D ( new_AGEMA_signal_11319 ), .Q ( new_AGEMA_signal_11320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3298 ( .C ( clk ), .D ( new_AGEMA_signal_11325 ), .Q ( new_AGEMA_signal_11326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3304 ( .C ( clk ), .D ( new_AGEMA_signal_11331 ), .Q ( new_AGEMA_signal_11332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3310 ( .C ( clk ), .D ( new_AGEMA_signal_11337 ), .Q ( new_AGEMA_signal_11338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3316 ( .C ( clk ), .D ( new_AGEMA_signal_11343 ), .Q ( new_AGEMA_signal_11344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3328 ( .C ( clk ), .D ( new_AGEMA_signal_11355 ), .Q ( new_AGEMA_signal_11356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3332 ( .C ( clk ), .D ( new_AGEMA_signal_11359 ), .Q ( new_AGEMA_signal_11360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3336 ( .C ( clk ), .D ( new_AGEMA_signal_11363 ), .Q ( new_AGEMA_signal_11364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3340 ( .C ( clk ), .D ( new_AGEMA_signal_11367 ), .Q ( new_AGEMA_signal_11368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3346 ( .C ( clk ), .D ( new_AGEMA_signal_11373 ), .Q ( new_AGEMA_signal_11374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3352 ( .C ( clk ), .D ( new_AGEMA_signal_11379 ), .Q ( new_AGEMA_signal_11380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3358 ( .C ( clk ), .D ( new_AGEMA_signal_11385 ), .Q ( new_AGEMA_signal_11386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3364 ( .C ( clk ), .D ( new_AGEMA_signal_11391 ), .Q ( new_AGEMA_signal_11392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3370 ( .C ( clk ), .D ( new_AGEMA_signal_11397 ), .Q ( new_AGEMA_signal_11398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3376 ( .C ( clk ), .D ( new_AGEMA_signal_11403 ), .Q ( new_AGEMA_signal_11404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3382 ( .C ( clk ), .D ( new_AGEMA_signal_11409 ), .Q ( new_AGEMA_signal_11410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3388 ( .C ( clk ), .D ( new_AGEMA_signal_11415 ), .Q ( new_AGEMA_signal_11416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3402 ( .C ( clk ), .D ( new_AGEMA_signal_11429 ), .Q ( new_AGEMA_signal_11430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3408 ( .C ( clk ), .D ( new_AGEMA_signal_11435 ), .Q ( new_AGEMA_signal_11436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3414 ( .C ( clk ), .D ( new_AGEMA_signal_11441 ), .Q ( new_AGEMA_signal_11442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3420 ( .C ( clk ), .D ( new_AGEMA_signal_11447 ), .Q ( new_AGEMA_signal_11448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3432 ( .C ( clk ), .D ( new_AGEMA_signal_11459 ), .Q ( new_AGEMA_signal_11460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3436 ( .C ( clk ), .D ( new_AGEMA_signal_11463 ), .Q ( new_AGEMA_signal_11464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3440 ( .C ( clk ), .D ( new_AGEMA_signal_11467 ), .Q ( new_AGEMA_signal_11468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3444 ( .C ( clk ), .D ( new_AGEMA_signal_11471 ), .Q ( new_AGEMA_signal_11472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3448 ( .C ( clk ), .D ( new_AGEMA_signal_11475 ), .Q ( new_AGEMA_signal_11476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3452 ( .C ( clk ), .D ( new_AGEMA_signal_11479 ), .Q ( new_AGEMA_signal_11480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3456 ( .C ( clk ), .D ( new_AGEMA_signal_11483 ), .Q ( new_AGEMA_signal_11484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3460 ( .C ( clk ), .D ( new_AGEMA_signal_11487 ), .Q ( new_AGEMA_signal_11488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3476 ( .C ( clk ), .D ( new_AGEMA_signal_11503 ), .Q ( new_AGEMA_signal_11504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3484 ( .C ( clk ), .D ( new_AGEMA_signal_11511 ), .Q ( new_AGEMA_signal_11512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3492 ( .C ( clk ), .D ( new_AGEMA_signal_11519 ), .Q ( new_AGEMA_signal_11520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3500 ( .C ( clk ), .D ( new_AGEMA_signal_11527 ), .Q ( new_AGEMA_signal_11528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3506 ( .C ( clk ), .D ( new_AGEMA_signal_11533 ), .Q ( new_AGEMA_signal_11534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3512 ( .C ( clk ), .D ( new_AGEMA_signal_11539 ), .Q ( new_AGEMA_signal_11540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3518 ( .C ( clk ), .D ( new_AGEMA_signal_11545 ), .Q ( new_AGEMA_signal_11546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3524 ( .C ( clk ), .D ( new_AGEMA_signal_11551 ), .Q ( new_AGEMA_signal_11552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3528 ( .C ( clk ), .D ( new_AGEMA_signal_11555 ), .Q ( new_AGEMA_signal_11556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3532 ( .C ( clk ), .D ( new_AGEMA_signal_11559 ), .Q ( new_AGEMA_signal_11560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3536 ( .C ( clk ), .D ( new_AGEMA_signal_11563 ), .Q ( new_AGEMA_signal_11564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3540 ( .C ( clk ), .D ( new_AGEMA_signal_11567 ), .Q ( new_AGEMA_signal_11568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3544 ( .C ( clk ), .D ( new_AGEMA_signal_11571 ), .Q ( new_AGEMA_signal_11572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3548 ( .C ( clk ), .D ( new_AGEMA_signal_11575 ), .Q ( new_AGEMA_signal_11576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3552 ( .C ( clk ), .D ( new_AGEMA_signal_11579 ), .Q ( new_AGEMA_signal_11580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3556 ( .C ( clk ), .D ( new_AGEMA_signal_11583 ), .Q ( new_AGEMA_signal_11584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3576 ( .C ( clk ), .D ( new_AGEMA_signal_11603 ), .Q ( new_AGEMA_signal_11604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3580 ( .C ( clk ), .D ( new_AGEMA_signal_11607 ), .Q ( new_AGEMA_signal_11608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3584 ( .C ( clk ), .D ( new_AGEMA_signal_11611 ), .Q ( new_AGEMA_signal_11612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3588 ( .C ( clk ), .D ( new_AGEMA_signal_11615 ), .Q ( new_AGEMA_signal_11616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3592 ( .C ( clk ), .D ( new_AGEMA_signal_11619 ), .Q ( new_AGEMA_signal_11620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3596 ( .C ( clk ), .D ( new_AGEMA_signal_11623 ), .Q ( new_AGEMA_signal_11624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3600 ( .C ( clk ), .D ( new_AGEMA_signal_11627 ), .Q ( new_AGEMA_signal_11628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3604 ( .C ( clk ), .D ( new_AGEMA_signal_11631 ), .Q ( new_AGEMA_signal_11632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3618 ( .C ( clk ), .D ( new_AGEMA_signal_11645 ), .Q ( new_AGEMA_signal_11646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3624 ( .C ( clk ), .D ( new_AGEMA_signal_11651 ), .Q ( new_AGEMA_signal_11652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3630 ( .C ( clk ), .D ( new_AGEMA_signal_11657 ), .Q ( new_AGEMA_signal_11658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3636 ( .C ( clk ), .D ( new_AGEMA_signal_11663 ), .Q ( new_AGEMA_signal_11664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3640 ( .C ( clk ), .D ( new_AGEMA_signal_11667 ), .Q ( new_AGEMA_signal_11668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3644 ( .C ( clk ), .D ( new_AGEMA_signal_11671 ), .Q ( new_AGEMA_signal_11672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3648 ( .C ( clk ), .D ( new_AGEMA_signal_11675 ), .Q ( new_AGEMA_signal_11676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3652 ( .C ( clk ), .D ( new_AGEMA_signal_11679 ), .Q ( new_AGEMA_signal_11680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3664 ( .C ( clk ), .D ( new_AGEMA_signal_11691 ), .Q ( new_AGEMA_signal_11692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3668 ( .C ( clk ), .D ( new_AGEMA_signal_11695 ), .Q ( new_AGEMA_signal_11696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3672 ( .C ( clk ), .D ( new_AGEMA_signal_11699 ), .Q ( new_AGEMA_signal_11700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3676 ( .C ( clk ), .D ( new_AGEMA_signal_11703 ), .Q ( new_AGEMA_signal_11704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3680 ( .C ( clk ), .D ( new_AGEMA_signal_11707 ), .Q ( new_AGEMA_signal_11708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3684 ( .C ( clk ), .D ( new_AGEMA_signal_11711 ), .Q ( new_AGEMA_signal_11712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3688 ( .C ( clk ), .D ( new_AGEMA_signal_11715 ), .Q ( new_AGEMA_signal_11716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3692 ( .C ( clk ), .D ( new_AGEMA_signal_11719 ), .Q ( new_AGEMA_signal_11720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3696 ( .C ( clk ), .D ( new_AGEMA_signal_11723 ), .Q ( new_AGEMA_signal_11724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3700 ( .C ( clk ), .D ( new_AGEMA_signal_11727 ), .Q ( new_AGEMA_signal_11728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3704 ( .C ( clk ), .D ( new_AGEMA_signal_11731 ), .Q ( new_AGEMA_signal_11732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3708 ( .C ( clk ), .D ( new_AGEMA_signal_11735 ), .Q ( new_AGEMA_signal_11736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3720 ( .C ( clk ), .D ( new_AGEMA_signal_11747 ), .Q ( new_AGEMA_signal_11748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3724 ( .C ( clk ), .D ( new_AGEMA_signal_11751 ), .Q ( new_AGEMA_signal_11752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3728 ( .C ( clk ), .D ( new_AGEMA_signal_11755 ), .Q ( new_AGEMA_signal_11756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3732 ( .C ( clk ), .D ( new_AGEMA_signal_11759 ), .Q ( new_AGEMA_signal_11760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3746 ( .C ( clk ), .D ( new_AGEMA_signal_11773 ), .Q ( new_AGEMA_signal_11774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3752 ( .C ( clk ), .D ( new_AGEMA_signal_11779 ), .Q ( new_AGEMA_signal_11780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3758 ( .C ( clk ), .D ( new_AGEMA_signal_11785 ), .Q ( new_AGEMA_signal_11786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3764 ( .C ( clk ), .D ( new_AGEMA_signal_11791 ), .Q ( new_AGEMA_signal_11792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3770 ( .C ( clk ), .D ( new_AGEMA_signal_11797 ), .Q ( new_AGEMA_signal_11798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3776 ( .C ( clk ), .D ( new_AGEMA_signal_11803 ), .Q ( new_AGEMA_signal_11804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3782 ( .C ( clk ), .D ( new_AGEMA_signal_11809 ), .Q ( new_AGEMA_signal_11810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3788 ( .C ( clk ), .D ( new_AGEMA_signal_11815 ), .Q ( new_AGEMA_signal_11816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3792 ( .C ( clk ), .D ( new_AGEMA_signal_11819 ), .Q ( new_AGEMA_signal_11820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3796 ( .C ( clk ), .D ( new_AGEMA_signal_11823 ), .Q ( new_AGEMA_signal_11824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3800 ( .C ( clk ), .D ( new_AGEMA_signal_11827 ), .Q ( new_AGEMA_signal_11828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3804 ( .C ( clk ), .D ( new_AGEMA_signal_11831 ), .Q ( new_AGEMA_signal_11832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3820 ( .C ( clk ), .D ( new_AGEMA_signal_11847 ), .Q ( new_AGEMA_signal_11848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3828 ( .C ( clk ), .D ( new_AGEMA_signal_11855 ), .Q ( new_AGEMA_signal_11856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3836 ( .C ( clk ), .D ( new_AGEMA_signal_11863 ), .Q ( new_AGEMA_signal_11864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3844 ( .C ( clk ), .D ( new_AGEMA_signal_11871 ), .Q ( new_AGEMA_signal_11872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3856 ( .C ( clk ), .D ( new_AGEMA_signal_11883 ), .Q ( new_AGEMA_signal_11884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3860 ( .C ( clk ), .D ( new_AGEMA_signal_11887 ), .Q ( new_AGEMA_signal_11888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3864 ( .C ( clk ), .D ( new_AGEMA_signal_11891 ), .Q ( new_AGEMA_signal_11892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3868 ( .C ( clk ), .D ( new_AGEMA_signal_11895 ), .Q ( new_AGEMA_signal_11896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3872 ( .C ( clk ), .D ( new_AGEMA_signal_11899 ), .Q ( new_AGEMA_signal_11900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3876 ( .C ( clk ), .D ( new_AGEMA_signal_11903 ), .Q ( new_AGEMA_signal_11904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3880 ( .C ( clk ), .D ( new_AGEMA_signal_11907 ), .Q ( new_AGEMA_signal_11908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3884 ( .C ( clk ), .D ( new_AGEMA_signal_11911 ), .Q ( new_AGEMA_signal_11912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3888 ( .C ( clk ), .D ( new_AGEMA_signal_11915 ), .Q ( new_AGEMA_signal_11916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3892 ( .C ( clk ), .D ( new_AGEMA_signal_11919 ), .Q ( new_AGEMA_signal_11920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3896 ( .C ( clk ), .D ( new_AGEMA_signal_11923 ), .Q ( new_AGEMA_signal_11924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3900 ( .C ( clk ), .D ( new_AGEMA_signal_11927 ), .Q ( new_AGEMA_signal_11928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3904 ( .C ( clk ), .D ( new_AGEMA_signal_11931 ), .Q ( new_AGEMA_signal_11932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3908 ( .C ( clk ), .D ( new_AGEMA_signal_11935 ), .Q ( new_AGEMA_signal_11936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3912 ( .C ( clk ), .D ( new_AGEMA_signal_11939 ), .Q ( new_AGEMA_signal_11940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3916 ( .C ( clk ), .D ( new_AGEMA_signal_11943 ), .Q ( new_AGEMA_signal_11944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3920 ( .C ( clk ), .D ( new_AGEMA_signal_11947 ), .Q ( new_AGEMA_signal_11948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3924 ( .C ( clk ), .D ( new_AGEMA_signal_11951 ), .Q ( new_AGEMA_signal_11952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3928 ( .C ( clk ), .D ( new_AGEMA_signal_11955 ), .Q ( new_AGEMA_signal_11956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3932 ( .C ( clk ), .D ( new_AGEMA_signal_11959 ), .Q ( new_AGEMA_signal_11960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3940 ( .C ( clk ), .D ( new_AGEMA_signal_11967 ), .Q ( new_AGEMA_signal_11968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3948 ( .C ( clk ), .D ( new_AGEMA_signal_11975 ), .Q ( new_AGEMA_signal_11976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3956 ( .C ( clk ), .D ( new_AGEMA_signal_11983 ), .Q ( new_AGEMA_signal_11984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3964 ( .C ( clk ), .D ( new_AGEMA_signal_11991 ), .Q ( new_AGEMA_signal_11992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3976 ( .C ( clk ), .D ( new_AGEMA_signal_12003 ), .Q ( new_AGEMA_signal_12004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3980 ( .C ( clk ), .D ( new_AGEMA_signal_12007 ), .Q ( new_AGEMA_signal_12008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3984 ( .C ( clk ), .D ( new_AGEMA_signal_12011 ), .Q ( new_AGEMA_signal_12012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3988 ( .C ( clk ), .D ( new_AGEMA_signal_12015 ), .Q ( new_AGEMA_signal_12016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4002 ( .C ( clk ), .D ( new_AGEMA_signal_12029 ), .Q ( new_AGEMA_signal_12030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4008 ( .C ( clk ), .D ( new_AGEMA_signal_12035 ), .Q ( new_AGEMA_signal_12036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4014 ( .C ( clk ), .D ( new_AGEMA_signal_12041 ), .Q ( new_AGEMA_signal_12042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4020 ( .C ( clk ), .D ( new_AGEMA_signal_12047 ), .Q ( new_AGEMA_signal_12048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4034 ( .C ( clk ), .D ( new_AGEMA_signal_12061 ), .Q ( new_AGEMA_signal_12062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4042 ( .C ( clk ), .D ( new_AGEMA_signal_12069 ), .Q ( new_AGEMA_signal_12070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4050 ( .C ( clk ), .D ( new_AGEMA_signal_12077 ), .Q ( new_AGEMA_signal_12078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4058 ( .C ( clk ), .D ( new_AGEMA_signal_12085 ), .Q ( new_AGEMA_signal_12086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4090 ( .C ( clk ), .D ( new_AGEMA_signal_12117 ), .Q ( new_AGEMA_signal_12118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4098 ( .C ( clk ), .D ( new_AGEMA_signal_12125 ), .Q ( new_AGEMA_signal_12126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4106 ( .C ( clk ), .D ( new_AGEMA_signal_12133 ), .Q ( new_AGEMA_signal_12134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4114 ( .C ( clk ), .D ( new_AGEMA_signal_12141 ), .Q ( new_AGEMA_signal_12142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4128 ( .C ( clk ), .D ( new_AGEMA_signal_12155 ), .Q ( new_AGEMA_signal_12156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4134 ( .C ( clk ), .D ( new_AGEMA_signal_12161 ), .Q ( new_AGEMA_signal_12162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4140 ( .C ( clk ), .D ( new_AGEMA_signal_12167 ), .Q ( new_AGEMA_signal_12168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4146 ( .C ( clk ), .D ( new_AGEMA_signal_12173 ), .Q ( new_AGEMA_signal_12174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4170 ( .C ( clk ), .D ( new_AGEMA_signal_12197 ), .Q ( new_AGEMA_signal_12198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4178 ( .C ( clk ), .D ( new_AGEMA_signal_12205 ), .Q ( new_AGEMA_signal_12206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4186 ( .C ( clk ), .D ( new_AGEMA_signal_12213 ), .Q ( new_AGEMA_signal_12214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4194 ( .C ( clk ), .D ( new_AGEMA_signal_12221 ), .Q ( new_AGEMA_signal_12222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4216 ( .C ( clk ), .D ( new_AGEMA_signal_12243 ), .Q ( new_AGEMA_signal_12244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4222 ( .C ( clk ), .D ( new_AGEMA_signal_12249 ), .Q ( new_AGEMA_signal_12250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4228 ( .C ( clk ), .D ( new_AGEMA_signal_12255 ), .Q ( new_AGEMA_signal_12256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4234 ( .C ( clk ), .D ( new_AGEMA_signal_12261 ), .Q ( new_AGEMA_signal_12262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4240 ( .C ( clk ), .D ( new_AGEMA_signal_12267 ), .Q ( new_AGEMA_signal_12268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4246 ( .C ( clk ), .D ( new_AGEMA_signal_12273 ), .Q ( new_AGEMA_signal_12274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4252 ( .C ( clk ), .D ( new_AGEMA_signal_12279 ), .Q ( new_AGEMA_signal_12280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4258 ( .C ( clk ), .D ( new_AGEMA_signal_12285 ), .Q ( new_AGEMA_signal_12286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4264 ( .C ( clk ), .D ( new_AGEMA_signal_12291 ), .Q ( new_AGEMA_signal_12292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4270 ( .C ( clk ), .D ( new_AGEMA_signal_12297 ), .Q ( new_AGEMA_signal_12298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4276 ( .C ( clk ), .D ( new_AGEMA_signal_12303 ), .Q ( new_AGEMA_signal_12304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4282 ( .C ( clk ), .D ( new_AGEMA_signal_12309 ), .Q ( new_AGEMA_signal_12310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4288 ( .C ( clk ), .D ( new_AGEMA_signal_12315 ), .Q ( new_AGEMA_signal_12316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4294 ( .C ( clk ), .D ( new_AGEMA_signal_12321 ), .Q ( new_AGEMA_signal_12322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4300 ( .C ( clk ), .D ( new_AGEMA_signal_12327 ), .Q ( new_AGEMA_signal_12328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4306 ( .C ( clk ), .D ( new_AGEMA_signal_12333 ), .Q ( new_AGEMA_signal_12334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4312 ( .C ( clk ), .D ( new_AGEMA_signal_12339 ), .Q ( new_AGEMA_signal_12340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4318 ( .C ( clk ), .D ( new_AGEMA_signal_12345 ), .Q ( new_AGEMA_signal_12346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4324 ( .C ( clk ), .D ( new_AGEMA_signal_12351 ), .Q ( new_AGEMA_signal_12352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4330 ( .C ( clk ), .D ( new_AGEMA_signal_12357 ), .Q ( new_AGEMA_signal_12358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4354 ( .C ( clk ), .D ( new_AGEMA_signal_12381 ), .Q ( new_AGEMA_signal_12382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4362 ( .C ( clk ), .D ( new_AGEMA_signal_12389 ), .Q ( new_AGEMA_signal_12390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4370 ( .C ( clk ), .D ( new_AGEMA_signal_12397 ), .Q ( new_AGEMA_signal_12398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4378 ( .C ( clk ), .D ( new_AGEMA_signal_12405 ), .Q ( new_AGEMA_signal_12406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4400 ( .C ( clk ), .D ( new_AGEMA_signal_12427 ), .Q ( new_AGEMA_signal_12428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4406 ( .C ( clk ), .D ( new_AGEMA_signal_12433 ), .Q ( new_AGEMA_signal_12434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4412 ( .C ( clk ), .D ( new_AGEMA_signal_12439 ), .Q ( new_AGEMA_signal_12440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4418 ( .C ( clk ), .D ( new_AGEMA_signal_12445 ), .Q ( new_AGEMA_signal_12446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4426 ( .C ( clk ), .D ( new_AGEMA_signal_12453 ), .Q ( new_AGEMA_signal_12454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4434 ( .C ( clk ), .D ( new_AGEMA_signal_12461 ), .Q ( new_AGEMA_signal_12462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4442 ( .C ( clk ), .D ( new_AGEMA_signal_12469 ), .Q ( new_AGEMA_signal_12470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4450 ( .C ( clk ), .D ( new_AGEMA_signal_12477 ), .Q ( new_AGEMA_signal_12478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4464 ( .C ( clk ), .D ( new_AGEMA_signal_12491 ), .Q ( new_AGEMA_signal_12492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4470 ( .C ( clk ), .D ( new_AGEMA_signal_12497 ), .Q ( new_AGEMA_signal_12498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4476 ( .C ( clk ), .D ( new_AGEMA_signal_12503 ), .Q ( new_AGEMA_signal_12504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4482 ( .C ( clk ), .D ( new_AGEMA_signal_12509 ), .Q ( new_AGEMA_signal_12510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4504 ( .C ( clk ), .D ( new_AGEMA_signal_12531 ), .Q ( new_AGEMA_signal_12532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4510 ( .C ( clk ), .D ( new_AGEMA_signal_12537 ), .Q ( new_AGEMA_signal_12538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4516 ( .C ( clk ), .D ( new_AGEMA_signal_12543 ), .Q ( new_AGEMA_signal_12544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4522 ( .C ( clk ), .D ( new_AGEMA_signal_12549 ), .Q ( new_AGEMA_signal_12550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4528 ( .C ( clk ), .D ( new_AGEMA_signal_12555 ), .Q ( new_AGEMA_signal_12556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4534 ( .C ( clk ), .D ( new_AGEMA_signal_12561 ), .Q ( new_AGEMA_signal_12562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4540 ( .C ( clk ), .D ( new_AGEMA_signal_12567 ), .Q ( new_AGEMA_signal_12568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4546 ( .C ( clk ), .D ( new_AGEMA_signal_12573 ), .Q ( new_AGEMA_signal_12574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4554 ( .C ( clk ), .D ( new_AGEMA_signal_12581 ), .Q ( new_AGEMA_signal_12582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4562 ( .C ( clk ), .D ( new_AGEMA_signal_12589 ), .Q ( new_AGEMA_signal_12590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4570 ( .C ( clk ), .D ( new_AGEMA_signal_12597 ), .Q ( new_AGEMA_signal_12598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4578 ( .C ( clk ), .D ( new_AGEMA_signal_12605 ), .Q ( new_AGEMA_signal_12606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4586 ( .C ( clk ), .D ( new_AGEMA_signal_12613 ), .Q ( new_AGEMA_signal_12614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4594 ( .C ( clk ), .D ( new_AGEMA_signal_12621 ), .Q ( new_AGEMA_signal_12622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4602 ( .C ( clk ), .D ( new_AGEMA_signal_12629 ), .Q ( new_AGEMA_signal_12630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4610 ( .C ( clk ), .D ( new_AGEMA_signal_12637 ), .Q ( new_AGEMA_signal_12638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4616 ( .C ( clk ), .D ( new_AGEMA_signal_12643 ), .Q ( new_AGEMA_signal_12644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4622 ( .C ( clk ), .D ( new_AGEMA_signal_12649 ), .Q ( new_AGEMA_signal_12650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4628 ( .C ( clk ), .D ( new_AGEMA_signal_12655 ), .Q ( new_AGEMA_signal_12656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4634 ( .C ( clk ), .D ( new_AGEMA_signal_12661 ), .Q ( new_AGEMA_signal_12662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4640 ( .C ( clk ), .D ( new_AGEMA_signal_12667 ), .Q ( new_AGEMA_signal_12668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4646 ( .C ( clk ), .D ( new_AGEMA_signal_12673 ), .Q ( new_AGEMA_signal_12674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4652 ( .C ( clk ), .D ( new_AGEMA_signal_12679 ), .Q ( new_AGEMA_signal_12680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4658 ( .C ( clk ), .D ( new_AGEMA_signal_12685 ), .Q ( new_AGEMA_signal_12686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4776 ( .C ( clk ), .D ( new_AGEMA_signal_12803 ), .Q ( new_AGEMA_signal_12804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4784 ( .C ( clk ), .D ( new_AGEMA_signal_12811 ), .Q ( new_AGEMA_signal_12812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4792 ( .C ( clk ), .D ( new_AGEMA_signal_12819 ), .Q ( new_AGEMA_signal_12820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4800 ( .C ( clk ), .D ( new_AGEMA_signal_12827 ), .Q ( new_AGEMA_signal_12828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4808 ( .C ( clk ), .D ( new_AGEMA_signal_12835 ), .Q ( new_AGEMA_signal_12836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4816 ( .C ( clk ), .D ( new_AGEMA_signal_12843 ), .Q ( new_AGEMA_signal_12844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4824 ( .C ( clk ), .D ( new_AGEMA_signal_12851 ), .Q ( new_AGEMA_signal_12852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4832 ( .C ( clk ), .D ( new_AGEMA_signal_12859 ), .Q ( new_AGEMA_signal_12860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4840 ( .C ( clk ), .D ( new_AGEMA_signal_12867 ), .Q ( new_AGEMA_signal_12868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4848 ( .C ( clk ), .D ( new_AGEMA_signal_12875 ), .Q ( new_AGEMA_signal_12876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4856 ( .C ( clk ), .D ( new_AGEMA_signal_12883 ), .Q ( new_AGEMA_signal_12884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4864 ( .C ( clk ), .D ( new_AGEMA_signal_12891 ), .Q ( new_AGEMA_signal_12892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4872 ( .C ( clk ), .D ( new_AGEMA_signal_12899 ), .Q ( new_AGEMA_signal_12900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4880 ( .C ( clk ), .D ( new_AGEMA_signal_12907 ), .Q ( new_AGEMA_signal_12908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4888 ( .C ( clk ), .D ( new_AGEMA_signal_12915 ), .Q ( new_AGEMA_signal_12916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4896 ( .C ( clk ), .D ( new_AGEMA_signal_12923 ), .Q ( new_AGEMA_signal_12924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4930 ( .C ( clk ), .D ( new_AGEMA_signal_12957 ), .Q ( new_AGEMA_signal_12958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4940 ( .C ( clk ), .D ( new_AGEMA_signal_12967 ), .Q ( new_AGEMA_signal_12968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4950 ( .C ( clk ), .D ( new_AGEMA_signal_12977 ), .Q ( new_AGEMA_signal_12978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4960 ( .C ( clk ), .D ( new_AGEMA_signal_12987 ), .Q ( new_AGEMA_signal_12988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4968 ( .C ( clk ), .D ( new_AGEMA_signal_12995 ), .Q ( new_AGEMA_signal_12996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4976 ( .C ( clk ), .D ( new_AGEMA_signal_13003 ), .Q ( new_AGEMA_signal_13004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4984 ( .C ( clk ), .D ( new_AGEMA_signal_13011 ), .Q ( new_AGEMA_signal_13012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4992 ( .C ( clk ), .D ( new_AGEMA_signal_13019 ), .Q ( new_AGEMA_signal_13020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5000 ( .C ( clk ), .D ( new_AGEMA_signal_13027 ), .Q ( new_AGEMA_signal_13028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5008 ( .C ( clk ), .D ( new_AGEMA_signal_13035 ), .Q ( new_AGEMA_signal_13036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5016 ( .C ( clk ), .D ( new_AGEMA_signal_13043 ), .Q ( new_AGEMA_signal_13044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5024 ( .C ( clk ), .D ( new_AGEMA_signal_13051 ), .Q ( new_AGEMA_signal_13052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5032 ( .C ( clk ), .D ( new_AGEMA_signal_13059 ), .Q ( new_AGEMA_signal_13060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5040 ( .C ( clk ), .D ( new_AGEMA_signal_13067 ), .Q ( new_AGEMA_signal_13068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5048 ( .C ( clk ), .D ( new_AGEMA_signal_13075 ), .Q ( new_AGEMA_signal_13076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5056 ( .C ( clk ), .D ( new_AGEMA_signal_13083 ), .Q ( new_AGEMA_signal_13084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5130 ( .C ( clk ), .D ( new_AGEMA_signal_13157 ), .Q ( new_AGEMA_signal_13158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5140 ( .C ( clk ), .D ( new_AGEMA_signal_13167 ), .Q ( new_AGEMA_signal_13168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5150 ( .C ( clk ), .D ( new_AGEMA_signal_13177 ), .Q ( new_AGEMA_signal_13178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5160 ( .C ( clk ), .D ( new_AGEMA_signal_13187 ), .Q ( new_AGEMA_signal_13188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5168 ( .C ( clk ), .D ( new_AGEMA_signal_13195 ), .Q ( new_AGEMA_signal_13196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5176 ( .C ( clk ), .D ( new_AGEMA_signal_13203 ), .Q ( new_AGEMA_signal_13204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5184 ( .C ( clk ), .D ( new_AGEMA_signal_13211 ), .Q ( new_AGEMA_signal_13212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5192 ( .C ( clk ), .D ( new_AGEMA_signal_13219 ), .Q ( new_AGEMA_signal_13220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C ( clk ), .D ( new_AGEMA_signal_13251 ), .Q ( new_AGEMA_signal_13252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C ( clk ), .D ( new_AGEMA_signal_13259 ), .Q ( new_AGEMA_signal_13260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C ( clk ), .D ( new_AGEMA_signal_13267 ), .Q ( new_AGEMA_signal_13268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C ( clk ), .D ( new_AGEMA_signal_13275 ), .Q ( new_AGEMA_signal_13276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5256 ( .C ( clk ), .D ( new_AGEMA_signal_13283 ), .Q ( new_AGEMA_signal_13284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5264 ( .C ( clk ), .D ( new_AGEMA_signal_13291 ), .Q ( new_AGEMA_signal_13292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5272 ( .C ( clk ), .D ( new_AGEMA_signal_13299 ), .Q ( new_AGEMA_signal_13300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5280 ( .C ( clk ), .D ( new_AGEMA_signal_13307 ), .Q ( new_AGEMA_signal_13308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5328 ( .C ( clk ), .D ( new_AGEMA_signal_13355 ), .Q ( new_AGEMA_signal_13356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5336 ( .C ( clk ), .D ( new_AGEMA_signal_13363 ), .Q ( new_AGEMA_signal_13364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5344 ( .C ( clk ), .D ( new_AGEMA_signal_13371 ), .Q ( new_AGEMA_signal_13372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5352 ( .C ( clk ), .D ( new_AGEMA_signal_13379 ), .Q ( new_AGEMA_signal_13380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5592 ( .C ( clk ), .D ( new_AGEMA_signal_13619 ), .Q ( new_AGEMA_signal_13620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5602 ( .C ( clk ), .D ( new_AGEMA_signal_13629 ), .Q ( new_AGEMA_signal_13630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5612 ( .C ( clk ), .D ( new_AGEMA_signal_13639 ), .Q ( new_AGEMA_signal_13640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5622 ( .C ( clk ), .D ( new_AGEMA_signal_13649 ), .Q ( new_AGEMA_signal_13650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6376 ( .C ( clk ), .D ( new_AGEMA_signal_14403 ), .Q ( new_AGEMA_signal_14404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6390 ( .C ( clk ), .D ( new_AGEMA_signal_14417 ), .Q ( new_AGEMA_signal_14418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6404 ( .C ( clk ), .D ( new_AGEMA_signal_14431 ), .Q ( new_AGEMA_signal_14432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6418 ( .C ( clk ), .D ( new_AGEMA_signal_14445 ), .Q ( new_AGEMA_signal_14446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6464 ( .C ( clk ), .D ( new_AGEMA_signal_14491 ), .Q ( new_AGEMA_signal_14492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6478 ( .C ( clk ), .D ( new_AGEMA_signal_14505 ), .Q ( new_AGEMA_signal_14506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6492 ( .C ( clk ), .D ( new_AGEMA_signal_14519 ), .Q ( new_AGEMA_signal_14520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6506 ( .C ( clk ), .D ( new_AGEMA_signal_14533 ), .Q ( new_AGEMA_signal_14534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6608 ( .C ( clk ), .D ( new_AGEMA_signal_14635 ), .Q ( new_AGEMA_signal_14636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6624 ( .C ( clk ), .D ( new_AGEMA_signal_14651 ), .Q ( new_AGEMA_signal_14652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6640 ( .C ( clk ), .D ( new_AGEMA_signal_14667 ), .Q ( new_AGEMA_signal_14668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6656 ( .C ( clk ), .D ( new_AGEMA_signal_14683 ), .Q ( new_AGEMA_signal_14684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6696 ( .C ( clk ), .D ( new_AGEMA_signal_14723 ), .Q ( new_AGEMA_signal_14724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6712 ( .C ( clk ), .D ( new_AGEMA_signal_14739 ), .Q ( new_AGEMA_signal_14740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6728 ( .C ( clk ), .D ( new_AGEMA_signal_14755 ), .Q ( new_AGEMA_signal_14756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6744 ( .C ( clk ), .D ( new_AGEMA_signal_14771 ), .Q ( new_AGEMA_signal_14772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7000 ( .C ( clk ), .D ( new_AGEMA_signal_15027 ), .Q ( new_AGEMA_signal_15028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7018 ( .C ( clk ), .D ( new_AGEMA_signal_15045 ), .Q ( new_AGEMA_signal_15046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7036 ( .C ( clk ), .D ( new_AGEMA_signal_15063 ), .Q ( new_AGEMA_signal_15064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7054 ( .C ( clk ), .D ( new_AGEMA_signal_15081 ), .Q ( new_AGEMA_signal_15082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7200 ( .C ( clk ), .D ( new_AGEMA_signal_15227 ), .Q ( new_AGEMA_signal_15228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7220 ( .C ( clk ), .D ( new_AGEMA_signal_15247 ), .Q ( new_AGEMA_signal_15248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7240 ( .C ( clk ), .D ( new_AGEMA_signal_15267 ), .Q ( new_AGEMA_signal_15268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7260 ( .C ( clk ), .D ( new_AGEMA_signal_15287 ), .Q ( new_AGEMA_signal_15288 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_3097 ( .C ( clk ), .D ( new_AGEMA_signal_11124 ), .Q ( new_AGEMA_signal_11125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3101 ( .C ( clk ), .D ( new_AGEMA_signal_11128 ), .Q ( new_AGEMA_signal_11129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3105 ( .C ( clk ), .D ( new_AGEMA_signal_11132 ), .Q ( new_AGEMA_signal_11133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3109 ( .C ( clk ), .D ( new_AGEMA_signal_11136 ), .Q ( new_AGEMA_signal_11137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3113 ( .C ( clk ), .D ( new_AGEMA_signal_11140 ), .Q ( new_AGEMA_signal_11141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3117 ( .C ( clk ), .D ( new_AGEMA_signal_11144 ), .Q ( new_AGEMA_signal_11145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3121 ( .C ( clk ), .D ( new_AGEMA_signal_11148 ), .Q ( new_AGEMA_signal_11149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3125 ( .C ( clk ), .D ( new_AGEMA_signal_11152 ), .Q ( new_AGEMA_signal_11153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3133 ( .C ( clk ), .D ( new_AGEMA_signal_11160 ), .Q ( new_AGEMA_signal_11161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3141 ( .C ( clk ), .D ( new_AGEMA_signal_11168 ), .Q ( new_AGEMA_signal_11169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3149 ( .C ( clk ), .D ( new_AGEMA_signal_11176 ), .Q ( new_AGEMA_signal_11177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3157 ( .C ( clk ), .D ( new_AGEMA_signal_11184 ), .Q ( new_AGEMA_signal_11185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3159 ( .C ( clk ), .D ( n1978 ), .Q ( new_AGEMA_signal_11187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3161 ( .C ( clk ), .D ( new_AGEMA_signal_2562 ), .Q ( new_AGEMA_signal_11189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3163 ( .C ( clk ), .D ( new_AGEMA_signal_2563 ), .Q ( new_AGEMA_signal_11191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3165 ( .C ( clk ), .D ( new_AGEMA_signal_2564 ), .Q ( new_AGEMA_signal_11193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3173 ( .C ( clk ), .D ( new_AGEMA_signal_11200 ), .Q ( new_AGEMA_signal_11201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3181 ( .C ( clk ), .D ( new_AGEMA_signal_11208 ), .Q ( new_AGEMA_signal_11209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3189 ( .C ( clk ), .D ( new_AGEMA_signal_11216 ), .Q ( new_AGEMA_signal_11217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3197 ( .C ( clk ), .D ( new_AGEMA_signal_11224 ), .Q ( new_AGEMA_signal_11225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3203 ( .C ( clk ), .D ( new_AGEMA_signal_11230 ), .Q ( new_AGEMA_signal_11231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3209 ( .C ( clk ), .D ( new_AGEMA_signal_11236 ), .Q ( new_AGEMA_signal_11237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3215 ( .C ( clk ), .D ( new_AGEMA_signal_11242 ), .Q ( new_AGEMA_signal_11243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3221 ( .C ( clk ), .D ( new_AGEMA_signal_11248 ), .Q ( new_AGEMA_signal_11249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3225 ( .C ( clk ), .D ( new_AGEMA_signal_11252 ), .Q ( new_AGEMA_signal_11253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3229 ( .C ( clk ), .D ( new_AGEMA_signal_11256 ), .Q ( new_AGEMA_signal_11257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3233 ( .C ( clk ), .D ( new_AGEMA_signal_11260 ), .Q ( new_AGEMA_signal_11261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3237 ( .C ( clk ), .D ( new_AGEMA_signal_11264 ), .Q ( new_AGEMA_signal_11265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3243 ( .C ( clk ), .D ( new_AGEMA_signal_11270 ), .Q ( new_AGEMA_signal_11271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3249 ( .C ( clk ), .D ( new_AGEMA_signal_11276 ), .Q ( new_AGEMA_signal_11277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3255 ( .C ( clk ), .D ( new_AGEMA_signal_11282 ), .Q ( new_AGEMA_signal_11283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3261 ( .C ( clk ), .D ( new_AGEMA_signal_11288 ), .Q ( new_AGEMA_signal_11289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3263 ( .C ( clk ), .D ( new_AGEMA_signal_10902 ), .Q ( new_AGEMA_signal_11291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3265 ( .C ( clk ), .D ( new_AGEMA_signal_10906 ), .Q ( new_AGEMA_signal_11293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3267 ( .C ( clk ), .D ( new_AGEMA_signal_10910 ), .Q ( new_AGEMA_signal_11295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3269 ( .C ( clk ), .D ( new_AGEMA_signal_10914 ), .Q ( new_AGEMA_signal_11297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3275 ( .C ( clk ), .D ( new_AGEMA_signal_11302 ), .Q ( new_AGEMA_signal_11303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3281 ( .C ( clk ), .D ( new_AGEMA_signal_11308 ), .Q ( new_AGEMA_signal_11309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3287 ( .C ( clk ), .D ( new_AGEMA_signal_11314 ), .Q ( new_AGEMA_signal_11315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3293 ( .C ( clk ), .D ( new_AGEMA_signal_11320 ), .Q ( new_AGEMA_signal_11321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3299 ( .C ( clk ), .D ( new_AGEMA_signal_11326 ), .Q ( new_AGEMA_signal_11327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3305 ( .C ( clk ), .D ( new_AGEMA_signal_11332 ), .Q ( new_AGEMA_signal_11333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3311 ( .C ( clk ), .D ( new_AGEMA_signal_11338 ), .Q ( new_AGEMA_signal_11339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3317 ( .C ( clk ), .D ( new_AGEMA_signal_11344 ), .Q ( new_AGEMA_signal_11345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3319 ( .C ( clk ), .D ( n2091 ), .Q ( new_AGEMA_signal_11347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3321 ( .C ( clk ), .D ( new_AGEMA_signal_2616 ), .Q ( new_AGEMA_signal_11349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3323 ( .C ( clk ), .D ( new_AGEMA_signal_2617 ), .Q ( new_AGEMA_signal_11351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3325 ( .C ( clk ), .D ( new_AGEMA_signal_2618 ), .Q ( new_AGEMA_signal_11353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3329 ( .C ( clk ), .D ( new_AGEMA_signal_11356 ), .Q ( new_AGEMA_signal_11357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3333 ( .C ( clk ), .D ( new_AGEMA_signal_11360 ), .Q ( new_AGEMA_signal_11361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3337 ( .C ( clk ), .D ( new_AGEMA_signal_11364 ), .Q ( new_AGEMA_signal_11365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3341 ( .C ( clk ), .D ( new_AGEMA_signal_11368 ), .Q ( new_AGEMA_signal_11369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3347 ( .C ( clk ), .D ( new_AGEMA_signal_11374 ), .Q ( new_AGEMA_signal_11375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3353 ( .C ( clk ), .D ( new_AGEMA_signal_11380 ), .Q ( new_AGEMA_signal_11381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3359 ( .C ( clk ), .D ( new_AGEMA_signal_11386 ), .Q ( new_AGEMA_signal_11387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3365 ( .C ( clk ), .D ( new_AGEMA_signal_11392 ), .Q ( new_AGEMA_signal_11393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3371 ( .C ( clk ), .D ( new_AGEMA_signal_11398 ), .Q ( new_AGEMA_signal_11399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3377 ( .C ( clk ), .D ( new_AGEMA_signal_11404 ), .Q ( new_AGEMA_signal_11405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3383 ( .C ( clk ), .D ( new_AGEMA_signal_11410 ), .Q ( new_AGEMA_signal_11411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3389 ( .C ( clk ), .D ( new_AGEMA_signal_11416 ), .Q ( new_AGEMA_signal_11417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3391 ( .C ( clk ), .D ( n2543 ), .Q ( new_AGEMA_signal_11419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3393 ( .C ( clk ), .D ( new_AGEMA_signal_2634 ), .Q ( new_AGEMA_signal_11421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3395 ( .C ( clk ), .D ( new_AGEMA_signal_2635 ), .Q ( new_AGEMA_signal_11423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3397 ( .C ( clk ), .D ( new_AGEMA_signal_2636 ), .Q ( new_AGEMA_signal_11425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3403 ( .C ( clk ), .D ( new_AGEMA_signal_11430 ), .Q ( new_AGEMA_signal_11431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3409 ( .C ( clk ), .D ( new_AGEMA_signal_11436 ), .Q ( new_AGEMA_signal_11437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3415 ( .C ( clk ), .D ( new_AGEMA_signal_11442 ), .Q ( new_AGEMA_signal_11443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3421 ( .C ( clk ), .D ( new_AGEMA_signal_11448 ), .Q ( new_AGEMA_signal_11449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3423 ( .C ( clk ), .D ( n2159 ), .Q ( new_AGEMA_signal_11451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3425 ( .C ( clk ), .D ( new_AGEMA_signal_2646 ), .Q ( new_AGEMA_signal_11453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3427 ( .C ( clk ), .D ( new_AGEMA_signal_2647 ), .Q ( new_AGEMA_signal_11455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3429 ( .C ( clk ), .D ( new_AGEMA_signal_2648 ), .Q ( new_AGEMA_signal_11457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3433 ( .C ( clk ), .D ( new_AGEMA_signal_11460 ), .Q ( new_AGEMA_signal_11461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3437 ( .C ( clk ), .D ( new_AGEMA_signal_11464 ), .Q ( new_AGEMA_signal_11465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3441 ( .C ( clk ), .D ( new_AGEMA_signal_11468 ), .Q ( new_AGEMA_signal_11469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3445 ( .C ( clk ), .D ( new_AGEMA_signal_11472 ), .Q ( new_AGEMA_signal_11473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3449 ( .C ( clk ), .D ( new_AGEMA_signal_11476 ), .Q ( new_AGEMA_signal_11477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3453 ( .C ( clk ), .D ( new_AGEMA_signal_11480 ), .Q ( new_AGEMA_signal_11481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3457 ( .C ( clk ), .D ( new_AGEMA_signal_11484 ), .Q ( new_AGEMA_signal_11485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3461 ( .C ( clk ), .D ( new_AGEMA_signal_11488 ), .Q ( new_AGEMA_signal_11489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3463 ( .C ( clk ), .D ( new_AGEMA_signal_10876 ), .Q ( new_AGEMA_signal_11491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3465 ( .C ( clk ), .D ( new_AGEMA_signal_10878 ), .Q ( new_AGEMA_signal_11493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3467 ( .C ( clk ), .D ( new_AGEMA_signal_10880 ), .Q ( new_AGEMA_signal_11495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3469 ( .C ( clk ), .D ( new_AGEMA_signal_10882 ), .Q ( new_AGEMA_signal_11497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3477 ( .C ( clk ), .D ( new_AGEMA_signal_11504 ), .Q ( new_AGEMA_signal_11505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3485 ( .C ( clk ), .D ( new_AGEMA_signal_11512 ), .Q ( new_AGEMA_signal_11513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3493 ( .C ( clk ), .D ( new_AGEMA_signal_11520 ), .Q ( new_AGEMA_signal_11521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3501 ( .C ( clk ), .D ( new_AGEMA_signal_11528 ), .Q ( new_AGEMA_signal_11529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3507 ( .C ( clk ), .D ( new_AGEMA_signal_11534 ), .Q ( new_AGEMA_signal_11535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3513 ( .C ( clk ), .D ( new_AGEMA_signal_11540 ), .Q ( new_AGEMA_signal_11541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3519 ( .C ( clk ), .D ( new_AGEMA_signal_11546 ), .Q ( new_AGEMA_signal_11547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3525 ( .C ( clk ), .D ( new_AGEMA_signal_11552 ), .Q ( new_AGEMA_signal_11553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3529 ( .C ( clk ), .D ( new_AGEMA_signal_11556 ), .Q ( new_AGEMA_signal_11557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3533 ( .C ( clk ), .D ( new_AGEMA_signal_11560 ), .Q ( new_AGEMA_signal_11561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3537 ( .C ( clk ), .D ( new_AGEMA_signal_11564 ), .Q ( new_AGEMA_signal_11565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3541 ( .C ( clk ), .D ( new_AGEMA_signal_11568 ), .Q ( new_AGEMA_signal_11569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3545 ( .C ( clk ), .D ( new_AGEMA_signal_11572 ), .Q ( new_AGEMA_signal_11573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3549 ( .C ( clk ), .D ( new_AGEMA_signal_11576 ), .Q ( new_AGEMA_signal_11577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3553 ( .C ( clk ), .D ( new_AGEMA_signal_11580 ), .Q ( new_AGEMA_signal_11581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3557 ( .C ( clk ), .D ( new_AGEMA_signal_11584 ), .Q ( new_AGEMA_signal_11585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3559 ( .C ( clk ), .D ( n2270 ), .Q ( new_AGEMA_signal_11587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3561 ( .C ( clk ), .D ( new_AGEMA_signal_2274 ), .Q ( new_AGEMA_signal_11589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3563 ( .C ( clk ), .D ( new_AGEMA_signal_2275 ), .Q ( new_AGEMA_signal_11591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3565 ( .C ( clk ), .D ( new_AGEMA_signal_2276 ), .Q ( new_AGEMA_signal_11593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3567 ( .C ( clk ), .D ( n2285 ), .Q ( new_AGEMA_signal_11595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3569 ( .C ( clk ), .D ( new_AGEMA_signal_2700 ), .Q ( new_AGEMA_signal_11597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3571 ( .C ( clk ), .D ( new_AGEMA_signal_2701 ), .Q ( new_AGEMA_signal_11599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3573 ( .C ( clk ), .D ( new_AGEMA_signal_2702 ), .Q ( new_AGEMA_signal_11601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3577 ( .C ( clk ), .D ( new_AGEMA_signal_11604 ), .Q ( new_AGEMA_signal_11605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3581 ( .C ( clk ), .D ( new_AGEMA_signal_11608 ), .Q ( new_AGEMA_signal_11609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3585 ( .C ( clk ), .D ( new_AGEMA_signal_11612 ), .Q ( new_AGEMA_signal_11613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3589 ( .C ( clk ), .D ( new_AGEMA_signal_11616 ), .Q ( new_AGEMA_signal_11617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3593 ( .C ( clk ), .D ( new_AGEMA_signal_11620 ), .Q ( new_AGEMA_signal_11621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3597 ( .C ( clk ), .D ( new_AGEMA_signal_11624 ), .Q ( new_AGEMA_signal_11625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3601 ( .C ( clk ), .D ( new_AGEMA_signal_11628 ), .Q ( new_AGEMA_signal_11629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3605 ( .C ( clk ), .D ( new_AGEMA_signal_11632 ), .Q ( new_AGEMA_signal_11633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3607 ( .C ( clk ), .D ( n2334 ), .Q ( new_AGEMA_signal_11635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3609 ( .C ( clk ), .D ( new_AGEMA_signal_2307 ), .Q ( new_AGEMA_signal_11637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3611 ( .C ( clk ), .D ( new_AGEMA_signal_2308 ), .Q ( new_AGEMA_signal_11639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3613 ( .C ( clk ), .D ( new_AGEMA_signal_2309 ), .Q ( new_AGEMA_signal_11641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3619 ( .C ( clk ), .D ( new_AGEMA_signal_11646 ), .Q ( new_AGEMA_signal_11647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3625 ( .C ( clk ), .D ( new_AGEMA_signal_11652 ), .Q ( new_AGEMA_signal_11653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3631 ( .C ( clk ), .D ( new_AGEMA_signal_11658 ), .Q ( new_AGEMA_signal_11659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3637 ( .C ( clk ), .D ( new_AGEMA_signal_11664 ), .Q ( new_AGEMA_signal_11665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3641 ( .C ( clk ), .D ( new_AGEMA_signal_11668 ), .Q ( new_AGEMA_signal_11669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3645 ( .C ( clk ), .D ( new_AGEMA_signal_11672 ), .Q ( new_AGEMA_signal_11673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3649 ( .C ( clk ), .D ( new_AGEMA_signal_11676 ), .Q ( new_AGEMA_signal_11677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3653 ( .C ( clk ), .D ( new_AGEMA_signal_11680 ), .Q ( new_AGEMA_signal_11681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3655 ( .C ( clk ), .D ( new_AGEMA_signal_10892 ), .Q ( new_AGEMA_signal_11683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3657 ( .C ( clk ), .D ( new_AGEMA_signal_10894 ), .Q ( new_AGEMA_signal_11685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3659 ( .C ( clk ), .D ( new_AGEMA_signal_10896 ), .Q ( new_AGEMA_signal_11687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3661 ( .C ( clk ), .D ( new_AGEMA_signal_10898 ), .Q ( new_AGEMA_signal_11689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3665 ( .C ( clk ), .D ( new_AGEMA_signal_11692 ), .Q ( new_AGEMA_signal_11693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3669 ( .C ( clk ), .D ( new_AGEMA_signal_11696 ), .Q ( new_AGEMA_signal_11697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3673 ( .C ( clk ), .D ( new_AGEMA_signal_11700 ), .Q ( new_AGEMA_signal_11701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3677 ( .C ( clk ), .D ( new_AGEMA_signal_11704 ), .Q ( new_AGEMA_signal_11705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3681 ( .C ( clk ), .D ( new_AGEMA_signal_11708 ), .Q ( new_AGEMA_signal_11709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3685 ( .C ( clk ), .D ( new_AGEMA_signal_11712 ), .Q ( new_AGEMA_signal_11713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3689 ( .C ( clk ), .D ( new_AGEMA_signal_11716 ), .Q ( new_AGEMA_signal_11717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3693 ( .C ( clk ), .D ( new_AGEMA_signal_11720 ), .Q ( new_AGEMA_signal_11721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3697 ( .C ( clk ), .D ( new_AGEMA_signal_11724 ), .Q ( new_AGEMA_signal_11725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3701 ( .C ( clk ), .D ( new_AGEMA_signal_11728 ), .Q ( new_AGEMA_signal_11729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3705 ( .C ( clk ), .D ( new_AGEMA_signal_11732 ), .Q ( new_AGEMA_signal_11733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3709 ( .C ( clk ), .D ( new_AGEMA_signal_11736 ), .Q ( new_AGEMA_signal_11737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3711 ( .C ( clk ), .D ( n2435 ), .Q ( new_AGEMA_signal_11739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3713 ( .C ( clk ), .D ( new_AGEMA_signal_2364 ), .Q ( new_AGEMA_signal_11741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3715 ( .C ( clk ), .D ( new_AGEMA_signal_2365 ), .Q ( new_AGEMA_signal_11743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3717 ( .C ( clk ), .D ( new_AGEMA_signal_2366 ), .Q ( new_AGEMA_signal_11745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3721 ( .C ( clk ), .D ( new_AGEMA_signal_11748 ), .Q ( new_AGEMA_signal_11749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3725 ( .C ( clk ), .D ( new_AGEMA_signal_11752 ), .Q ( new_AGEMA_signal_11753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3729 ( .C ( clk ), .D ( new_AGEMA_signal_11756 ), .Q ( new_AGEMA_signal_11757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3733 ( .C ( clk ), .D ( new_AGEMA_signal_11760 ), .Q ( new_AGEMA_signal_11761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3735 ( .C ( clk ), .D ( new_AGEMA_signal_10740 ), .Q ( new_AGEMA_signal_11763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3737 ( .C ( clk ), .D ( new_AGEMA_signal_10742 ), .Q ( new_AGEMA_signal_11765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3739 ( .C ( clk ), .D ( new_AGEMA_signal_10744 ), .Q ( new_AGEMA_signal_11767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3741 ( .C ( clk ), .D ( new_AGEMA_signal_10746 ), .Q ( new_AGEMA_signal_11769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3747 ( .C ( clk ), .D ( new_AGEMA_signal_11774 ), .Q ( new_AGEMA_signal_11775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3753 ( .C ( clk ), .D ( new_AGEMA_signal_11780 ), .Q ( new_AGEMA_signal_11781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3759 ( .C ( clk ), .D ( new_AGEMA_signal_11786 ), .Q ( new_AGEMA_signal_11787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3765 ( .C ( clk ), .D ( new_AGEMA_signal_11792 ), .Q ( new_AGEMA_signal_11793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3771 ( .C ( clk ), .D ( new_AGEMA_signal_11798 ), .Q ( new_AGEMA_signal_11799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3777 ( .C ( clk ), .D ( new_AGEMA_signal_11804 ), .Q ( new_AGEMA_signal_11805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3783 ( .C ( clk ), .D ( new_AGEMA_signal_11810 ), .Q ( new_AGEMA_signal_11811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3789 ( .C ( clk ), .D ( new_AGEMA_signal_11816 ), .Q ( new_AGEMA_signal_11817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3793 ( .C ( clk ), .D ( new_AGEMA_signal_11820 ), .Q ( new_AGEMA_signal_11821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3797 ( .C ( clk ), .D ( new_AGEMA_signal_11824 ), .Q ( new_AGEMA_signal_11825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3801 ( .C ( clk ), .D ( new_AGEMA_signal_11828 ), .Q ( new_AGEMA_signal_11829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3805 ( .C ( clk ), .D ( new_AGEMA_signal_11832 ), .Q ( new_AGEMA_signal_11833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3807 ( .C ( clk ), .D ( new_AGEMA_signal_10696 ), .Q ( new_AGEMA_signal_11835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3809 ( .C ( clk ), .D ( new_AGEMA_signal_10702 ), .Q ( new_AGEMA_signal_11837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3811 ( .C ( clk ), .D ( new_AGEMA_signal_10708 ), .Q ( new_AGEMA_signal_11839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3813 ( .C ( clk ), .D ( new_AGEMA_signal_10714 ), .Q ( new_AGEMA_signal_11841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3821 ( .C ( clk ), .D ( new_AGEMA_signal_11848 ), .Q ( new_AGEMA_signal_11849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3829 ( .C ( clk ), .D ( new_AGEMA_signal_11856 ), .Q ( new_AGEMA_signal_11857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3837 ( .C ( clk ), .D ( new_AGEMA_signal_11864 ), .Q ( new_AGEMA_signal_11865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3845 ( .C ( clk ), .D ( new_AGEMA_signal_11872 ), .Q ( new_AGEMA_signal_11873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3847 ( .C ( clk ), .D ( n2547 ), .Q ( new_AGEMA_signal_11875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3849 ( .C ( clk ), .D ( new_AGEMA_signal_2418 ), .Q ( new_AGEMA_signal_11877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3851 ( .C ( clk ), .D ( new_AGEMA_signal_2419 ), .Q ( new_AGEMA_signal_11879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3853 ( .C ( clk ), .D ( new_AGEMA_signal_2420 ), .Q ( new_AGEMA_signal_11881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3857 ( .C ( clk ), .D ( new_AGEMA_signal_11884 ), .Q ( new_AGEMA_signal_11885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3861 ( .C ( clk ), .D ( new_AGEMA_signal_11888 ), .Q ( new_AGEMA_signal_11889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3865 ( .C ( clk ), .D ( new_AGEMA_signal_11892 ), .Q ( new_AGEMA_signal_11893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3869 ( .C ( clk ), .D ( new_AGEMA_signal_11896 ), .Q ( new_AGEMA_signal_11897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3873 ( .C ( clk ), .D ( new_AGEMA_signal_11900 ), .Q ( new_AGEMA_signal_11901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3877 ( .C ( clk ), .D ( new_AGEMA_signal_11904 ), .Q ( new_AGEMA_signal_11905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3881 ( .C ( clk ), .D ( new_AGEMA_signal_11908 ), .Q ( new_AGEMA_signal_11909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3885 ( .C ( clk ), .D ( new_AGEMA_signal_11912 ), .Q ( new_AGEMA_signal_11913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3889 ( .C ( clk ), .D ( new_AGEMA_signal_11916 ), .Q ( new_AGEMA_signal_11917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3893 ( .C ( clk ), .D ( new_AGEMA_signal_11920 ), .Q ( new_AGEMA_signal_11921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3897 ( .C ( clk ), .D ( new_AGEMA_signal_11924 ), .Q ( new_AGEMA_signal_11925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3901 ( .C ( clk ), .D ( new_AGEMA_signal_11928 ), .Q ( new_AGEMA_signal_11929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3905 ( .C ( clk ), .D ( new_AGEMA_signal_11932 ), .Q ( new_AGEMA_signal_11933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3909 ( .C ( clk ), .D ( new_AGEMA_signal_11936 ), .Q ( new_AGEMA_signal_11937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3913 ( .C ( clk ), .D ( new_AGEMA_signal_11940 ), .Q ( new_AGEMA_signal_11941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3917 ( .C ( clk ), .D ( new_AGEMA_signal_11944 ), .Q ( new_AGEMA_signal_11945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3921 ( .C ( clk ), .D ( new_AGEMA_signal_11948 ), .Q ( new_AGEMA_signal_11949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3925 ( .C ( clk ), .D ( new_AGEMA_signal_11952 ), .Q ( new_AGEMA_signal_11953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3929 ( .C ( clk ), .D ( new_AGEMA_signal_11956 ), .Q ( new_AGEMA_signal_11957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3933 ( .C ( clk ), .D ( new_AGEMA_signal_11960 ), .Q ( new_AGEMA_signal_11961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3941 ( .C ( clk ), .D ( new_AGEMA_signal_11968 ), .Q ( new_AGEMA_signal_11969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3949 ( .C ( clk ), .D ( new_AGEMA_signal_11976 ), .Q ( new_AGEMA_signal_11977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3957 ( .C ( clk ), .D ( new_AGEMA_signal_11984 ), .Q ( new_AGEMA_signal_11985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3965 ( .C ( clk ), .D ( new_AGEMA_signal_11992 ), .Q ( new_AGEMA_signal_11993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3967 ( .C ( clk ), .D ( n2758 ), .Q ( new_AGEMA_signal_11995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3969 ( .C ( clk ), .D ( new_AGEMA_signal_2853 ), .Q ( new_AGEMA_signal_11997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3971 ( .C ( clk ), .D ( new_AGEMA_signal_2854 ), .Q ( new_AGEMA_signal_11999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3973 ( .C ( clk ), .D ( new_AGEMA_signal_2855 ), .Q ( new_AGEMA_signal_12001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3977 ( .C ( clk ), .D ( new_AGEMA_signal_12004 ), .Q ( new_AGEMA_signal_12005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3981 ( .C ( clk ), .D ( new_AGEMA_signal_12008 ), .Q ( new_AGEMA_signal_12009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3985 ( .C ( clk ), .D ( new_AGEMA_signal_12012 ), .Q ( new_AGEMA_signal_12013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3989 ( .C ( clk ), .D ( new_AGEMA_signal_12016 ), .Q ( new_AGEMA_signal_12017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3991 ( .C ( clk ), .D ( n2797 ), .Q ( new_AGEMA_signal_12019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3993 ( .C ( clk ), .D ( new_AGEMA_signal_2865 ), .Q ( new_AGEMA_signal_12021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3995 ( .C ( clk ), .D ( new_AGEMA_signal_2866 ), .Q ( new_AGEMA_signal_12023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3997 ( .C ( clk ), .D ( new_AGEMA_signal_2867 ), .Q ( new_AGEMA_signal_12025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4003 ( .C ( clk ), .D ( new_AGEMA_signal_12030 ), .Q ( new_AGEMA_signal_12031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4009 ( .C ( clk ), .D ( new_AGEMA_signal_12036 ), .Q ( new_AGEMA_signal_12037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4015 ( .C ( clk ), .D ( new_AGEMA_signal_12042 ), .Q ( new_AGEMA_signal_12043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4021 ( .C ( clk ), .D ( new_AGEMA_signal_12048 ), .Q ( new_AGEMA_signal_12049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4035 ( .C ( clk ), .D ( new_AGEMA_signal_12062 ), .Q ( new_AGEMA_signal_12063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4043 ( .C ( clk ), .D ( new_AGEMA_signal_12070 ), .Q ( new_AGEMA_signal_12071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4051 ( .C ( clk ), .D ( new_AGEMA_signal_12078 ), .Q ( new_AGEMA_signal_12079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4059 ( .C ( clk ), .D ( new_AGEMA_signal_12086 ), .Q ( new_AGEMA_signal_12087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4071 ( .C ( clk ), .D ( n2012 ), .Q ( new_AGEMA_signal_12099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4075 ( .C ( clk ), .D ( new_AGEMA_signal_2577 ), .Q ( new_AGEMA_signal_12103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4079 ( .C ( clk ), .D ( new_AGEMA_signal_2578 ), .Q ( new_AGEMA_signal_12107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4083 ( .C ( clk ), .D ( new_AGEMA_signal_2579 ), .Q ( new_AGEMA_signal_12111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4091 ( .C ( clk ), .D ( new_AGEMA_signal_12118 ), .Q ( new_AGEMA_signal_12119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4099 ( .C ( clk ), .D ( new_AGEMA_signal_12126 ), .Q ( new_AGEMA_signal_12127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4107 ( .C ( clk ), .D ( new_AGEMA_signal_12134 ), .Q ( new_AGEMA_signal_12135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4115 ( .C ( clk ), .D ( new_AGEMA_signal_12142 ), .Q ( new_AGEMA_signal_12143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4129 ( .C ( clk ), .D ( new_AGEMA_signal_12156 ), .Q ( new_AGEMA_signal_12157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4135 ( .C ( clk ), .D ( new_AGEMA_signal_12162 ), .Q ( new_AGEMA_signal_12163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4141 ( .C ( clk ), .D ( new_AGEMA_signal_12168 ), .Q ( new_AGEMA_signal_12169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4147 ( .C ( clk ), .D ( new_AGEMA_signal_12174 ), .Q ( new_AGEMA_signal_12175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4151 ( .C ( clk ), .D ( n2652 ), .Q ( new_AGEMA_signal_12179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4155 ( .C ( clk ), .D ( new_AGEMA_signal_2604 ), .Q ( new_AGEMA_signal_12183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4159 ( .C ( clk ), .D ( new_AGEMA_signal_2605 ), .Q ( new_AGEMA_signal_12187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4163 ( .C ( clk ), .D ( new_AGEMA_signal_2606 ), .Q ( new_AGEMA_signal_12191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4171 ( .C ( clk ), .D ( new_AGEMA_signal_12198 ), .Q ( new_AGEMA_signal_12199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4179 ( .C ( clk ), .D ( new_AGEMA_signal_12206 ), .Q ( new_AGEMA_signal_12207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4187 ( .C ( clk ), .D ( new_AGEMA_signal_12214 ), .Q ( new_AGEMA_signal_12215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4195 ( .C ( clk ), .D ( new_AGEMA_signal_12222 ), .Q ( new_AGEMA_signal_12223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4199 ( .C ( clk ), .D ( n2143 ), .Q ( new_AGEMA_signal_12227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4203 ( .C ( clk ), .D ( new_AGEMA_signal_2640 ), .Q ( new_AGEMA_signal_12231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4207 ( .C ( clk ), .D ( new_AGEMA_signal_2641 ), .Q ( new_AGEMA_signal_12235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4211 ( .C ( clk ), .D ( new_AGEMA_signal_2642 ), .Q ( new_AGEMA_signal_12239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4217 ( .C ( clk ), .D ( new_AGEMA_signal_12244 ), .Q ( new_AGEMA_signal_12245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4223 ( .C ( clk ), .D ( new_AGEMA_signal_12250 ), .Q ( new_AGEMA_signal_12251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4229 ( .C ( clk ), .D ( new_AGEMA_signal_12256 ), .Q ( new_AGEMA_signal_12257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4235 ( .C ( clk ), .D ( new_AGEMA_signal_12262 ), .Q ( new_AGEMA_signal_12263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4241 ( .C ( clk ), .D ( new_AGEMA_signal_12268 ), .Q ( new_AGEMA_signal_12269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4247 ( .C ( clk ), .D ( new_AGEMA_signal_12274 ), .Q ( new_AGEMA_signal_12275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4253 ( .C ( clk ), .D ( new_AGEMA_signal_12280 ), .Q ( new_AGEMA_signal_12281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4259 ( .C ( clk ), .D ( new_AGEMA_signal_12286 ), .Q ( new_AGEMA_signal_12287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4265 ( .C ( clk ), .D ( new_AGEMA_signal_12292 ), .Q ( new_AGEMA_signal_12293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4271 ( .C ( clk ), .D ( new_AGEMA_signal_12298 ), .Q ( new_AGEMA_signal_12299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4277 ( .C ( clk ), .D ( new_AGEMA_signal_12304 ), .Q ( new_AGEMA_signal_12305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4283 ( .C ( clk ), .D ( new_AGEMA_signal_12310 ), .Q ( new_AGEMA_signal_12311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4289 ( .C ( clk ), .D ( new_AGEMA_signal_12316 ), .Q ( new_AGEMA_signal_12317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4295 ( .C ( clk ), .D ( new_AGEMA_signal_12322 ), .Q ( new_AGEMA_signal_12323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4301 ( .C ( clk ), .D ( new_AGEMA_signal_12328 ), .Q ( new_AGEMA_signal_12329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4307 ( .C ( clk ), .D ( new_AGEMA_signal_12334 ), .Q ( new_AGEMA_signal_12335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4313 ( .C ( clk ), .D ( new_AGEMA_signal_12340 ), .Q ( new_AGEMA_signal_12341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4319 ( .C ( clk ), .D ( new_AGEMA_signal_12346 ), .Q ( new_AGEMA_signal_12347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4325 ( .C ( clk ), .D ( new_AGEMA_signal_12352 ), .Q ( new_AGEMA_signal_12353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4331 ( .C ( clk ), .D ( new_AGEMA_signal_12358 ), .Q ( new_AGEMA_signal_12359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4335 ( .C ( clk ), .D ( n2297 ), .Q ( new_AGEMA_signal_12363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4339 ( .C ( clk ), .D ( new_AGEMA_signal_2709 ), .Q ( new_AGEMA_signal_12367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4343 ( .C ( clk ), .D ( new_AGEMA_signal_2710 ), .Q ( new_AGEMA_signal_12371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4347 ( .C ( clk ), .D ( new_AGEMA_signal_2711 ), .Q ( new_AGEMA_signal_12375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4355 ( .C ( clk ), .D ( new_AGEMA_signal_12382 ), .Q ( new_AGEMA_signal_12383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4363 ( .C ( clk ), .D ( new_AGEMA_signal_12390 ), .Q ( new_AGEMA_signal_12391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4371 ( .C ( clk ), .D ( new_AGEMA_signal_12398 ), .Q ( new_AGEMA_signal_12399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4379 ( .C ( clk ), .D ( new_AGEMA_signal_12406 ), .Q ( new_AGEMA_signal_12407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4383 ( .C ( clk ), .D ( n2336 ), .Q ( new_AGEMA_signal_12411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4387 ( .C ( clk ), .D ( new_AGEMA_signal_2994 ), .Q ( new_AGEMA_signal_12415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4391 ( .C ( clk ), .D ( new_AGEMA_signal_2995 ), .Q ( new_AGEMA_signal_12419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4395 ( .C ( clk ), .D ( new_AGEMA_signal_2996 ), .Q ( new_AGEMA_signal_12423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4401 ( .C ( clk ), .D ( new_AGEMA_signal_12428 ), .Q ( new_AGEMA_signal_12429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4407 ( .C ( clk ), .D ( new_AGEMA_signal_12434 ), .Q ( new_AGEMA_signal_12435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4413 ( .C ( clk ), .D ( new_AGEMA_signal_12440 ), .Q ( new_AGEMA_signal_12441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4419 ( .C ( clk ), .D ( new_AGEMA_signal_12446 ), .Q ( new_AGEMA_signal_12447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4427 ( .C ( clk ), .D ( new_AGEMA_signal_12454 ), .Q ( new_AGEMA_signal_12455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4435 ( .C ( clk ), .D ( new_AGEMA_signal_12462 ), .Q ( new_AGEMA_signal_12463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4443 ( .C ( clk ), .D ( new_AGEMA_signal_12470 ), .Q ( new_AGEMA_signal_12471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4451 ( .C ( clk ), .D ( new_AGEMA_signal_12478 ), .Q ( new_AGEMA_signal_12479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4465 ( .C ( clk ), .D ( new_AGEMA_signal_12492 ), .Q ( new_AGEMA_signal_12493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4471 ( .C ( clk ), .D ( new_AGEMA_signal_12498 ), .Q ( new_AGEMA_signal_12499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4477 ( .C ( clk ), .D ( new_AGEMA_signal_12504 ), .Q ( new_AGEMA_signal_12505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4483 ( .C ( clk ), .D ( new_AGEMA_signal_12510 ), .Q ( new_AGEMA_signal_12511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4505 ( .C ( clk ), .D ( new_AGEMA_signal_12532 ), .Q ( new_AGEMA_signal_12533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4511 ( .C ( clk ), .D ( new_AGEMA_signal_12538 ), .Q ( new_AGEMA_signal_12539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4517 ( .C ( clk ), .D ( new_AGEMA_signal_12544 ), .Q ( new_AGEMA_signal_12545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4523 ( .C ( clk ), .D ( new_AGEMA_signal_12550 ), .Q ( new_AGEMA_signal_12551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4529 ( .C ( clk ), .D ( new_AGEMA_signal_12556 ), .Q ( new_AGEMA_signal_12557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4535 ( .C ( clk ), .D ( new_AGEMA_signal_12562 ), .Q ( new_AGEMA_signal_12563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4541 ( .C ( clk ), .D ( new_AGEMA_signal_12568 ), .Q ( new_AGEMA_signal_12569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4547 ( .C ( clk ), .D ( new_AGEMA_signal_12574 ), .Q ( new_AGEMA_signal_12575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4555 ( .C ( clk ), .D ( new_AGEMA_signal_12582 ), .Q ( new_AGEMA_signal_12583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4563 ( .C ( clk ), .D ( new_AGEMA_signal_12590 ), .Q ( new_AGEMA_signal_12591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4571 ( .C ( clk ), .D ( new_AGEMA_signal_12598 ), .Q ( new_AGEMA_signal_12599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4579 ( .C ( clk ), .D ( new_AGEMA_signal_12606 ), .Q ( new_AGEMA_signal_12607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4587 ( .C ( clk ), .D ( new_AGEMA_signal_12614 ), .Q ( new_AGEMA_signal_12615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4595 ( .C ( clk ), .D ( new_AGEMA_signal_12622 ), .Q ( new_AGEMA_signal_12623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4603 ( .C ( clk ), .D ( new_AGEMA_signal_12630 ), .Q ( new_AGEMA_signal_12631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4611 ( .C ( clk ), .D ( new_AGEMA_signal_12638 ), .Q ( new_AGEMA_signal_12639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4617 ( .C ( clk ), .D ( new_AGEMA_signal_12644 ), .Q ( new_AGEMA_signal_12645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4623 ( .C ( clk ), .D ( new_AGEMA_signal_12650 ), .Q ( new_AGEMA_signal_12651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4629 ( .C ( clk ), .D ( new_AGEMA_signal_12656 ), .Q ( new_AGEMA_signal_12657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4635 ( .C ( clk ), .D ( new_AGEMA_signal_12662 ), .Q ( new_AGEMA_signal_12663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4641 ( .C ( clk ), .D ( new_AGEMA_signal_12668 ), .Q ( new_AGEMA_signal_12669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4647 ( .C ( clk ), .D ( new_AGEMA_signal_12674 ), .Q ( new_AGEMA_signal_12675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4653 ( .C ( clk ), .D ( new_AGEMA_signal_12680 ), .Q ( new_AGEMA_signal_12681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4659 ( .C ( clk ), .D ( new_AGEMA_signal_12686 ), .Q ( new_AGEMA_signal_12687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4671 ( .C ( clk ), .D ( n2658 ), .Q ( new_AGEMA_signal_12699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4675 ( .C ( clk ), .D ( new_AGEMA_signal_2550 ), .Q ( new_AGEMA_signal_12703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4679 ( .C ( clk ), .D ( new_AGEMA_signal_2551 ), .Q ( new_AGEMA_signal_12707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4683 ( .C ( clk ), .D ( new_AGEMA_signal_2552 ), .Q ( new_AGEMA_signal_12711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4687 ( .C ( clk ), .D ( n2698 ), .Q ( new_AGEMA_signal_12715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4691 ( .C ( clk ), .D ( new_AGEMA_signal_2835 ), .Q ( new_AGEMA_signal_12719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4695 ( .C ( clk ), .D ( new_AGEMA_signal_2836 ), .Q ( new_AGEMA_signal_12723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4699 ( .C ( clk ), .D ( new_AGEMA_signal_2837 ), .Q ( new_AGEMA_signal_12727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4703 ( .C ( clk ), .D ( n2800 ), .Q ( new_AGEMA_signal_12731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4707 ( .C ( clk ), .D ( new_AGEMA_signal_2859 ), .Q ( new_AGEMA_signal_12735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4711 ( .C ( clk ), .D ( new_AGEMA_signal_2860 ), .Q ( new_AGEMA_signal_12739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4715 ( .C ( clk ), .D ( new_AGEMA_signal_2861 ), .Q ( new_AGEMA_signal_12743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4727 ( .C ( clk ), .D ( n1936 ), .Q ( new_AGEMA_signal_12755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4733 ( .C ( clk ), .D ( new_AGEMA_signal_2526 ), .Q ( new_AGEMA_signal_12761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4739 ( .C ( clk ), .D ( new_AGEMA_signal_2527 ), .Q ( new_AGEMA_signal_12767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4745 ( .C ( clk ), .D ( new_AGEMA_signal_2528 ), .Q ( new_AGEMA_signal_12773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4777 ( .C ( clk ), .D ( new_AGEMA_signal_12804 ), .Q ( new_AGEMA_signal_12805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4785 ( .C ( clk ), .D ( new_AGEMA_signal_12812 ), .Q ( new_AGEMA_signal_12813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4793 ( .C ( clk ), .D ( new_AGEMA_signal_12820 ), .Q ( new_AGEMA_signal_12821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4801 ( .C ( clk ), .D ( new_AGEMA_signal_12828 ), .Q ( new_AGEMA_signal_12829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4809 ( .C ( clk ), .D ( new_AGEMA_signal_12836 ), .Q ( new_AGEMA_signal_12837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4817 ( .C ( clk ), .D ( new_AGEMA_signal_12844 ), .Q ( new_AGEMA_signal_12845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4825 ( .C ( clk ), .D ( new_AGEMA_signal_12852 ), .Q ( new_AGEMA_signal_12853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4833 ( .C ( clk ), .D ( new_AGEMA_signal_12860 ), .Q ( new_AGEMA_signal_12861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4841 ( .C ( clk ), .D ( new_AGEMA_signal_12868 ), .Q ( new_AGEMA_signal_12869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4849 ( .C ( clk ), .D ( new_AGEMA_signal_12876 ), .Q ( new_AGEMA_signal_12877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4857 ( .C ( clk ), .D ( new_AGEMA_signal_12884 ), .Q ( new_AGEMA_signal_12885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4865 ( .C ( clk ), .D ( new_AGEMA_signal_12892 ), .Q ( new_AGEMA_signal_12893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4873 ( .C ( clk ), .D ( new_AGEMA_signal_12900 ), .Q ( new_AGEMA_signal_12901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4881 ( .C ( clk ), .D ( new_AGEMA_signal_12908 ), .Q ( new_AGEMA_signal_12909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4889 ( .C ( clk ), .D ( new_AGEMA_signal_12916 ), .Q ( new_AGEMA_signal_12917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4897 ( .C ( clk ), .D ( new_AGEMA_signal_12924 ), .Q ( new_AGEMA_signal_12925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4903 ( .C ( clk ), .D ( n2099 ), .Q ( new_AGEMA_signal_12931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4909 ( .C ( clk ), .D ( new_AGEMA_signal_2613 ), .Q ( new_AGEMA_signal_12937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4915 ( .C ( clk ), .D ( new_AGEMA_signal_2614 ), .Q ( new_AGEMA_signal_12943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4921 ( .C ( clk ), .D ( new_AGEMA_signal_2615 ), .Q ( new_AGEMA_signal_12949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4931 ( .C ( clk ), .D ( new_AGEMA_signal_12958 ), .Q ( new_AGEMA_signal_12959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4941 ( .C ( clk ), .D ( new_AGEMA_signal_12968 ), .Q ( new_AGEMA_signal_12969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4951 ( .C ( clk ), .D ( new_AGEMA_signal_12978 ), .Q ( new_AGEMA_signal_12979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4961 ( .C ( clk ), .D ( new_AGEMA_signal_12988 ), .Q ( new_AGEMA_signal_12989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4969 ( .C ( clk ), .D ( new_AGEMA_signal_12996 ), .Q ( new_AGEMA_signal_12997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4977 ( .C ( clk ), .D ( new_AGEMA_signal_13004 ), .Q ( new_AGEMA_signal_13005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4985 ( .C ( clk ), .D ( new_AGEMA_signal_13012 ), .Q ( new_AGEMA_signal_13013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4993 ( .C ( clk ), .D ( new_AGEMA_signal_13020 ), .Q ( new_AGEMA_signal_13021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5001 ( .C ( clk ), .D ( new_AGEMA_signal_13028 ), .Q ( new_AGEMA_signal_13029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5009 ( .C ( clk ), .D ( new_AGEMA_signal_13036 ), .Q ( new_AGEMA_signal_13037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5017 ( .C ( clk ), .D ( new_AGEMA_signal_13044 ), .Q ( new_AGEMA_signal_13045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5025 ( .C ( clk ), .D ( new_AGEMA_signal_13052 ), .Q ( new_AGEMA_signal_13053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5033 ( .C ( clk ), .D ( new_AGEMA_signal_13060 ), .Q ( new_AGEMA_signal_13061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5041 ( .C ( clk ), .D ( new_AGEMA_signal_13068 ), .Q ( new_AGEMA_signal_13069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5049 ( .C ( clk ), .D ( new_AGEMA_signal_13076 ), .Q ( new_AGEMA_signal_13077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5057 ( .C ( clk ), .D ( new_AGEMA_signal_13084 ), .Q ( new_AGEMA_signal_13085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5087 ( .C ( clk ), .D ( n2301 ), .Q ( new_AGEMA_signal_13115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5093 ( .C ( clk ), .D ( new_AGEMA_signal_2715 ), .Q ( new_AGEMA_signal_13121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5099 ( .C ( clk ), .D ( new_AGEMA_signal_2716 ), .Q ( new_AGEMA_signal_13127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5105 ( .C ( clk ), .D ( new_AGEMA_signal_2717 ), .Q ( new_AGEMA_signal_13133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5131 ( .C ( clk ), .D ( new_AGEMA_signal_13158 ), .Q ( new_AGEMA_signal_13159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5141 ( .C ( clk ), .D ( new_AGEMA_signal_13168 ), .Q ( new_AGEMA_signal_13169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5151 ( .C ( clk ), .D ( new_AGEMA_signal_13178 ), .Q ( new_AGEMA_signal_13179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5161 ( .C ( clk ), .D ( new_AGEMA_signal_13188 ), .Q ( new_AGEMA_signal_13189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5169 ( .C ( clk ), .D ( new_AGEMA_signal_13196 ), .Q ( new_AGEMA_signal_13197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5177 ( .C ( clk ), .D ( new_AGEMA_signal_13204 ), .Q ( new_AGEMA_signal_13205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5185 ( .C ( clk ), .D ( new_AGEMA_signal_13212 ), .Q ( new_AGEMA_signal_13213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C ( clk ), .D ( new_AGEMA_signal_13220 ), .Q ( new_AGEMA_signal_13221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C ( clk ), .D ( new_AGEMA_signal_13252 ), .Q ( new_AGEMA_signal_13253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C ( clk ), .D ( new_AGEMA_signal_13260 ), .Q ( new_AGEMA_signal_13261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C ( clk ), .D ( new_AGEMA_signal_13268 ), .Q ( new_AGEMA_signal_13269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C ( clk ), .D ( new_AGEMA_signal_13276 ), .Q ( new_AGEMA_signal_13277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5257 ( .C ( clk ), .D ( new_AGEMA_signal_13284 ), .Q ( new_AGEMA_signal_13285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5265 ( .C ( clk ), .D ( new_AGEMA_signal_13292 ), .Q ( new_AGEMA_signal_13293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5273 ( .C ( clk ), .D ( new_AGEMA_signal_13300 ), .Q ( new_AGEMA_signal_13301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5281 ( .C ( clk ), .D ( new_AGEMA_signal_13308 ), .Q ( new_AGEMA_signal_13309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5287 ( .C ( clk ), .D ( new_AGEMA_signal_10630 ), .Q ( new_AGEMA_signal_13315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5293 ( .C ( clk ), .D ( new_AGEMA_signal_10634 ), .Q ( new_AGEMA_signal_13321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5299 ( .C ( clk ), .D ( new_AGEMA_signal_10638 ), .Q ( new_AGEMA_signal_13327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5305 ( .C ( clk ), .D ( new_AGEMA_signal_10642 ), .Q ( new_AGEMA_signal_13333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5329 ( .C ( clk ), .D ( new_AGEMA_signal_13356 ), .Q ( new_AGEMA_signal_13357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5337 ( .C ( clk ), .D ( new_AGEMA_signal_13364 ), .Q ( new_AGEMA_signal_13365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5345 ( .C ( clk ), .D ( new_AGEMA_signal_13372 ), .Q ( new_AGEMA_signal_13373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5353 ( .C ( clk ), .D ( new_AGEMA_signal_13380 ), .Q ( new_AGEMA_signal_13381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5455 ( .C ( clk ), .D ( new_AGEMA_signal_11078 ), .Q ( new_AGEMA_signal_13483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5463 ( .C ( clk ), .D ( new_AGEMA_signal_11082 ), .Q ( new_AGEMA_signal_13491 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5471 ( .C ( clk ), .D ( new_AGEMA_signal_11086 ), .Q ( new_AGEMA_signal_13499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5479 ( .C ( clk ), .D ( new_AGEMA_signal_11090 ), .Q ( new_AGEMA_signal_13507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5527 ( .C ( clk ), .D ( n2102 ), .Q ( new_AGEMA_signal_13555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5535 ( .C ( clk ), .D ( new_AGEMA_signal_2625 ), .Q ( new_AGEMA_signal_13563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5543 ( .C ( clk ), .D ( new_AGEMA_signal_2626 ), .Q ( new_AGEMA_signal_13571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5551 ( .C ( clk ), .D ( new_AGEMA_signal_2627 ), .Q ( new_AGEMA_signal_13579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5559 ( .C ( clk ), .D ( new_AGEMA_signal_10468 ), .Q ( new_AGEMA_signal_13587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5567 ( .C ( clk ), .D ( new_AGEMA_signal_10470 ), .Q ( new_AGEMA_signal_13595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5575 ( .C ( clk ), .D ( new_AGEMA_signal_10472 ), .Q ( new_AGEMA_signal_13603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5583 ( .C ( clk ), .D ( new_AGEMA_signal_10474 ), .Q ( new_AGEMA_signal_13611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5593 ( .C ( clk ), .D ( new_AGEMA_signal_13620 ), .Q ( new_AGEMA_signal_13621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5603 ( .C ( clk ), .D ( new_AGEMA_signal_13630 ), .Q ( new_AGEMA_signal_13631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5613 ( .C ( clk ), .D ( new_AGEMA_signal_13640 ), .Q ( new_AGEMA_signal_13641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5623 ( .C ( clk ), .D ( new_AGEMA_signal_13650 ), .Q ( new_AGEMA_signal_13651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5631 ( .C ( clk ), .D ( new_AGEMA_signal_10838 ), .Q ( new_AGEMA_signal_13659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5639 ( .C ( clk ), .D ( new_AGEMA_signal_10842 ), .Q ( new_AGEMA_signal_13667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5647 ( .C ( clk ), .D ( new_AGEMA_signal_10846 ), .Q ( new_AGEMA_signal_13675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5655 ( .C ( clk ), .D ( new_AGEMA_signal_10850 ), .Q ( new_AGEMA_signal_13683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5727 ( .C ( clk ), .D ( n2367 ), .Q ( new_AGEMA_signal_13755 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5735 ( .C ( clk ), .D ( new_AGEMA_signal_2316 ), .Q ( new_AGEMA_signal_13763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5743 ( .C ( clk ), .D ( new_AGEMA_signal_2317 ), .Q ( new_AGEMA_signal_13771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5751 ( .C ( clk ), .D ( new_AGEMA_signal_2318 ), .Q ( new_AGEMA_signal_13779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5791 ( .C ( clk ), .D ( n2591 ), .Q ( new_AGEMA_signal_13819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5799 ( .C ( clk ), .D ( new_AGEMA_signal_2808 ), .Q ( new_AGEMA_signal_13827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5807 ( .C ( clk ), .D ( new_AGEMA_signal_2809 ), .Q ( new_AGEMA_signal_13835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5815 ( .C ( clk ), .D ( new_AGEMA_signal_2810 ), .Q ( new_AGEMA_signal_13843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5967 ( .C ( clk ), .D ( n2105 ), .Q ( new_AGEMA_signal_13995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5977 ( .C ( clk ), .D ( new_AGEMA_signal_2610 ), .Q ( new_AGEMA_signal_14005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5987 ( .C ( clk ), .D ( new_AGEMA_signal_2611 ), .Q ( new_AGEMA_signal_14015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5997 ( .C ( clk ), .D ( new_AGEMA_signal_2612 ), .Q ( new_AGEMA_signal_14025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6327 ( .C ( clk ), .D ( n2106 ), .Q ( new_AGEMA_signal_14355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6339 ( .C ( clk ), .D ( new_AGEMA_signal_2187 ), .Q ( new_AGEMA_signal_14367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6351 ( .C ( clk ), .D ( new_AGEMA_signal_2188 ), .Q ( new_AGEMA_signal_14379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6363 ( .C ( clk ), .D ( new_AGEMA_signal_2189 ), .Q ( new_AGEMA_signal_14391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6377 ( .C ( clk ), .D ( new_AGEMA_signal_14404 ), .Q ( new_AGEMA_signal_14405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6391 ( .C ( clk ), .D ( new_AGEMA_signal_14418 ), .Q ( new_AGEMA_signal_14419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6405 ( .C ( clk ), .D ( new_AGEMA_signal_14432 ), .Q ( new_AGEMA_signal_14433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6419 ( .C ( clk ), .D ( new_AGEMA_signal_14446 ), .Q ( new_AGEMA_signal_14447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6465 ( .C ( clk ), .D ( new_AGEMA_signal_14492 ), .Q ( new_AGEMA_signal_14493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6479 ( .C ( clk ), .D ( new_AGEMA_signal_14506 ), .Q ( new_AGEMA_signal_14507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6493 ( .C ( clk ), .D ( new_AGEMA_signal_14520 ), .Q ( new_AGEMA_signal_14521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6507 ( .C ( clk ), .D ( new_AGEMA_signal_14534 ), .Q ( new_AGEMA_signal_14535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6609 ( .C ( clk ), .D ( new_AGEMA_signal_14636 ), .Q ( new_AGEMA_signal_14637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6625 ( .C ( clk ), .D ( new_AGEMA_signal_14652 ), .Q ( new_AGEMA_signal_14653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6641 ( .C ( clk ), .D ( new_AGEMA_signal_14668 ), .Q ( new_AGEMA_signal_14669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6657 ( .C ( clk ), .D ( new_AGEMA_signal_14684 ), .Q ( new_AGEMA_signal_14685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6697 ( .C ( clk ), .D ( new_AGEMA_signal_14724 ), .Q ( new_AGEMA_signal_14725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6713 ( .C ( clk ), .D ( new_AGEMA_signal_14740 ), .Q ( new_AGEMA_signal_14741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6729 ( .C ( clk ), .D ( new_AGEMA_signal_14756 ), .Q ( new_AGEMA_signal_14757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6745 ( .C ( clk ), .D ( new_AGEMA_signal_14772 ), .Q ( new_AGEMA_signal_14773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6895 ( .C ( clk ), .D ( n2155 ), .Q ( new_AGEMA_signal_14923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6911 ( .C ( clk ), .D ( new_AGEMA_signal_2193 ), .Q ( new_AGEMA_signal_14939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6927 ( .C ( clk ), .D ( new_AGEMA_signal_2194 ), .Q ( new_AGEMA_signal_14955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6943 ( .C ( clk ), .D ( new_AGEMA_signal_2195 ), .Q ( new_AGEMA_signal_14971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7001 ( .C ( clk ), .D ( new_AGEMA_signal_15028 ), .Q ( new_AGEMA_signal_15029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7019 ( .C ( clk ), .D ( new_AGEMA_signal_15046 ), .Q ( new_AGEMA_signal_15047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7037 ( .C ( clk ), .D ( new_AGEMA_signal_15064 ), .Q ( new_AGEMA_signal_15065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7055 ( .C ( clk ), .D ( new_AGEMA_signal_15082 ), .Q ( new_AGEMA_signal_15083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7201 ( .C ( clk ), .D ( new_AGEMA_signal_15228 ), .Q ( new_AGEMA_signal_15229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7221 ( .C ( clk ), .D ( new_AGEMA_signal_15248 ), .Q ( new_AGEMA_signal_15249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7241 ( .C ( clk ), .D ( new_AGEMA_signal_15268 ), .Q ( new_AGEMA_signal_15269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7261 ( .C ( clk ), .D ( new_AGEMA_signal_15288 ), .Q ( new_AGEMA_signal_15289 ) ) ;

    /* cells in depth 10 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1983 ( .a ({new_AGEMA_signal_10330, new_AGEMA_signal_10326, new_AGEMA_signal_10322, new_AGEMA_signal_10318}), .b ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, n1928}), .clk ( clk ), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, n1934}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U1998 ( .a ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, n1931}), .b ({new_AGEMA_signal_10346, new_AGEMA_signal_10342, new_AGEMA_signal_10338, new_AGEMA_signal_10334}), .clk ( clk ), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n1932}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2015 ( .a ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, n1939}), .b ({new_AGEMA_signal_10354, new_AGEMA_signal_10352, new_AGEMA_signal_10350, new_AGEMA_signal_10348}), .clk ( clk ), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, n1940}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2033 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, n1948}), .b ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, n1947}), .clk ( clk ), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, n1961}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2050 ( .a ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, n1954}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, n1953}), .clk ( clk ), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, n1955}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2066 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10360, new_AGEMA_signal_10358, new_AGEMA_signal_10356}), .b ({new_AGEMA_signal_2084, new_AGEMA_signal_2083, new_AGEMA_signal_2082, n1965}), .clk ( clk ), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, n1967}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2085 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, n1970}), .b ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, n1969}), .clk ( clk ), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, n1984}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2103 ( .a ({new_AGEMA_signal_10378, new_AGEMA_signal_10374, new_AGEMA_signal_10370, new_AGEMA_signal_10366}), .b ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, n1975}), .clk ( clk ), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, n1977}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2108 ( .a ({new_AGEMA_signal_10386, new_AGEMA_signal_10384, new_AGEMA_signal_10382, new_AGEMA_signal_10380}), .b ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, n1980}), .clk ( clk ), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, n1981}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2115 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10398, new_AGEMA_signal_10394, new_AGEMA_signal_10390}), .b ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, n1986}), .clk ( clk ), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, n1987}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2127 ( .a ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, n1997}), .b ({new_AGEMA_signal_10410, new_AGEMA_signal_10408, new_AGEMA_signal_10406, new_AGEMA_signal_10404}), .clk ( clk ), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n1998}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2146 ( .a ({new_AGEMA_signal_10426, new_AGEMA_signal_10422, new_AGEMA_signal_10418, new_AGEMA_signal_10414}), .b ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, n2007}), .clk ( clk ), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, n2010}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2162 ( .a ({new_AGEMA_signal_10442, new_AGEMA_signal_10438, new_AGEMA_signal_10434, new_AGEMA_signal_10430}), .b ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, n2021}), .clk ( clk ), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, n2024}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2177 ( .a ({new_AGEMA_signal_10450, new_AGEMA_signal_10448, new_AGEMA_signal_10446, new_AGEMA_signal_10444}), .b ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, n2032}), .clk ( clk ), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, n2035}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2186 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, n2041}), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10456, new_AGEMA_signal_10454, new_AGEMA_signal_10452}), .clk ( clk ), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, n2054}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2190 ( .a ({new_AGEMA_signal_10466, new_AGEMA_signal_10464, new_AGEMA_signal_10462, new_AGEMA_signal_10460}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, n2043}), .clk ( clk ), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, n2048}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2195 ( .a ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, n2046}), .b ({new_AGEMA_signal_10474, new_AGEMA_signal_10472, new_AGEMA_signal_10470, new_AGEMA_signal_10468}), .clk ( clk ), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, n2047}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2206 ( .a ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, n2058}), .b ({new_AGEMA_signal_10490, new_AGEMA_signal_10486, new_AGEMA_signal_10482, new_AGEMA_signal_10478}), .clk ( clk ), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, n2059}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2213 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, n2063}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10502, new_AGEMA_signal_10498, new_AGEMA_signal_10494}), .clk ( clk ), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2064}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2229 ( .a ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, n2076}), .b ({new_AGEMA_signal_10522, new_AGEMA_signal_10518, new_AGEMA_signal_10514, new_AGEMA_signal_10510}), .clk ( clk ), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, n2077}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2249 ( .a ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, n2090}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10528, new_AGEMA_signal_10526, new_AGEMA_signal_10524}), .clk ( clk ), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2255 ( .a ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, n2093}), .b ({new_AGEMA_signal_10538, new_AGEMA_signal_10536, new_AGEMA_signal_10534, new_AGEMA_signal_10532}), .clk ( clk ), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, n2095}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2274 ( .a ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, n2116}), .b ({new_AGEMA_signal_10546, new_AGEMA_signal_10544, new_AGEMA_signal_10542, new_AGEMA_signal_10540}), .clk ( clk ), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, n2117}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2283 ( .a ({new_AGEMA_signal_10562, new_AGEMA_signal_10558, new_AGEMA_signal_10554, new_AGEMA_signal_10550}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, n2120}), .clk ( clk ), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, n2123}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2300 ( .a ({new_AGEMA_signal_10570, new_AGEMA_signal_10568, new_AGEMA_signal_10566, new_AGEMA_signal_10564}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, n2134}), .clk ( clk ), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, n2135}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2309 ( .a ({new_AGEMA_signal_10586, new_AGEMA_signal_10582, new_AGEMA_signal_10578, new_AGEMA_signal_10574}), .b ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, n2140}), .clk ( clk ), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, n2141}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2327 ( .a ({new_AGEMA_signal_10610, new_AGEMA_signal_10604, new_AGEMA_signal_10598, new_AGEMA_signal_10592}), .b ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, n2161}), .clk ( clk ), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2166}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2331 ( .a ({new_AGEMA_signal_10626, new_AGEMA_signal_10622, new_AGEMA_signal_10618, new_AGEMA_signal_10614}), .b ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, n2164}), .clk ( clk ), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2165}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2346 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, n2179}), .b ({new_AGEMA_signal_10642, new_AGEMA_signal_10638, new_AGEMA_signal_10634, new_AGEMA_signal_10630}), .clk ( clk ), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, n2180}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2360 ( .a ({new_AGEMA_signal_10650, new_AGEMA_signal_10648, new_AGEMA_signal_10646, new_AGEMA_signal_10644}), .b ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, n2192}), .clk ( clk ), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, n2194}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2372 ( .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, n2203}), .b ({new_AGEMA_signal_10658, new_AGEMA_signal_10656, new_AGEMA_signal_10654, new_AGEMA_signal_10652}), .clk ( clk ), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, n2204}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2389 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, n2224}), .b ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, n2223}), .clk ( clk ), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2225}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2394 ( .a ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, n2229}), .b ({new_AGEMA_signal_10666, new_AGEMA_signal_10664, new_AGEMA_signal_10662, new_AGEMA_signal_10660}), .clk ( clk ), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, n2230}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2400 ( .a ({new_AGEMA_signal_10674, new_AGEMA_signal_10672, new_AGEMA_signal_10670, new_AGEMA_signal_10668}), .b ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, n2234}), .clk ( clk ), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2236}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2412 ( .a ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, n2246}), .b ({new_AGEMA_signal_10690, new_AGEMA_signal_10686, new_AGEMA_signal_10682, new_AGEMA_signal_10678}), .clk ( clk ), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, n2247}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2419 ( .a ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, n2254}), .b ({new_AGEMA_signal_10714, new_AGEMA_signal_10708, new_AGEMA_signal_10702, new_AGEMA_signal_10696}), .clk ( clk ), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, n2255}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2427 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, n2263}), .b ({new_AGEMA_signal_10730, new_AGEMA_signal_10726, new_AGEMA_signal_10722, new_AGEMA_signal_10718}), .clk ( clk ), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, n2264}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2435 ( .a ({new_AGEMA_signal_10738, new_AGEMA_signal_10736, new_AGEMA_signal_10734, new_AGEMA_signal_10732}), .b ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, n2267}), .clk ( clk ), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, n2271}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2446 ( .a ({new_AGEMA_signal_10402, new_AGEMA_signal_10398, new_AGEMA_signal_10394, new_AGEMA_signal_10390}), .b ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, n2279}), .clk ( clk ), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, n2280}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2451 ( .a ({new_AGEMA_signal_10746, new_AGEMA_signal_10744, new_AGEMA_signal_10742, new_AGEMA_signal_10740}), .b ({new_AGEMA_signal_2282, new_AGEMA_signal_2281, new_AGEMA_signal_2280, n2283}), .clk ( clk ), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, n2286}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2461 ( .a ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}), .b ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, n2289}), .clk ( clk ), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, n2304}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2466 ( .a ({new_AGEMA_signal_10754, new_AGEMA_signal_10752, new_AGEMA_signal_10750, new_AGEMA_signal_10748}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, n2292}), .clk ( clk ), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, n2295}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2488 ( .a ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, n2321}), .b ({new_AGEMA_signal_1817, new_AGEMA_signal_1816, new_AGEMA_signal_1815, n2320}), .clk ( clk ), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, n2322}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2499 ( .a ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, n2332}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, n2331}), .clk ( clk ), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, n2333}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2509 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10766, new_AGEMA_signal_10762, new_AGEMA_signal_10758}), .b ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, n2342}), .clk ( clk ), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, n2345}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2526 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, n2358}), .b ({new_AGEMA_signal_10778, new_AGEMA_signal_10776, new_AGEMA_signal_10774, new_AGEMA_signal_10772}), .clk ( clk ), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, n2361}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2549 ( .a ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, n2387}), .b ({new_AGEMA_signal_10786, new_AGEMA_signal_10784, new_AGEMA_signal_10782, new_AGEMA_signal_10780}), .clk ( clk ), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, n2388}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2556 ( .a ({new_AGEMA_signal_10802, new_AGEMA_signal_10798, new_AGEMA_signal_10794, new_AGEMA_signal_10790}), .b ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, n2392}), .clk ( clk ), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2393}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2567 ( .a ({new_AGEMA_signal_10818, new_AGEMA_signal_10814, new_AGEMA_signal_10810, new_AGEMA_signal_10806}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, n2404}), .clk ( clk ), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, n2405}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2571 ( .a ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, n2409}), .b ({new_AGEMA_signal_10834, new_AGEMA_signal_10830, new_AGEMA_signal_10826, new_AGEMA_signal_10822}), .clk ( clk ), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, n2410}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2576 ( .a ({new_AGEMA_signal_10850, new_AGEMA_signal_10846, new_AGEMA_signal_10842, new_AGEMA_signal_10838}), .b ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, n2414}), .clk ( clk ), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, n2421}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2579 ( .a ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, n2418}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10862, new_AGEMA_signal_10858, new_AGEMA_signal_10854}), .clk ( clk ), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2419}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2590 ( .a ({new_AGEMA_signal_10874, new_AGEMA_signal_10872, new_AGEMA_signal_10870, new_AGEMA_signal_10868}), .b ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, n2432}), .clk ( clk ), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, n2436}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2604 ( .a ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, n2449}), .b ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, n2448}), .clk ( clk ), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, n2450}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2610 ( .a ({new_AGEMA_signal_10882, new_AGEMA_signal_10880, new_AGEMA_signal_10878, new_AGEMA_signal_10876}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, n2455}), .clk ( clk ), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, n2456}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2613 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, n2460}), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10888, new_AGEMA_signal_10886, new_AGEMA_signal_10884}), .clk ( clk ), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2461}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2619 ( .a ({new_AGEMA_signal_10898, new_AGEMA_signal_10896, new_AGEMA_signal_10894, new_AGEMA_signal_10892}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, n2466}), .clk ( clk ), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, n2469}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2630 ( .a ({new_AGEMA_signal_10914, new_AGEMA_signal_10910, new_AGEMA_signal_10906, new_AGEMA_signal_10902}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, n2477}), .clk ( clk ), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, n2478}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2635 ( .a ({new_AGEMA_signal_10930, new_AGEMA_signal_10926, new_AGEMA_signal_10922, new_AGEMA_signal_10918}), .b ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, n2482}), .clk ( clk ), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, n2484}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2643 ( .a ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, n2490}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10936, new_AGEMA_signal_10934, new_AGEMA_signal_10932}), .clk ( clk ), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, n2491}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2649 ( .a ({new_AGEMA_signal_10946, new_AGEMA_signal_10944, new_AGEMA_signal_10942, new_AGEMA_signal_10940}), .b ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, n2496}), .clk ( clk ), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2500}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2656 ( .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, n2507}), .b ({new_AGEMA_signal_10954, new_AGEMA_signal_10952, new_AGEMA_signal_10950, new_AGEMA_signal_10948}), .clk ( clk ), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, n2508}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2670 ( .a ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, n2525}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, n2524}), .clk ( clk ), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, n2526}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2679 ( .a ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, n2537}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, n2536}), .clk ( clk ), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, n2539}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2682 ( .a ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, n2543}), .b ({new_AGEMA_signal_10962, new_AGEMA_signal_10960, new_AGEMA_signal_10958, new_AGEMA_signal_10956}), .clk ( clk ), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n2548}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2694 ( .a ({new_AGEMA_signal_10970, new_AGEMA_signal_10968, new_AGEMA_signal_10966, new_AGEMA_signal_10964}), .b ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, n2557}), .clk ( clk ), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, n2568}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2700 ( .a ({new_AGEMA_signal_10978, new_AGEMA_signal_10976, new_AGEMA_signal_10974, new_AGEMA_signal_10972}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, n2565}), .clk ( clk ), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, n2567}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2710 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10984, new_AGEMA_signal_10982, new_AGEMA_signal_10980}), .b ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, n2580}), .clk ( clk ), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, n2583}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2728 ( .a ({new_AGEMA_signal_10994, new_AGEMA_signal_10992, new_AGEMA_signal_10990, new_AGEMA_signal_10988}), .b ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, n2602}), .clk ( clk ), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2604}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2739 ( .a ({new_AGEMA_signal_11002, new_AGEMA_signal_11000, new_AGEMA_signal_10998, new_AGEMA_signal_10996}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, n2619}), .clk ( clk ), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, n2621}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2745 ( .a ({new_AGEMA_signal_11018, new_AGEMA_signal_11014, new_AGEMA_signal_11010, new_AGEMA_signal_11006}), .b ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, n2628}), .clk ( clk ), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, n2633}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2756 ( .a ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, n2649}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, n2648}), .clk ( clk ), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, n2660}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2759 ( .a ({new_AGEMA_signal_11026, new_AGEMA_signal_11024, new_AGEMA_signal_11022, new_AGEMA_signal_11020}), .b ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, n2652}), .clk ( clk ), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n2656}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2766 ( .a ({new_AGEMA_signal_11034, new_AGEMA_signal_11032, new_AGEMA_signal_11030, new_AGEMA_signal_11028}), .b ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, n2664}), .clk ( clk ), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, n2666}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2774 ( .a ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, n2681}), .b ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, n2680}), .clk ( clk ), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, n2706}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2777 ( .a ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, n2686}), .b ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, n2685}), .clk ( clk ), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, n2704}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2781 ( .a ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, n2692}), .b ({new_AGEMA_signal_11042, new_AGEMA_signal_11040, new_AGEMA_signal_11038, new_AGEMA_signal_11036}), .clk ( clk ), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n2696}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2794 ( .a ({new_AGEMA_signal_11050, new_AGEMA_signal_11048, new_AGEMA_signal_11046, new_AGEMA_signal_11044}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, n2716}), .clk ( clk ), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, n2718}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2801 ( .a ({new_AGEMA_signal_11058, new_AGEMA_signal_11056, new_AGEMA_signal_11054, new_AGEMA_signal_11052}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, n2728}), .clk ( clk ), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, n2730}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2805 ( .a ({new_AGEMA_signal_11074, new_AGEMA_signal_11070, new_AGEMA_signal_11066, new_AGEMA_signal_11062}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, n2735}), .clk ( clk ), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, n2745}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2809 ( .a ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, n2743}), .b ({new_AGEMA_signal_11090, new_AGEMA_signal_11086, new_AGEMA_signal_11082, new_AGEMA_signal_11078}), .clk ( clk ), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n2744}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2814 ( .a ({new_AGEMA_signal_10738, new_AGEMA_signal_10736, new_AGEMA_signal_10734, new_AGEMA_signal_10732}), .b ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, n2751}), .clk ( clk ), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, n2759}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2821 ( .a ({new_AGEMA_signal_11106, new_AGEMA_signal_11102, new_AGEMA_signal_11098, new_AGEMA_signal_11094}), .b ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, n2764}), .clk ( clk ), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, n2771}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2833 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, n2788}), .b ({new_AGEMA_signal_11122, new_AGEMA_signal_11118, new_AGEMA_signal_11114, new_AGEMA_signal_11110}), .clk ( clk ), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2798}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2850 ( .a ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, n2822}), .b ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, n2821}), .clk ( clk ), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n2826}) ) ;
    buf_clk new_AGEMA_reg_buffer_3098 ( .C ( clk ), .D ( new_AGEMA_signal_11125 ), .Q ( new_AGEMA_signal_11126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3102 ( .C ( clk ), .D ( new_AGEMA_signal_11129 ), .Q ( new_AGEMA_signal_11130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3106 ( .C ( clk ), .D ( new_AGEMA_signal_11133 ), .Q ( new_AGEMA_signal_11134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3110 ( .C ( clk ), .D ( new_AGEMA_signal_11137 ), .Q ( new_AGEMA_signal_11138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3114 ( .C ( clk ), .D ( new_AGEMA_signal_11141 ), .Q ( new_AGEMA_signal_11142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3118 ( .C ( clk ), .D ( new_AGEMA_signal_11145 ), .Q ( new_AGEMA_signal_11146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3122 ( .C ( clk ), .D ( new_AGEMA_signal_11149 ), .Q ( new_AGEMA_signal_11150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3126 ( .C ( clk ), .D ( new_AGEMA_signal_11153 ), .Q ( new_AGEMA_signal_11154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3134 ( .C ( clk ), .D ( new_AGEMA_signal_11161 ), .Q ( new_AGEMA_signal_11162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3142 ( .C ( clk ), .D ( new_AGEMA_signal_11169 ), .Q ( new_AGEMA_signal_11170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3150 ( .C ( clk ), .D ( new_AGEMA_signal_11177 ), .Q ( new_AGEMA_signal_11178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3158 ( .C ( clk ), .D ( new_AGEMA_signal_11185 ), .Q ( new_AGEMA_signal_11186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3160 ( .C ( clk ), .D ( new_AGEMA_signal_11187 ), .Q ( new_AGEMA_signal_11188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3162 ( .C ( clk ), .D ( new_AGEMA_signal_11189 ), .Q ( new_AGEMA_signal_11190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3164 ( .C ( clk ), .D ( new_AGEMA_signal_11191 ), .Q ( new_AGEMA_signal_11192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3166 ( .C ( clk ), .D ( new_AGEMA_signal_11193 ), .Q ( new_AGEMA_signal_11194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3174 ( .C ( clk ), .D ( new_AGEMA_signal_11201 ), .Q ( new_AGEMA_signal_11202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3182 ( .C ( clk ), .D ( new_AGEMA_signal_11209 ), .Q ( new_AGEMA_signal_11210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3190 ( .C ( clk ), .D ( new_AGEMA_signal_11217 ), .Q ( new_AGEMA_signal_11218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3198 ( .C ( clk ), .D ( new_AGEMA_signal_11225 ), .Q ( new_AGEMA_signal_11226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3204 ( .C ( clk ), .D ( new_AGEMA_signal_11231 ), .Q ( new_AGEMA_signal_11232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3210 ( .C ( clk ), .D ( new_AGEMA_signal_11237 ), .Q ( new_AGEMA_signal_11238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3216 ( .C ( clk ), .D ( new_AGEMA_signal_11243 ), .Q ( new_AGEMA_signal_11244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3222 ( .C ( clk ), .D ( new_AGEMA_signal_11249 ), .Q ( new_AGEMA_signal_11250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3226 ( .C ( clk ), .D ( new_AGEMA_signal_11253 ), .Q ( new_AGEMA_signal_11254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3230 ( .C ( clk ), .D ( new_AGEMA_signal_11257 ), .Q ( new_AGEMA_signal_11258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3234 ( .C ( clk ), .D ( new_AGEMA_signal_11261 ), .Q ( new_AGEMA_signal_11262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3238 ( .C ( clk ), .D ( new_AGEMA_signal_11265 ), .Q ( new_AGEMA_signal_11266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3244 ( .C ( clk ), .D ( new_AGEMA_signal_11271 ), .Q ( new_AGEMA_signal_11272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3250 ( .C ( clk ), .D ( new_AGEMA_signal_11277 ), .Q ( new_AGEMA_signal_11278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3256 ( .C ( clk ), .D ( new_AGEMA_signal_11283 ), .Q ( new_AGEMA_signal_11284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3262 ( .C ( clk ), .D ( new_AGEMA_signal_11289 ), .Q ( new_AGEMA_signal_11290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3264 ( .C ( clk ), .D ( new_AGEMA_signal_11291 ), .Q ( new_AGEMA_signal_11292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3266 ( .C ( clk ), .D ( new_AGEMA_signal_11293 ), .Q ( new_AGEMA_signal_11294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3268 ( .C ( clk ), .D ( new_AGEMA_signal_11295 ), .Q ( new_AGEMA_signal_11296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3270 ( .C ( clk ), .D ( new_AGEMA_signal_11297 ), .Q ( new_AGEMA_signal_11298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3276 ( .C ( clk ), .D ( new_AGEMA_signal_11303 ), .Q ( new_AGEMA_signal_11304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3282 ( .C ( clk ), .D ( new_AGEMA_signal_11309 ), .Q ( new_AGEMA_signal_11310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3288 ( .C ( clk ), .D ( new_AGEMA_signal_11315 ), .Q ( new_AGEMA_signal_11316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3294 ( .C ( clk ), .D ( new_AGEMA_signal_11321 ), .Q ( new_AGEMA_signal_11322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3300 ( .C ( clk ), .D ( new_AGEMA_signal_11327 ), .Q ( new_AGEMA_signal_11328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3306 ( .C ( clk ), .D ( new_AGEMA_signal_11333 ), .Q ( new_AGEMA_signal_11334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3312 ( .C ( clk ), .D ( new_AGEMA_signal_11339 ), .Q ( new_AGEMA_signal_11340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3318 ( .C ( clk ), .D ( new_AGEMA_signal_11345 ), .Q ( new_AGEMA_signal_11346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3320 ( .C ( clk ), .D ( new_AGEMA_signal_11347 ), .Q ( new_AGEMA_signal_11348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3322 ( .C ( clk ), .D ( new_AGEMA_signal_11349 ), .Q ( new_AGEMA_signal_11350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3324 ( .C ( clk ), .D ( new_AGEMA_signal_11351 ), .Q ( new_AGEMA_signal_11352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3326 ( .C ( clk ), .D ( new_AGEMA_signal_11353 ), .Q ( new_AGEMA_signal_11354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3330 ( .C ( clk ), .D ( new_AGEMA_signal_11357 ), .Q ( new_AGEMA_signal_11358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3334 ( .C ( clk ), .D ( new_AGEMA_signal_11361 ), .Q ( new_AGEMA_signal_11362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3338 ( .C ( clk ), .D ( new_AGEMA_signal_11365 ), .Q ( new_AGEMA_signal_11366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3342 ( .C ( clk ), .D ( new_AGEMA_signal_11369 ), .Q ( new_AGEMA_signal_11370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3348 ( .C ( clk ), .D ( new_AGEMA_signal_11375 ), .Q ( new_AGEMA_signal_11376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3354 ( .C ( clk ), .D ( new_AGEMA_signal_11381 ), .Q ( new_AGEMA_signal_11382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3360 ( .C ( clk ), .D ( new_AGEMA_signal_11387 ), .Q ( new_AGEMA_signal_11388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3366 ( .C ( clk ), .D ( new_AGEMA_signal_11393 ), .Q ( new_AGEMA_signal_11394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3372 ( .C ( clk ), .D ( new_AGEMA_signal_11399 ), .Q ( new_AGEMA_signal_11400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3378 ( .C ( clk ), .D ( new_AGEMA_signal_11405 ), .Q ( new_AGEMA_signal_11406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3384 ( .C ( clk ), .D ( new_AGEMA_signal_11411 ), .Q ( new_AGEMA_signal_11412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3390 ( .C ( clk ), .D ( new_AGEMA_signal_11417 ), .Q ( new_AGEMA_signal_11418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3392 ( .C ( clk ), .D ( new_AGEMA_signal_11419 ), .Q ( new_AGEMA_signal_11420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3394 ( .C ( clk ), .D ( new_AGEMA_signal_11421 ), .Q ( new_AGEMA_signal_11422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3396 ( .C ( clk ), .D ( new_AGEMA_signal_11423 ), .Q ( new_AGEMA_signal_11424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3398 ( .C ( clk ), .D ( new_AGEMA_signal_11425 ), .Q ( new_AGEMA_signal_11426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3404 ( .C ( clk ), .D ( new_AGEMA_signal_11431 ), .Q ( new_AGEMA_signal_11432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3410 ( .C ( clk ), .D ( new_AGEMA_signal_11437 ), .Q ( new_AGEMA_signal_11438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3416 ( .C ( clk ), .D ( new_AGEMA_signal_11443 ), .Q ( new_AGEMA_signal_11444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3422 ( .C ( clk ), .D ( new_AGEMA_signal_11449 ), .Q ( new_AGEMA_signal_11450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3424 ( .C ( clk ), .D ( new_AGEMA_signal_11451 ), .Q ( new_AGEMA_signal_11452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3426 ( .C ( clk ), .D ( new_AGEMA_signal_11453 ), .Q ( new_AGEMA_signal_11454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3428 ( .C ( clk ), .D ( new_AGEMA_signal_11455 ), .Q ( new_AGEMA_signal_11456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3430 ( .C ( clk ), .D ( new_AGEMA_signal_11457 ), .Q ( new_AGEMA_signal_11458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3434 ( .C ( clk ), .D ( new_AGEMA_signal_11461 ), .Q ( new_AGEMA_signal_11462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3438 ( .C ( clk ), .D ( new_AGEMA_signal_11465 ), .Q ( new_AGEMA_signal_11466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3442 ( .C ( clk ), .D ( new_AGEMA_signal_11469 ), .Q ( new_AGEMA_signal_11470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3446 ( .C ( clk ), .D ( new_AGEMA_signal_11473 ), .Q ( new_AGEMA_signal_11474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3450 ( .C ( clk ), .D ( new_AGEMA_signal_11477 ), .Q ( new_AGEMA_signal_11478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3454 ( .C ( clk ), .D ( new_AGEMA_signal_11481 ), .Q ( new_AGEMA_signal_11482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3458 ( .C ( clk ), .D ( new_AGEMA_signal_11485 ), .Q ( new_AGEMA_signal_11486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3462 ( .C ( clk ), .D ( new_AGEMA_signal_11489 ), .Q ( new_AGEMA_signal_11490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3464 ( .C ( clk ), .D ( new_AGEMA_signal_11491 ), .Q ( new_AGEMA_signal_11492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3466 ( .C ( clk ), .D ( new_AGEMA_signal_11493 ), .Q ( new_AGEMA_signal_11494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3468 ( .C ( clk ), .D ( new_AGEMA_signal_11495 ), .Q ( new_AGEMA_signal_11496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3470 ( .C ( clk ), .D ( new_AGEMA_signal_11497 ), .Q ( new_AGEMA_signal_11498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3478 ( .C ( clk ), .D ( new_AGEMA_signal_11505 ), .Q ( new_AGEMA_signal_11506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3486 ( .C ( clk ), .D ( new_AGEMA_signal_11513 ), .Q ( new_AGEMA_signal_11514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3494 ( .C ( clk ), .D ( new_AGEMA_signal_11521 ), .Q ( new_AGEMA_signal_11522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3502 ( .C ( clk ), .D ( new_AGEMA_signal_11529 ), .Q ( new_AGEMA_signal_11530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3508 ( .C ( clk ), .D ( new_AGEMA_signal_11535 ), .Q ( new_AGEMA_signal_11536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3514 ( .C ( clk ), .D ( new_AGEMA_signal_11541 ), .Q ( new_AGEMA_signal_11542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3520 ( .C ( clk ), .D ( new_AGEMA_signal_11547 ), .Q ( new_AGEMA_signal_11548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3526 ( .C ( clk ), .D ( new_AGEMA_signal_11553 ), .Q ( new_AGEMA_signal_11554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3530 ( .C ( clk ), .D ( new_AGEMA_signal_11557 ), .Q ( new_AGEMA_signal_11558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3534 ( .C ( clk ), .D ( new_AGEMA_signal_11561 ), .Q ( new_AGEMA_signal_11562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3538 ( .C ( clk ), .D ( new_AGEMA_signal_11565 ), .Q ( new_AGEMA_signal_11566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3542 ( .C ( clk ), .D ( new_AGEMA_signal_11569 ), .Q ( new_AGEMA_signal_11570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3546 ( .C ( clk ), .D ( new_AGEMA_signal_11573 ), .Q ( new_AGEMA_signal_11574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3550 ( .C ( clk ), .D ( new_AGEMA_signal_11577 ), .Q ( new_AGEMA_signal_11578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3554 ( .C ( clk ), .D ( new_AGEMA_signal_11581 ), .Q ( new_AGEMA_signal_11582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3558 ( .C ( clk ), .D ( new_AGEMA_signal_11585 ), .Q ( new_AGEMA_signal_11586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3560 ( .C ( clk ), .D ( new_AGEMA_signal_11587 ), .Q ( new_AGEMA_signal_11588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3562 ( .C ( clk ), .D ( new_AGEMA_signal_11589 ), .Q ( new_AGEMA_signal_11590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3564 ( .C ( clk ), .D ( new_AGEMA_signal_11591 ), .Q ( new_AGEMA_signal_11592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3566 ( .C ( clk ), .D ( new_AGEMA_signal_11593 ), .Q ( new_AGEMA_signal_11594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3568 ( .C ( clk ), .D ( new_AGEMA_signal_11595 ), .Q ( new_AGEMA_signal_11596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3570 ( .C ( clk ), .D ( new_AGEMA_signal_11597 ), .Q ( new_AGEMA_signal_11598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3572 ( .C ( clk ), .D ( new_AGEMA_signal_11599 ), .Q ( new_AGEMA_signal_11600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3574 ( .C ( clk ), .D ( new_AGEMA_signal_11601 ), .Q ( new_AGEMA_signal_11602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3578 ( .C ( clk ), .D ( new_AGEMA_signal_11605 ), .Q ( new_AGEMA_signal_11606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3582 ( .C ( clk ), .D ( new_AGEMA_signal_11609 ), .Q ( new_AGEMA_signal_11610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3586 ( .C ( clk ), .D ( new_AGEMA_signal_11613 ), .Q ( new_AGEMA_signal_11614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3590 ( .C ( clk ), .D ( new_AGEMA_signal_11617 ), .Q ( new_AGEMA_signal_11618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3594 ( .C ( clk ), .D ( new_AGEMA_signal_11621 ), .Q ( new_AGEMA_signal_11622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3598 ( .C ( clk ), .D ( new_AGEMA_signal_11625 ), .Q ( new_AGEMA_signal_11626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3602 ( .C ( clk ), .D ( new_AGEMA_signal_11629 ), .Q ( new_AGEMA_signal_11630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3606 ( .C ( clk ), .D ( new_AGEMA_signal_11633 ), .Q ( new_AGEMA_signal_11634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3608 ( .C ( clk ), .D ( new_AGEMA_signal_11635 ), .Q ( new_AGEMA_signal_11636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3610 ( .C ( clk ), .D ( new_AGEMA_signal_11637 ), .Q ( new_AGEMA_signal_11638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3612 ( .C ( clk ), .D ( new_AGEMA_signal_11639 ), .Q ( new_AGEMA_signal_11640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3614 ( .C ( clk ), .D ( new_AGEMA_signal_11641 ), .Q ( new_AGEMA_signal_11642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3620 ( .C ( clk ), .D ( new_AGEMA_signal_11647 ), .Q ( new_AGEMA_signal_11648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3626 ( .C ( clk ), .D ( new_AGEMA_signal_11653 ), .Q ( new_AGEMA_signal_11654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3632 ( .C ( clk ), .D ( new_AGEMA_signal_11659 ), .Q ( new_AGEMA_signal_11660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3638 ( .C ( clk ), .D ( new_AGEMA_signal_11665 ), .Q ( new_AGEMA_signal_11666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3642 ( .C ( clk ), .D ( new_AGEMA_signal_11669 ), .Q ( new_AGEMA_signal_11670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3646 ( .C ( clk ), .D ( new_AGEMA_signal_11673 ), .Q ( new_AGEMA_signal_11674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3650 ( .C ( clk ), .D ( new_AGEMA_signal_11677 ), .Q ( new_AGEMA_signal_11678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3654 ( .C ( clk ), .D ( new_AGEMA_signal_11681 ), .Q ( new_AGEMA_signal_11682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3656 ( .C ( clk ), .D ( new_AGEMA_signal_11683 ), .Q ( new_AGEMA_signal_11684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3658 ( .C ( clk ), .D ( new_AGEMA_signal_11685 ), .Q ( new_AGEMA_signal_11686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3660 ( .C ( clk ), .D ( new_AGEMA_signal_11687 ), .Q ( new_AGEMA_signal_11688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3662 ( .C ( clk ), .D ( new_AGEMA_signal_11689 ), .Q ( new_AGEMA_signal_11690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3666 ( .C ( clk ), .D ( new_AGEMA_signal_11693 ), .Q ( new_AGEMA_signal_11694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3670 ( .C ( clk ), .D ( new_AGEMA_signal_11697 ), .Q ( new_AGEMA_signal_11698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3674 ( .C ( clk ), .D ( new_AGEMA_signal_11701 ), .Q ( new_AGEMA_signal_11702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3678 ( .C ( clk ), .D ( new_AGEMA_signal_11705 ), .Q ( new_AGEMA_signal_11706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3682 ( .C ( clk ), .D ( new_AGEMA_signal_11709 ), .Q ( new_AGEMA_signal_11710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3686 ( .C ( clk ), .D ( new_AGEMA_signal_11713 ), .Q ( new_AGEMA_signal_11714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3690 ( .C ( clk ), .D ( new_AGEMA_signal_11717 ), .Q ( new_AGEMA_signal_11718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3694 ( .C ( clk ), .D ( new_AGEMA_signal_11721 ), .Q ( new_AGEMA_signal_11722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3698 ( .C ( clk ), .D ( new_AGEMA_signal_11725 ), .Q ( new_AGEMA_signal_11726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3702 ( .C ( clk ), .D ( new_AGEMA_signal_11729 ), .Q ( new_AGEMA_signal_11730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3706 ( .C ( clk ), .D ( new_AGEMA_signal_11733 ), .Q ( new_AGEMA_signal_11734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3710 ( .C ( clk ), .D ( new_AGEMA_signal_11737 ), .Q ( new_AGEMA_signal_11738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3712 ( .C ( clk ), .D ( new_AGEMA_signal_11739 ), .Q ( new_AGEMA_signal_11740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3714 ( .C ( clk ), .D ( new_AGEMA_signal_11741 ), .Q ( new_AGEMA_signal_11742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3716 ( .C ( clk ), .D ( new_AGEMA_signal_11743 ), .Q ( new_AGEMA_signal_11744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3718 ( .C ( clk ), .D ( new_AGEMA_signal_11745 ), .Q ( new_AGEMA_signal_11746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3722 ( .C ( clk ), .D ( new_AGEMA_signal_11749 ), .Q ( new_AGEMA_signal_11750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3726 ( .C ( clk ), .D ( new_AGEMA_signal_11753 ), .Q ( new_AGEMA_signal_11754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3730 ( .C ( clk ), .D ( new_AGEMA_signal_11757 ), .Q ( new_AGEMA_signal_11758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3734 ( .C ( clk ), .D ( new_AGEMA_signal_11761 ), .Q ( new_AGEMA_signal_11762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3736 ( .C ( clk ), .D ( new_AGEMA_signal_11763 ), .Q ( new_AGEMA_signal_11764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3738 ( .C ( clk ), .D ( new_AGEMA_signal_11765 ), .Q ( new_AGEMA_signal_11766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3740 ( .C ( clk ), .D ( new_AGEMA_signal_11767 ), .Q ( new_AGEMA_signal_11768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3742 ( .C ( clk ), .D ( new_AGEMA_signal_11769 ), .Q ( new_AGEMA_signal_11770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3748 ( .C ( clk ), .D ( new_AGEMA_signal_11775 ), .Q ( new_AGEMA_signal_11776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3754 ( .C ( clk ), .D ( new_AGEMA_signal_11781 ), .Q ( new_AGEMA_signal_11782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3760 ( .C ( clk ), .D ( new_AGEMA_signal_11787 ), .Q ( new_AGEMA_signal_11788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3766 ( .C ( clk ), .D ( new_AGEMA_signal_11793 ), .Q ( new_AGEMA_signal_11794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3772 ( .C ( clk ), .D ( new_AGEMA_signal_11799 ), .Q ( new_AGEMA_signal_11800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3778 ( .C ( clk ), .D ( new_AGEMA_signal_11805 ), .Q ( new_AGEMA_signal_11806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3784 ( .C ( clk ), .D ( new_AGEMA_signal_11811 ), .Q ( new_AGEMA_signal_11812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3790 ( .C ( clk ), .D ( new_AGEMA_signal_11817 ), .Q ( new_AGEMA_signal_11818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3794 ( .C ( clk ), .D ( new_AGEMA_signal_11821 ), .Q ( new_AGEMA_signal_11822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3798 ( .C ( clk ), .D ( new_AGEMA_signal_11825 ), .Q ( new_AGEMA_signal_11826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3802 ( .C ( clk ), .D ( new_AGEMA_signal_11829 ), .Q ( new_AGEMA_signal_11830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3806 ( .C ( clk ), .D ( new_AGEMA_signal_11833 ), .Q ( new_AGEMA_signal_11834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3808 ( .C ( clk ), .D ( new_AGEMA_signal_11835 ), .Q ( new_AGEMA_signal_11836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3810 ( .C ( clk ), .D ( new_AGEMA_signal_11837 ), .Q ( new_AGEMA_signal_11838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3812 ( .C ( clk ), .D ( new_AGEMA_signal_11839 ), .Q ( new_AGEMA_signal_11840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3814 ( .C ( clk ), .D ( new_AGEMA_signal_11841 ), .Q ( new_AGEMA_signal_11842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3822 ( .C ( clk ), .D ( new_AGEMA_signal_11849 ), .Q ( new_AGEMA_signal_11850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3830 ( .C ( clk ), .D ( new_AGEMA_signal_11857 ), .Q ( new_AGEMA_signal_11858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3838 ( .C ( clk ), .D ( new_AGEMA_signal_11865 ), .Q ( new_AGEMA_signal_11866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3846 ( .C ( clk ), .D ( new_AGEMA_signal_11873 ), .Q ( new_AGEMA_signal_11874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3848 ( .C ( clk ), .D ( new_AGEMA_signal_11875 ), .Q ( new_AGEMA_signal_11876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3850 ( .C ( clk ), .D ( new_AGEMA_signal_11877 ), .Q ( new_AGEMA_signal_11878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3852 ( .C ( clk ), .D ( new_AGEMA_signal_11879 ), .Q ( new_AGEMA_signal_11880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3854 ( .C ( clk ), .D ( new_AGEMA_signal_11881 ), .Q ( new_AGEMA_signal_11882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3858 ( .C ( clk ), .D ( new_AGEMA_signal_11885 ), .Q ( new_AGEMA_signal_11886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3862 ( .C ( clk ), .D ( new_AGEMA_signal_11889 ), .Q ( new_AGEMA_signal_11890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3866 ( .C ( clk ), .D ( new_AGEMA_signal_11893 ), .Q ( new_AGEMA_signal_11894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3870 ( .C ( clk ), .D ( new_AGEMA_signal_11897 ), .Q ( new_AGEMA_signal_11898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3874 ( .C ( clk ), .D ( new_AGEMA_signal_11901 ), .Q ( new_AGEMA_signal_11902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3878 ( .C ( clk ), .D ( new_AGEMA_signal_11905 ), .Q ( new_AGEMA_signal_11906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3882 ( .C ( clk ), .D ( new_AGEMA_signal_11909 ), .Q ( new_AGEMA_signal_11910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3886 ( .C ( clk ), .D ( new_AGEMA_signal_11913 ), .Q ( new_AGEMA_signal_11914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3890 ( .C ( clk ), .D ( new_AGEMA_signal_11917 ), .Q ( new_AGEMA_signal_11918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3894 ( .C ( clk ), .D ( new_AGEMA_signal_11921 ), .Q ( new_AGEMA_signal_11922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3898 ( .C ( clk ), .D ( new_AGEMA_signal_11925 ), .Q ( new_AGEMA_signal_11926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3902 ( .C ( clk ), .D ( new_AGEMA_signal_11929 ), .Q ( new_AGEMA_signal_11930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3906 ( .C ( clk ), .D ( new_AGEMA_signal_11933 ), .Q ( new_AGEMA_signal_11934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3910 ( .C ( clk ), .D ( new_AGEMA_signal_11937 ), .Q ( new_AGEMA_signal_11938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3914 ( .C ( clk ), .D ( new_AGEMA_signal_11941 ), .Q ( new_AGEMA_signal_11942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3918 ( .C ( clk ), .D ( new_AGEMA_signal_11945 ), .Q ( new_AGEMA_signal_11946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3922 ( .C ( clk ), .D ( new_AGEMA_signal_11949 ), .Q ( new_AGEMA_signal_11950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3926 ( .C ( clk ), .D ( new_AGEMA_signal_11953 ), .Q ( new_AGEMA_signal_11954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3930 ( .C ( clk ), .D ( new_AGEMA_signal_11957 ), .Q ( new_AGEMA_signal_11958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3934 ( .C ( clk ), .D ( new_AGEMA_signal_11961 ), .Q ( new_AGEMA_signal_11962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3942 ( .C ( clk ), .D ( new_AGEMA_signal_11969 ), .Q ( new_AGEMA_signal_11970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3950 ( .C ( clk ), .D ( new_AGEMA_signal_11977 ), .Q ( new_AGEMA_signal_11978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3958 ( .C ( clk ), .D ( new_AGEMA_signal_11985 ), .Q ( new_AGEMA_signal_11986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3966 ( .C ( clk ), .D ( new_AGEMA_signal_11993 ), .Q ( new_AGEMA_signal_11994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3968 ( .C ( clk ), .D ( new_AGEMA_signal_11995 ), .Q ( new_AGEMA_signal_11996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3970 ( .C ( clk ), .D ( new_AGEMA_signal_11997 ), .Q ( new_AGEMA_signal_11998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3972 ( .C ( clk ), .D ( new_AGEMA_signal_11999 ), .Q ( new_AGEMA_signal_12000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3974 ( .C ( clk ), .D ( new_AGEMA_signal_12001 ), .Q ( new_AGEMA_signal_12002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3978 ( .C ( clk ), .D ( new_AGEMA_signal_12005 ), .Q ( new_AGEMA_signal_12006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3982 ( .C ( clk ), .D ( new_AGEMA_signal_12009 ), .Q ( new_AGEMA_signal_12010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3986 ( .C ( clk ), .D ( new_AGEMA_signal_12013 ), .Q ( new_AGEMA_signal_12014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3990 ( .C ( clk ), .D ( new_AGEMA_signal_12017 ), .Q ( new_AGEMA_signal_12018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3992 ( .C ( clk ), .D ( new_AGEMA_signal_12019 ), .Q ( new_AGEMA_signal_12020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3994 ( .C ( clk ), .D ( new_AGEMA_signal_12021 ), .Q ( new_AGEMA_signal_12022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3996 ( .C ( clk ), .D ( new_AGEMA_signal_12023 ), .Q ( new_AGEMA_signal_12024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_3998 ( .C ( clk ), .D ( new_AGEMA_signal_12025 ), .Q ( new_AGEMA_signal_12026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4004 ( .C ( clk ), .D ( new_AGEMA_signal_12031 ), .Q ( new_AGEMA_signal_12032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4010 ( .C ( clk ), .D ( new_AGEMA_signal_12037 ), .Q ( new_AGEMA_signal_12038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4016 ( .C ( clk ), .D ( new_AGEMA_signal_12043 ), .Q ( new_AGEMA_signal_12044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4022 ( .C ( clk ), .D ( new_AGEMA_signal_12049 ), .Q ( new_AGEMA_signal_12050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4036 ( .C ( clk ), .D ( new_AGEMA_signal_12063 ), .Q ( new_AGEMA_signal_12064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4044 ( .C ( clk ), .D ( new_AGEMA_signal_12071 ), .Q ( new_AGEMA_signal_12072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4052 ( .C ( clk ), .D ( new_AGEMA_signal_12079 ), .Q ( new_AGEMA_signal_12080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4060 ( .C ( clk ), .D ( new_AGEMA_signal_12087 ), .Q ( new_AGEMA_signal_12088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4072 ( .C ( clk ), .D ( new_AGEMA_signal_12099 ), .Q ( new_AGEMA_signal_12100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4076 ( .C ( clk ), .D ( new_AGEMA_signal_12103 ), .Q ( new_AGEMA_signal_12104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4080 ( .C ( clk ), .D ( new_AGEMA_signal_12107 ), .Q ( new_AGEMA_signal_12108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4084 ( .C ( clk ), .D ( new_AGEMA_signal_12111 ), .Q ( new_AGEMA_signal_12112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4092 ( .C ( clk ), .D ( new_AGEMA_signal_12119 ), .Q ( new_AGEMA_signal_12120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4100 ( .C ( clk ), .D ( new_AGEMA_signal_12127 ), .Q ( new_AGEMA_signal_12128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4108 ( .C ( clk ), .D ( new_AGEMA_signal_12135 ), .Q ( new_AGEMA_signal_12136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4116 ( .C ( clk ), .D ( new_AGEMA_signal_12143 ), .Q ( new_AGEMA_signal_12144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4130 ( .C ( clk ), .D ( new_AGEMA_signal_12157 ), .Q ( new_AGEMA_signal_12158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4136 ( .C ( clk ), .D ( new_AGEMA_signal_12163 ), .Q ( new_AGEMA_signal_12164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4142 ( .C ( clk ), .D ( new_AGEMA_signal_12169 ), .Q ( new_AGEMA_signal_12170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4148 ( .C ( clk ), .D ( new_AGEMA_signal_12175 ), .Q ( new_AGEMA_signal_12176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4152 ( .C ( clk ), .D ( new_AGEMA_signal_12179 ), .Q ( new_AGEMA_signal_12180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4156 ( .C ( clk ), .D ( new_AGEMA_signal_12183 ), .Q ( new_AGEMA_signal_12184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4160 ( .C ( clk ), .D ( new_AGEMA_signal_12187 ), .Q ( new_AGEMA_signal_12188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4164 ( .C ( clk ), .D ( new_AGEMA_signal_12191 ), .Q ( new_AGEMA_signal_12192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4172 ( .C ( clk ), .D ( new_AGEMA_signal_12199 ), .Q ( new_AGEMA_signal_12200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4180 ( .C ( clk ), .D ( new_AGEMA_signal_12207 ), .Q ( new_AGEMA_signal_12208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4188 ( .C ( clk ), .D ( new_AGEMA_signal_12215 ), .Q ( new_AGEMA_signal_12216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4196 ( .C ( clk ), .D ( new_AGEMA_signal_12223 ), .Q ( new_AGEMA_signal_12224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4200 ( .C ( clk ), .D ( new_AGEMA_signal_12227 ), .Q ( new_AGEMA_signal_12228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4204 ( .C ( clk ), .D ( new_AGEMA_signal_12231 ), .Q ( new_AGEMA_signal_12232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4208 ( .C ( clk ), .D ( new_AGEMA_signal_12235 ), .Q ( new_AGEMA_signal_12236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4212 ( .C ( clk ), .D ( new_AGEMA_signal_12239 ), .Q ( new_AGEMA_signal_12240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4218 ( .C ( clk ), .D ( new_AGEMA_signal_12245 ), .Q ( new_AGEMA_signal_12246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4224 ( .C ( clk ), .D ( new_AGEMA_signal_12251 ), .Q ( new_AGEMA_signal_12252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4230 ( .C ( clk ), .D ( new_AGEMA_signal_12257 ), .Q ( new_AGEMA_signal_12258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4236 ( .C ( clk ), .D ( new_AGEMA_signal_12263 ), .Q ( new_AGEMA_signal_12264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4242 ( .C ( clk ), .D ( new_AGEMA_signal_12269 ), .Q ( new_AGEMA_signal_12270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4248 ( .C ( clk ), .D ( new_AGEMA_signal_12275 ), .Q ( new_AGEMA_signal_12276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4254 ( .C ( clk ), .D ( new_AGEMA_signal_12281 ), .Q ( new_AGEMA_signal_12282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4260 ( .C ( clk ), .D ( new_AGEMA_signal_12287 ), .Q ( new_AGEMA_signal_12288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4266 ( .C ( clk ), .D ( new_AGEMA_signal_12293 ), .Q ( new_AGEMA_signal_12294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4272 ( .C ( clk ), .D ( new_AGEMA_signal_12299 ), .Q ( new_AGEMA_signal_12300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4278 ( .C ( clk ), .D ( new_AGEMA_signal_12305 ), .Q ( new_AGEMA_signal_12306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4284 ( .C ( clk ), .D ( new_AGEMA_signal_12311 ), .Q ( new_AGEMA_signal_12312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4290 ( .C ( clk ), .D ( new_AGEMA_signal_12317 ), .Q ( new_AGEMA_signal_12318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4296 ( .C ( clk ), .D ( new_AGEMA_signal_12323 ), .Q ( new_AGEMA_signal_12324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4302 ( .C ( clk ), .D ( new_AGEMA_signal_12329 ), .Q ( new_AGEMA_signal_12330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4308 ( .C ( clk ), .D ( new_AGEMA_signal_12335 ), .Q ( new_AGEMA_signal_12336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4314 ( .C ( clk ), .D ( new_AGEMA_signal_12341 ), .Q ( new_AGEMA_signal_12342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4320 ( .C ( clk ), .D ( new_AGEMA_signal_12347 ), .Q ( new_AGEMA_signal_12348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4326 ( .C ( clk ), .D ( new_AGEMA_signal_12353 ), .Q ( new_AGEMA_signal_12354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4332 ( .C ( clk ), .D ( new_AGEMA_signal_12359 ), .Q ( new_AGEMA_signal_12360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4336 ( .C ( clk ), .D ( new_AGEMA_signal_12363 ), .Q ( new_AGEMA_signal_12364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4340 ( .C ( clk ), .D ( new_AGEMA_signal_12367 ), .Q ( new_AGEMA_signal_12368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4344 ( .C ( clk ), .D ( new_AGEMA_signal_12371 ), .Q ( new_AGEMA_signal_12372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4348 ( .C ( clk ), .D ( new_AGEMA_signal_12375 ), .Q ( new_AGEMA_signal_12376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4356 ( .C ( clk ), .D ( new_AGEMA_signal_12383 ), .Q ( new_AGEMA_signal_12384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4364 ( .C ( clk ), .D ( new_AGEMA_signal_12391 ), .Q ( new_AGEMA_signal_12392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4372 ( .C ( clk ), .D ( new_AGEMA_signal_12399 ), .Q ( new_AGEMA_signal_12400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4380 ( .C ( clk ), .D ( new_AGEMA_signal_12407 ), .Q ( new_AGEMA_signal_12408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4384 ( .C ( clk ), .D ( new_AGEMA_signal_12411 ), .Q ( new_AGEMA_signal_12412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4388 ( .C ( clk ), .D ( new_AGEMA_signal_12415 ), .Q ( new_AGEMA_signal_12416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4392 ( .C ( clk ), .D ( new_AGEMA_signal_12419 ), .Q ( new_AGEMA_signal_12420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4396 ( .C ( clk ), .D ( new_AGEMA_signal_12423 ), .Q ( new_AGEMA_signal_12424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4402 ( .C ( clk ), .D ( new_AGEMA_signal_12429 ), .Q ( new_AGEMA_signal_12430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4408 ( .C ( clk ), .D ( new_AGEMA_signal_12435 ), .Q ( new_AGEMA_signal_12436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4414 ( .C ( clk ), .D ( new_AGEMA_signal_12441 ), .Q ( new_AGEMA_signal_12442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4420 ( .C ( clk ), .D ( new_AGEMA_signal_12447 ), .Q ( new_AGEMA_signal_12448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4428 ( .C ( clk ), .D ( new_AGEMA_signal_12455 ), .Q ( new_AGEMA_signal_12456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4436 ( .C ( clk ), .D ( new_AGEMA_signal_12463 ), .Q ( new_AGEMA_signal_12464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4444 ( .C ( clk ), .D ( new_AGEMA_signal_12471 ), .Q ( new_AGEMA_signal_12472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4452 ( .C ( clk ), .D ( new_AGEMA_signal_12479 ), .Q ( new_AGEMA_signal_12480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4466 ( .C ( clk ), .D ( new_AGEMA_signal_12493 ), .Q ( new_AGEMA_signal_12494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4472 ( .C ( clk ), .D ( new_AGEMA_signal_12499 ), .Q ( new_AGEMA_signal_12500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4478 ( .C ( clk ), .D ( new_AGEMA_signal_12505 ), .Q ( new_AGEMA_signal_12506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4484 ( .C ( clk ), .D ( new_AGEMA_signal_12511 ), .Q ( new_AGEMA_signal_12512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4506 ( .C ( clk ), .D ( new_AGEMA_signal_12533 ), .Q ( new_AGEMA_signal_12534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4512 ( .C ( clk ), .D ( new_AGEMA_signal_12539 ), .Q ( new_AGEMA_signal_12540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4518 ( .C ( clk ), .D ( new_AGEMA_signal_12545 ), .Q ( new_AGEMA_signal_12546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4524 ( .C ( clk ), .D ( new_AGEMA_signal_12551 ), .Q ( new_AGEMA_signal_12552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4530 ( .C ( clk ), .D ( new_AGEMA_signal_12557 ), .Q ( new_AGEMA_signal_12558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4536 ( .C ( clk ), .D ( new_AGEMA_signal_12563 ), .Q ( new_AGEMA_signal_12564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4542 ( .C ( clk ), .D ( new_AGEMA_signal_12569 ), .Q ( new_AGEMA_signal_12570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4548 ( .C ( clk ), .D ( new_AGEMA_signal_12575 ), .Q ( new_AGEMA_signal_12576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4556 ( .C ( clk ), .D ( new_AGEMA_signal_12583 ), .Q ( new_AGEMA_signal_12584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4564 ( .C ( clk ), .D ( new_AGEMA_signal_12591 ), .Q ( new_AGEMA_signal_12592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4572 ( .C ( clk ), .D ( new_AGEMA_signal_12599 ), .Q ( new_AGEMA_signal_12600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4580 ( .C ( clk ), .D ( new_AGEMA_signal_12607 ), .Q ( new_AGEMA_signal_12608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4588 ( .C ( clk ), .D ( new_AGEMA_signal_12615 ), .Q ( new_AGEMA_signal_12616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4596 ( .C ( clk ), .D ( new_AGEMA_signal_12623 ), .Q ( new_AGEMA_signal_12624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4604 ( .C ( clk ), .D ( new_AGEMA_signal_12631 ), .Q ( new_AGEMA_signal_12632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4612 ( .C ( clk ), .D ( new_AGEMA_signal_12639 ), .Q ( new_AGEMA_signal_12640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4618 ( .C ( clk ), .D ( new_AGEMA_signal_12645 ), .Q ( new_AGEMA_signal_12646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4624 ( .C ( clk ), .D ( new_AGEMA_signal_12651 ), .Q ( new_AGEMA_signal_12652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4630 ( .C ( clk ), .D ( new_AGEMA_signal_12657 ), .Q ( new_AGEMA_signal_12658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4636 ( .C ( clk ), .D ( new_AGEMA_signal_12663 ), .Q ( new_AGEMA_signal_12664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4642 ( .C ( clk ), .D ( new_AGEMA_signal_12669 ), .Q ( new_AGEMA_signal_12670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4648 ( .C ( clk ), .D ( new_AGEMA_signal_12675 ), .Q ( new_AGEMA_signal_12676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4654 ( .C ( clk ), .D ( new_AGEMA_signal_12681 ), .Q ( new_AGEMA_signal_12682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4660 ( .C ( clk ), .D ( new_AGEMA_signal_12687 ), .Q ( new_AGEMA_signal_12688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4672 ( .C ( clk ), .D ( new_AGEMA_signal_12699 ), .Q ( new_AGEMA_signal_12700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4676 ( .C ( clk ), .D ( new_AGEMA_signal_12703 ), .Q ( new_AGEMA_signal_12704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4680 ( .C ( clk ), .D ( new_AGEMA_signal_12707 ), .Q ( new_AGEMA_signal_12708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4684 ( .C ( clk ), .D ( new_AGEMA_signal_12711 ), .Q ( new_AGEMA_signal_12712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4688 ( .C ( clk ), .D ( new_AGEMA_signal_12715 ), .Q ( new_AGEMA_signal_12716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4692 ( .C ( clk ), .D ( new_AGEMA_signal_12719 ), .Q ( new_AGEMA_signal_12720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4696 ( .C ( clk ), .D ( new_AGEMA_signal_12723 ), .Q ( new_AGEMA_signal_12724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4700 ( .C ( clk ), .D ( new_AGEMA_signal_12727 ), .Q ( new_AGEMA_signal_12728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4704 ( .C ( clk ), .D ( new_AGEMA_signal_12731 ), .Q ( new_AGEMA_signal_12732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4708 ( .C ( clk ), .D ( new_AGEMA_signal_12735 ), .Q ( new_AGEMA_signal_12736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4712 ( .C ( clk ), .D ( new_AGEMA_signal_12739 ), .Q ( new_AGEMA_signal_12740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4716 ( .C ( clk ), .D ( new_AGEMA_signal_12743 ), .Q ( new_AGEMA_signal_12744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4728 ( .C ( clk ), .D ( new_AGEMA_signal_12755 ), .Q ( new_AGEMA_signal_12756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4734 ( .C ( clk ), .D ( new_AGEMA_signal_12761 ), .Q ( new_AGEMA_signal_12762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4740 ( .C ( clk ), .D ( new_AGEMA_signal_12767 ), .Q ( new_AGEMA_signal_12768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4746 ( .C ( clk ), .D ( new_AGEMA_signal_12773 ), .Q ( new_AGEMA_signal_12774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4778 ( .C ( clk ), .D ( new_AGEMA_signal_12805 ), .Q ( new_AGEMA_signal_12806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4786 ( .C ( clk ), .D ( new_AGEMA_signal_12813 ), .Q ( new_AGEMA_signal_12814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4794 ( .C ( clk ), .D ( new_AGEMA_signal_12821 ), .Q ( new_AGEMA_signal_12822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4802 ( .C ( clk ), .D ( new_AGEMA_signal_12829 ), .Q ( new_AGEMA_signal_12830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4810 ( .C ( clk ), .D ( new_AGEMA_signal_12837 ), .Q ( new_AGEMA_signal_12838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4818 ( .C ( clk ), .D ( new_AGEMA_signal_12845 ), .Q ( new_AGEMA_signal_12846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4826 ( .C ( clk ), .D ( new_AGEMA_signal_12853 ), .Q ( new_AGEMA_signal_12854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4834 ( .C ( clk ), .D ( new_AGEMA_signal_12861 ), .Q ( new_AGEMA_signal_12862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4842 ( .C ( clk ), .D ( new_AGEMA_signal_12869 ), .Q ( new_AGEMA_signal_12870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4850 ( .C ( clk ), .D ( new_AGEMA_signal_12877 ), .Q ( new_AGEMA_signal_12878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4858 ( .C ( clk ), .D ( new_AGEMA_signal_12885 ), .Q ( new_AGEMA_signal_12886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4866 ( .C ( clk ), .D ( new_AGEMA_signal_12893 ), .Q ( new_AGEMA_signal_12894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4874 ( .C ( clk ), .D ( new_AGEMA_signal_12901 ), .Q ( new_AGEMA_signal_12902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4882 ( .C ( clk ), .D ( new_AGEMA_signal_12909 ), .Q ( new_AGEMA_signal_12910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4890 ( .C ( clk ), .D ( new_AGEMA_signal_12917 ), .Q ( new_AGEMA_signal_12918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4898 ( .C ( clk ), .D ( new_AGEMA_signal_12925 ), .Q ( new_AGEMA_signal_12926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4904 ( .C ( clk ), .D ( new_AGEMA_signal_12931 ), .Q ( new_AGEMA_signal_12932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4910 ( .C ( clk ), .D ( new_AGEMA_signal_12937 ), .Q ( new_AGEMA_signal_12938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4916 ( .C ( clk ), .D ( new_AGEMA_signal_12943 ), .Q ( new_AGEMA_signal_12944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4922 ( .C ( clk ), .D ( new_AGEMA_signal_12949 ), .Q ( new_AGEMA_signal_12950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4932 ( .C ( clk ), .D ( new_AGEMA_signal_12959 ), .Q ( new_AGEMA_signal_12960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4942 ( .C ( clk ), .D ( new_AGEMA_signal_12969 ), .Q ( new_AGEMA_signal_12970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4952 ( .C ( clk ), .D ( new_AGEMA_signal_12979 ), .Q ( new_AGEMA_signal_12980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4962 ( .C ( clk ), .D ( new_AGEMA_signal_12989 ), .Q ( new_AGEMA_signal_12990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4970 ( .C ( clk ), .D ( new_AGEMA_signal_12997 ), .Q ( new_AGEMA_signal_12998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4978 ( .C ( clk ), .D ( new_AGEMA_signal_13005 ), .Q ( new_AGEMA_signal_13006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4986 ( .C ( clk ), .D ( new_AGEMA_signal_13013 ), .Q ( new_AGEMA_signal_13014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4994 ( .C ( clk ), .D ( new_AGEMA_signal_13021 ), .Q ( new_AGEMA_signal_13022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5002 ( .C ( clk ), .D ( new_AGEMA_signal_13029 ), .Q ( new_AGEMA_signal_13030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5010 ( .C ( clk ), .D ( new_AGEMA_signal_13037 ), .Q ( new_AGEMA_signal_13038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5018 ( .C ( clk ), .D ( new_AGEMA_signal_13045 ), .Q ( new_AGEMA_signal_13046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5026 ( .C ( clk ), .D ( new_AGEMA_signal_13053 ), .Q ( new_AGEMA_signal_13054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5034 ( .C ( clk ), .D ( new_AGEMA_signal_13061 ), .Q ( new_AGEMA_signal_13062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5042 ( .C ( clk ), .D ( new_AGEMA_signal_13069 ), .Q ( new_AGEMA_signal_13070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5050 ( .C ( clk ), .D ( new_AGEMA_signal_13077 ), .Q ( new_AGEMA_signal_13078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5058 ( .C ( clk ), .D ( new_AGEMA_signal_13085 ), .Q ( new_AGEMA_signal_13086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5088 ( .C ( clk ), .D ( new_AGEMA_signal_13115 ), .Q ( new_AGEMA_signal_13116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5094 ( .C ( clk ), .D ( new_AGEMA_signal_13121 ), .Q ( new_AGEMA_signal_13122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5100 ( .C ( clk ), .D ( new_AGEMA_signal_13127 ), .Q ( new_AGEMA_signal_13128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5106 ( .C ( clk ), .D ( new_AGEMA_signal_13133 ), .Q ( new_AGEMA_signal_13134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5132 ( .C ( clk ), .D ( new_AGEMA_signal_13159 ), .Q ( new_AGEMA_signal_13160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5142 ( .C ( clk ), .D ( new_AGEMA_signal_13169 ), .Q ( new_AGEMA_signal_13170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5152 ( .C ( clk ), .D ( new_AGEMA_signal_13179 ), .Q ( new_AGEMA_signal_13180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5162 ( .C ( clk ), .D ( new_AGEMA_signal_13189 ), .Q ( new_AGEMA_signal_13190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5170 ( .C ( clk ), .D ( new_AGEMA_signal_13197 ), .Q ( new_AGEMA_signal_13198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5178 ( .C ( clk ), .D ( new_AGEMA_signal_13205 ), .Q ( new_AGEMA_signal_13206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5186 ( .C ( clk ), .D ( new_AGEMA_signal_13213 ), .Q ( new_AGEMA_signal_13214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C ( clk ), .D ( new_AGEMA_signal_13221 ), .Q ( new_AGEMA_signal_13222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C ( clk ), .D ( new_AGEMA_signal_13253 ), .Q ( new_AGEMA_signal_13254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C ( clk ), .D ( new_AGEMA_signal_13261 ), .Q ( new_AGEMA_signal_13262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C ( clk ), .D ( new_AGEMA_signal_13269 ), .Q ( new_AGEMA_signal_13270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C ( clk ), .D ( new_AGEMA_signal_13277 ), .Q ( new_AGEMA_signal_13278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5258 ( .C ( clk ), .D ( new_AGEMA_signal_13285 ), .Q ( new_AGEMA_signal_13286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5266 ( .C ( clk ), .D ( new_AGEMA_signal_13293 ), .Q ( new_AGEMA_signal_13294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5274 ( .C ( clk ), .D ( new_AGEMA_signal_13301 ), .Q ( new_AGEMA_signal_13302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5282 ( .C ( clk ), .D ( new_AGEMA_signal_13309 ), .Q ( new_AGEMA_signal_13310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5288 ( .C ( clk ), .D ( new_AGEMA_signal_13315 ), .Q ( new_AGEMA_signal_13316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5294 ( .C ( clk ), .D ( new_AGEMA_signal_13321 ), .Q ( new_AGEMA_signal_13322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5300 ( .C ( clk ), .D ( new_AGEMA_signal_13327 ), .Q ( new_AGEMA_signal_13328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5306 ( .C ( clk ), .D ( new_AGEMA_signal_13333 ), .Q ( new_AGEMA_signal_13334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5330 ( .C ( clk ), .D ( new_AGEMA_signal_13357 ), .Q ( new_AGEMA_signal_13358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5338 ( .C ( clk ), .D ( new_AGEMA_signal_13365 ), .Q ( new_AGEMA_signal_13366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5346 ( .C ( clk ), .D ( new_AGEMA_signal_13373 ), .Q ( new_AGEMA_signal_13374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5354 ( .C ( clk ), .D ( new_AGEMA_signal_13381 ), .Q ( new_AGEMA_signal_13382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5456 ( .C ( clk ), .D ( new_AGEMA_signal_13483 ), .Q ( new_AGEMA_signal_13484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5464 ( .C ( clk ), .D ( new_AGEMA_signal_13491 ), .Q ( new_AGEMA_signal_13492 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5472 ( .C ( clk ), .D ( new_AGEMA_signal_13499 ), .Q ( new_AGEMA_signal_13500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5480 ( .C ( clk ), .D ( new_AGEMA_signal_13507 ), .Q ( new_AGEMA_signal_13508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5528 ( .C ( clk ), .D ( new_AGEMA_signal_13555 ), .Q ( new_AGEMA_signal_13556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5536 ( .C ( clk ), .D ( new_AGEMA_signal_13563 ), .Q ( new_AGEMA_signal_13564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5544 ( .C ( clk ), .D ( new_AGEMA_signal_13571 ), .Q ( new_AGEMA_signal_13572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5552 ( .C ( clk ), .D ( new_AGEMA_signal_13579 ), .Q ( new_AGEMA_signal_13580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5560 ( .C ( clk ), .D ( new_AGEMA_signal_13587 ), .Q ( new_AGEMA_signal_13588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5568 ( .C ( clk ), .D ( new_AGEMA_signal_13595 ), .Q ( new_AGEMA_signal_13596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5576 ( .C ( clk ), .D ( new_AGEMA_signal_13603 ), .Q ( new_AGEMA_signal_13604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5584 ( .C ( clk ), .D ( new_AGEMA_signal_13611 ), .Q ( new_AGEMA_signal_13612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5594 ( .C ( clk ), .D ( new_AGEMA_signal_13621 ), .Q ( new_AGEMA_signal_13622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5604 ( .C ( clk ), .D ( new_AGEMA_signal_13631 ), .Q ( new_AGEMA_signal_13632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5614 ( .C ( clk ), .D ( new_AGEMA_signal_13641 ), .Q ( new_AGEMA_signal_13642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5624 ( .C ( clk ), .D ( new_AGEMA_signal_13651 ), .Q ( new_AGEMA_signal_13652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5632 ( .C ( clk ), .D ( new_AGEMA_signal_13659 ), .Q ( new_AGEMA_signal_13660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5640 ( .C ( clk ), .D ( new_AGEMA_signal_13667 ), .Q ( new_AGEMA_signal_13668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5648 ( .C ( clk ), .D ( new_AGEMA_signal_13675 ), .Q ( new_AGEMA_signal_13676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5656 ( .C ( clk ), .D ( new_AGEMA_signal_13683 ), .Q ( new_AGEMA_signal_13684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5728 ( .C ( clk ), .D ( new_AGEMA_signal_13755 ), .Q ( new_AGEMA_signal_13756 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5736 ( .C ( clk ), .D ( new_AGEMA_signal_13763 ), .Q ( new_AGEMA_signal_13764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5744 ( .C ( clk ), .D ( new_AGEMA_signal_13771 ), .Q ( new_AGEMA_signal_13772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5752 ( .C ( clk ), .D ( new_AGEMA_signal_13779 ), .Q ( new_AGEMA_signal_13780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5792 ( .C ( clk ), .D ( new_AGEMA_signal_13819 ), .Q ( new_AGEMA_signal_13820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5800 ( .C ( clk ), .D ( new_AGEMA_signal_13827 ), .Q ( new_AGEMA_signal_13828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5808 ( .C ( clk ), .D ( new_AGEMA_signal_13835 ), .Q ( new_AGEMA_signal_13836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5816 ( .C ( clk ), .D ( new_AGEMA_signal_13843 ), .Q ( new_AGEMA_signal_13844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5968 ( .C ( clk ), .D ( new_AGEMA_signal_13995 ), .Q ( new_AGEMA_signal_13996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5978 ( .C ( clk ), .D ( new_AGEMA_signal_14005 ), .Q ( new_AGEMA_signal_14006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5988 ( .C ( clk ), .D ( new_AGEMA_signal_14015 ), .Q ( new_AGEMA_signal_14016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5998 ( .C ( clk ), .D ( new_AGEMA_signal_14025 ), .Q ( new_AGEMA_signal_14026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6328 ( .C ( clk ), .D ( new_AGEMA_signal_14355 ), .Q ( new_AGEMA_signal_14356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6340 ( .C ( clk ), .D ( new_AGEMA_signal_14367 ), .Q ( new_AGEMA_signal_14368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6352 ( .C ( clk ), .D ( new_AGEMA_signal_14379 ), .Q ( new_AGEMA_signal_14380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6364 ( .C ( clk ), .D ( new_AGEMA_signal_14391 ), .Q ( new_AGEMA_signal_14392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6378 ( .C ( clk ), .D ( new_AGEMA_signal_14405 ), .Q ( new_AGEMA_signal_14406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6392 ( .C ( clk ), .D ( new_AGEMA_signal_14419 ), .Q ( new_AGEMA_signal_14420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6406 ( .C ( clk ), .D ( new_AGEMA_signal_14433 ), .Q ( new_AGEMA_signal_14434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6420 ( .C ( clk ), .D ( new_AGEMA_signal_14447 ), .Q ( new_AGEMA_signal_14448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6466 ( .C ( clk ), .D ( new_AGEMA_signal_14493 ), .Q ( new_AGEMA_signal_14494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6480 ( .C ( clk ), .D ( new_AGEMA_signal_14507 ), .Q ( new_AGEMA_signal_14508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6494 ( .C ( clk ), .D ( new_AGEMA_signal_14521 ), .Q ( new_AGEMA_signal_14522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6508 ( .C ( clk ), .D ( new_AGEMA_signal_14535 ), .Q ( new_AGEMA_signal_14536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6610 ( .C ( clk ), .D ( new_AGEMA_signal_14637 ), .Q ( new_AGEMA_signal_14638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6626 ( .C ( clk ), .D ( new_AGEMA_signal_14653 ), .Q ( new_AGEMA_signal_14654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6642 ( .C ( clk ), .D ( new_AGEMA_signal_14669 ), .Q ( new_AGEMA_signal_14670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6658 ( .C ( clk ), .D ( new_AGEMA_signal_14685 ), .Q ( new_AGEMA_signal_14686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6698 ( .C ( clk ), .D ( new_AGEMA_signal_14725 ), .Q ( new_AGEMA_signal_14726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6714 ( .C ( clk ), .D ( new_AGEMA_signal_14741 ), .Q ( new_AGEMA_signal_14742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6730 ( .C ( clk ), .D ( new_AGEMA_signal_14757 ), .Q ( new_AGEMA_signal_14758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6746 ( .C ( clk ), .D ( new_AGEMA_signal_14773 ), .Q ( new_AGEMA_signal_14774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6896 ( .C ( clk ), .D ( new_AGEMA_signal_14923 ), .Q ( new_AGEMA_signal_14924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6912 ( .C ( clk ), .D ( new_AGEMA_signal_14939 ), .Q ( new_AGEMA_signal_14940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6928 ( .C ( clk ), .D ( new_AGEMA_signal_14955 ), .Q ( new_AGEMA_signal_14956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6944 ( .C ( clk ), .D ( new_AGEMA_signal_14971 ), .Q ( new_AGEMA_signal_14972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7002 ( .C ( clk ), .D ( new_AGEMA_signal_15029 ), .Q ( new_AGEMA_signal_15030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7020 ( .C ( clk ), .D ( new_AGEMA_signal_15047 ), .Q ( new_AGEMA_signal_15048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7038 ( .C ( clk ), .D ( new_AGEMA_signal_15065 ), .Q ( new_AGEMA_signal_15066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7056 ( .C ( clk ), .D ( new_AGEMA_signal_15083 ), .Q ( new_AGEMA_signal_15084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7202 ( .C ( clk ), .D ( new_AGEMA_signal_15229 ), .Q ( new_AGEMA_signal_15230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7222 ( .C ( clk ), .D ( new_AGEMA_signal_15249 ), .Q ( new_AGEMA_signal_15250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7242 ( .C ( clk ), .D ( new_AGEMA_signal_15269 ), .Q ( new_AGEMA_signal_15270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7262 ( .C ( clk ), .D ( new_AGEMA_signal_15289 ), .Q ( new_AGEMA_signal_15290 ) ) ;

    /* cells in depth 11 */
    buf_clk new_AGEMA_reg_buffer_4023 ( .C ( clk ), .D ( n1934 ), .Q ( new_AGEMA_signal_12051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4025 ( .C ( clk ), .D ( new_AGEMA_signal_2871 ), .Q ( new_AGEMA_signal_12053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4027 ( .C ( clk ), .D ( new_AGEMA_signal_2872 ), .Q ( new_AGEMA_signal_12055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4029 ( .C ( clk ), .D ( new_AGEMA_signal_2873 ), .Q ( new_AGEMA_signal_12057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4037 ( .C ( clk ), .D ( new_AGEMA_signal_12064 ), .Q ( new_AGEMA_signal_12065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4045 ( .C ( clk ), .D ( new_AGEMA_signal_12072 ), .Q ( new_AGEMA_signal_12073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4053 ( .C ( clk ), .D ( new_AGEMA_signal_12080 ), .Q ( new_AGEMA_signal_12081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4061 ( .C ( clk ), .D ( new_AGEMA_signal_12088 ), .Q ( new_AGEMA_signal_12089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4063 ( .C ( clk ), .D ( n1981 ), .Q ( new_AGEMA_signal_12091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4065 ( .C ( clk ), .D ( new_AGEMA_signal_2895 ), .Q ( new_AGEMA_signal_12093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4067 ( .C ( clk ), .D ( new_AGEMA_signal_2896 ), .Q ( new_AGEMA_signal_12095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4069 ( .C ( clk ), .D ( new_AGEMA_signal_2897 ), .Q ( new_AGEMA_signal_12097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4073 ( .C ( clk ), .D ( new_AGEMA_signal_12100 ), .Q ( new_AGEMA_signal_12101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4077 ( .C ( clk ), .D ( new_AGEMA_signal_12104 ), .Q ( new_AGEMA_signal_12105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4081 ( .C ( clk ), .D ( new_AGEMA_signal_12108 ), .Q ( new_AGEMA_signal_12109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4085 ( .C ( clk ), .D ( new_AGEMA_signal_12112 ), .Q ( new_AGEMA_signal_12113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4093 ( .C ( clk ), .D ( new_AGEMA_signal_12120 ), .Q ( new_AGEMA_signal_12121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4101 ( .C ( clk ), .D ( new_AGEMA_signal_12128 ), .Q ( new_AGEMA_signal_12129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4109 ( .C ( clk ), .D ( new_AGEMA_signal_12136 ), .Q ( new_AGEMA_signal_12137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4117 ( .C ( clk ), .D ( new_AGEMA_signal_12144 ), .Q ( new_AGEMA_signal_12145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4119 ( .C ( clk ), .D ( new_AGEMA_signal_11202 ), .Q ( new_AGEMA_signal_12147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4121 ( .C ( clk ), .D ( new_AGEMA_signal_11210 ), .Q ( new_AGEMA_signal_12149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4123 ( .C ( clk ), .D ( new_AGEMA_signal_11218 ), .Q ( new_AGEMA_signal_12151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4125 ( .C ( clk ), .D ( new_AGEMA_signal_11226 ), .Q ( new_AGEMA_signal_12153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4131 ( .C ( clk ), .D ( new_AGEMA_signal_12158 ), .Q ( new_AGEMA_signal_12159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4137 ( .C ( clk ), .D ( new_AGEMA_signal_12164 ), .Q ( new_AGEMA_signal_12165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4143 ( .C ( clk ), .D ( new_AGEMA_signal_12170 ), .Q ( new_AGEMA_signal_12171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4149 ( .C ( clk ), .D ( new_AGEMA_signal_12176 ), .Q ( new_AGEMA_signal_12177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4153 ( .C ( clk ), .D ( new_AGEMA_signal_12180 ), .Q ( new_AGEMA_signal_12181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4157 ( .C ( clk ), .D ( new_AGEMA_signal_12184 ), .Q ( new_AGEMA_signal_12185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4161 ( .C ( clk ), .D ( new_AGEMA_signal_12188 ), .Q ( new_AGEMA_signal_12189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4165 ( .C ( clk ), .D ( new_AGEMA_signal_12192 ), .Q ( new_AGEMA_signal_12193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4173 ( .C ( clk ), .D ( new_AGEMA_signal_12200 ), .Q ( new_AGEMA_signal_12201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4181 ( .C ( clk ), .D ( new_AGEMA_signal_12208 ), .Q ( new_AGEMA_signal_12209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4189 ( .C ( clk ), .D ( new_AGEMA_signal_12216 ), .Q ( new_AGEMA_signal_12217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4197 ( .C ( clk ), .D ( new_AGEMA_signal_12224 ), .Q ( new_AGEMA_signal_12225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4201 ( .C ( clk ), .D ( new_AGEMA_signal_12228 ), .Q ( new_AGEMA_signal_12229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4205 ( .C ( clk ), .D ( new_AGEMA_signal_12232 ), .Q ( new_AGEMA_signal_12233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4209 ( .C ( clk ), .D ( new_AGEMA_signal_12236 ), .Q ( new_AGEMA_signal_12237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4213 ( .C ( clk ), .D ( new_AGEMA_signal_12240 ), .Q ( new_AGEMA_signal_12241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4219 ( .C ( clk ), .D ( new_AGEMA_signal_12246 ), .Q ( new_AGEMA_signal_12247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4225 ( .C ( clk ), .D ( new_AGEMA_signal_12252 ), .Q ( new_AGEMA_signal_12253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4231 ( .C ( clk ), .D ( new_AGEMA_signal_12258 ), .Q ( new_AGEMA_signal_12259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4237 ( .C ( clk ), .D ( new_AGEMA_signal_12264 ), .Q ( new_AGEMA_signal_12265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4243 ( .C ( clk ), .D ( new_AGEMA_signal_12270 ), .Q ( new_AGEMA_signal_12271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4249 ( .C ( clk ), .D ( new_AGEMA_signal_12276 ), .Q ( new_AGEMA_signal_12277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4255 ( .C ( clk ), .D ( new_AGEMA_signal_12282 ), .Q ( new_AGEMA_signal_12283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4261 ( .C ( clk ), .D ( new_AGEMA_signal_12288 ), .Q ( new_AGEMA_signal_12289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4267 ( .C ( clk ), .D ( new_AGEMA_signal_12294 ), .Q ( new_AGEMA_signal_12295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4273 ( .C ( clk ), .D ( new_AGEMA_signal_12300 ), .Q ( new_AGEMA_signal_12301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4279 ( .C ( clk ), .D ( new_AGEMA_signal_12306 ), .Q ( new_AGEMA_signal_12307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4285 ( .C ( clk ), .D ( new_AGEMA_signal_12312 ), .Q ( new_AGEMA_signal_12313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4291 ( .C ( clk ), .D ( new_AGEMA_signal_12318 ), .Q ( new_AGEMA_signal_12319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4297 ( .C ( clk ), .D ( new_AGEMA_signal_12324 ), .Q ( new_AGEMA_signal_12325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4303 ( .C ( clk ), .D ( new_AGEMA_signal_12330 ), .Q ( new_AGEMA_signal_12331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4309 ( .C ( clk ), .D ( new_AGEMA_signal_12336 ), .Q ( new_AGEMA_signal_12337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4315 ( .C ( clk ), .D ( new_AGEMA_signal_12342 ), .Q ( new_AGEMA_signal_12343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4321 ( .C ( clk ), .D ( new_AGEMA_signal_12348 ), .Q ( new_AGEMA_signal_12349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4327 ( .C ( clk ), .D ( new_AGEMA_signal_12354 ), .Q ( new_AGEMA_signal_12355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4333 ( .C ( clk ), .D ( new_AGEMA_signal_12360 ), .Q ( new_AGEMA_signal_12361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4337 ( .C ( clk ), .D ( new_AGEMA_signal_12364 ), .Q ( new_AGEMA_signal_12365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4341 ( .C ( clk ), .D ( new_AGEMA_signal_12368 ), .Q ( new_AGEMA_signal_12369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4345 ( .C ( clk ), .D ( new_AGEMA_signal_12372 ), .Q ( new_AGEMA_signal_12373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4349 ( .C ( clk ), .D ( new_AGEMA_signal_12376 ), .Q ( new_AGEMA_signal_12377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4357 ( .C ( clk ), .D ( new_AGEMA_signal_12384 ), .Q ( new_AGEMA_signal_12385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4365 ( .C ( clk ), .D ( new_AGEMA_signal_12392 ), .Q ( new_AGEMA_signal_12393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4373 ( .C ( clk ), .D ( new_AGEMA_signal_12400 ), .Q ( new_AGEMA_signal_12401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4381 ( .C ( clk ), .D ( new_AGEMA_signal_12408 ), .Q ( new_AGEMA_signal_12409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4385 ( .C ( clk ), .D ( new_AGEMA_signal_12412 ), .Q ( new_AGEMA_signal_12413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4389 ( .C ( clk ), .D ( new_AGEMA_signal_12416 ), .Q ( new_AGEMA_signal_12417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4393 ( .C ( clk ), .D ( new_AGEMA_signal_12420 ), .Q ( new_AGEMA_signal_12421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4397 ( .C ( clk ), .D ( new_AGEMA_signal_12424 ), .Q ( new_AGEMA_signal_12425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4403 ( .C ( clk ), .D ( new_AGEMA_signal_12430 ), .Q ( new_AGEMA_signal_12431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4409 ( .C ( clk ), .D ( new_AGEMA_signal_12436 ), .Q ( new_AGEMA_signal_12437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4415 ( .C ( clk ), .D ( new_AGEMA_signal_12442 ), .Q ( new_AGEMA_signal_12443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4421 ( .C ( clk ), .D ( new_AGEMA_signal_12448 ), .Q ( new_AGEMA_signal_12449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4429 ( .C ( clk ), .D ( new_AGEMA_signal_12456 ), .Q ( new_AGEMA_signal_12457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4437 ( .C ( clk ), .D ( new_AGEMA_signal_12464 ), .Q ( new_AGEMA_signal_12465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4445 ( .C ( clk ), .D ( new_AGEMA_signal_12472 ), .Q ( new_AGEMA_signal_12473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4453 ( .C ( clk ), .D ( new_AGEMA_signal_12480 ), .Q ( new_AGEMA_signal_12481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4455 ( .C ( clk ), .D ( new_AGEMA_signal_11764 ), .Q ( new_AGEMA_signal_12483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4457 ( .C ( clk ), .D ( new_AGEMA_signal_11766 ), .Q ( new_AGEMA_signal_12485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4459 ( .C ( clk ), .D ( new_AGEMA_signal_11768 ), .Q ( new_AGEMA_signal_12487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4461 ( .C ( clk ), .D ( new_AGEMA_signal_11770 ), .Q ( new_AGEMA_signal_12489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4467 ( .C ( clk ), .D ( new_AGEMA_signal_12494 ), .Q ( new_AGEMA_signal_12495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4473 ( .C ( clk ), .D ( new_AGEMA_signal_12500 ), .Q ( new_AGEMA_signal_12501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4479 ( .C ( clk ), .D ( new_AGEMA_signal_12506 ), .Q ( new_AGEMA_signal_12507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4485 ( .C ( clk ), .D ( new_AGEMA_signal_12512 ), .Q ( new_AGEMA_signal_12513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4487 ( .C ( clk ), .D ( n2410 ), .Q ( new_AGEMA_signal_12515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4489 ( .C ( clk ), .D ( new_AGEMA_signal_3012 ), .Q ( new_AGEMA_signal_12517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4491 ( .C ( clk ), .D ( new_AGEMA_signal_3013 ), .Q ( new_AGEMA_signal_12519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4493 ( .C ( clk ), .D ( new_AGEMA_signal_3014 ), .Q ( new_AGEMA_signal_12521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4495 ( .C ( clk ), .D ( n2421 ), .Q ( new_AGEMA_signal_12523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4497 ( .C ( clk ), .D ( new_AGEMA_signal_3015 ), .Q ( new_AGEMA_signal_12525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4499 ( .C ( clk ), .D ( new_AGEMA_signal_3016 ), .Q ( new_AGEMA_signal_12527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4501 ( .C ( clk ), .D ( new_AGEMA_signal_3017 ), .Q ( new_AGEMA_signal_12529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4507 ( .C ( clk ), .D ( new_AGEMA_signal_12534 ), .Q ( new_AGEMA_signal_12535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4513 ( .C ( clk ), .D ( new_AGEMA_signal_12540 ), .Q ( new_AGEMA_signal_12541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4519 ( .C ( clk ), .D ( new_AGEMA_signal_12546 ), .Q ( new_AGEMA_signal_12547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4525 ( .C ( clk ), .D ( new_AGEMA_signal_12552 ), .Q ( new_AGEMA_signal_12553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4531 ( .C ( clk ), .D ( new_AGEMA_signal_12558 ), .Q ( new_AGEMA_signal_12559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4537 ( .C ( clk ), .D ( new_AGEMA_signal_12564 ), .Q ( new_AGEMA_signal_12565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4543 ( .C ( clk ), .D ( new_AGEMA_signal_12570 ), .Q ( new_AGEMA_signal_12571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4549 ( .C ( clk ), .D ( new_AGEMA_signal_12576 ), .Q ( new_AGEMA_signal_12577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4557 ( .C ( clk ), .D ( new_AGEMA_signal_12584 ), .Q ( new_AGEMA_signal_12585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4565 ( .C ( clk ), .D ( new_AGEMA_signal_12592 ), .Q ( new_AGEMA_signal_12593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4573 ( .C ( clk ), .D ( new_AGEMA_signal_12600 ), .Q ( new_AGEMA_signal_12601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4581 ( .C ( clk ), .D ( new_AGEMA_signal_12608 ), .Q ( new_AGEMA_signal_12609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4589 ( .C ( clk ), .D ( new_AGEMA_signal_12616 ), .Q ( new_AGEMA_signal_12617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4597 ( .C ( clk ), .D ( new_AGEMA_signal_12624 ), .Q ( new_AGEMA_signal_12625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4605 ( .C ( clk ), .D ( new_AGEMA_signal_12632 ), .Q ( new_AGEMA_signal_12633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4613 ( .C ( clk ), .D ( new_AGEMA_signal_12640 ), .Q ( new_AGEMA_signal_12641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4619 ( .C ( clk ), .D ( new_AGEMA_signal_12646 ), .Q ( new_AGEMA_signal_12647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4625 ( .C ( clk ), .D ( new_AGEMA_signal_12652 ), .Q ( new_AGEMA_signal_12653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4631 ( .C ( clk ), .D ( new_AGEMA_signal_12658 ), .Q ( new_AGEMA_signal_12659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4637 ( .C ( clk ), .D ( new_AGEMA_signal_12664 ), .Q ( new_AGEMA_signal_12665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4643 ( .C ( clk ), .D ( new_AGEMA_signal_12670 ), .Q ( new_AGEMA_signal_12671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4649 ( .C ( clk ), .D ( new_AGEMA_signal_12676 ), .Q ( new_AGEMA_signal_12677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4655 ( .C ( clk ), .D ( new_AGEMA_signal_12682 ), .Q ( new_AGEMA_signal_12683 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4661 ( .C ( clk ), .D ( new_AGEMA_signal_12688 ), .Q ( new_AGEMA_signal_12689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4663 ( .C ( clk ), .D ( new_AGEMA_signal_11726 ), .Q ( new_AGEMA_signal_12691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4665 ( .C ( clk ), .D ( new_AGEMA_signal_11730 ), .Q ( new_AGEMA_signal_12693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4667 ( .C ( clk ), .D ( new_AGEMA_signal_11734 ), .Q ( new_AGEMA_signal_12695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4669 ( .C ( clk ), .D ( new_AGEMA_signal_11738 ), .Q ( new_AGEMA_signal_12697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4673 ( .C ( clk ), .D ( new_AGEMA_signal_12700 ), .Q ( new_AGEMA_signal_12701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4677 ( .C ( clk ), .D ( new_AGEMA_signal_12704 ), .Q ( new_AGEMA_signal_12705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4681 ( .C ( clk ), .D ( new_AGEMA_signal_12708 ), .Q ( new_AGEMA_signal_12709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4685 ( .C ( clk ), .D ( new_AGEMA_signal_12712 ), .Q ( new_AGEMA_signal_12713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4689 ( .C ( clk ), .D ( new_AGEMA_signal_12716 ), .Q ( new_AGEMA_signal_12717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4693 ( .C ( clk ), .D ( new_AGEMA_signal_12720 ), .Q ( new_AGEMA_signal_12721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4697 ( .C ( clk ), .D ( new_AGEMA_signal_12724 ), .Q ( new_AGEMA_signal_12725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4701 ( .C ( clk ), .D ( new_AGEMA_signal_12728 ), .Q ( new_AGEMA_signal_12729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4705 ( .C ( clk ), .D ( new_AGEMA_signal_12732 ), .Q ( new_AGEMA_signal_12733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4709 ( .C ( clk ), .D ( new_AGEMA_signal_12736 ), .Q ( new_AGEMA_signal_12737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4713 ( .C ( clk ), .D ( new_AGEMA_signal_12740 ), .Q ( new_AGEMA_signal_12741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4717 ( .C ( clk ), .D ( new_AGEMA_signal_12744 ), .Q ( new_AGEMA_signal_12745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4719 ( .C ( clk ), .D ( new_AGEMA_signal_11506 ), .Q ( new_AGEMA_signal_12747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4721 ( .C ( clk ), .D ( new_AGEMA_signal_11514 ), .Q ( new_AGEMA_signal_12749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4723 ( .C ( clk ), .D ( new_AGEMA_signal_11522 ), .Q ( new_AGEMA_signal_12751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4725 ( .C ( clk ), .D ( new_AGEMA_signal_11530 ), .Q ( new_AGEMA_signal_12753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4729 ( .C ( clk ), .D ( new_AGEMA_signal_12756 ), .Q ( new_AGEMA_signal_12757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4735 ( .C ( clk ), .D ( new_AGEMA_signal_12762 ), .Q ( new_AGEMA_signal_12763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4741 ( .C ( clk ), .D ( new_AGEMA_signal_12768 ), .Q ( new_AGEMA_signal_12769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4747 ( .C ( clk ), .D ( new_AGEMA_signal_12774 ), .Q ( new_AGEMA_signal_12775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4759 ( .C ( clk ), .D ( n1984 ), .Q ( new_AGEMA_signal_12787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4763 ( .C ( clk ), .D ( new_AGEMA_signal_3123 ), .Q ( new_AGEMA_signal_12791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4767 ( .C ( clk ), .D ( new_AGEMA_signal_3124 ), .Q ( new_AGEMA_signal_12795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4771 ( .C ( clk ), .D ( new_AGEMA_signal_3125 ), .Q ( new_AGEMA_signal_12799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4779 ( .C ( clk ), .D ( new_AGEMA_signal_12806 ), .Q ( new_AGEMA_signal_12807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4787 ( .C ( clk ), .D ( new_AGEMA_signal_12814 ), .Q ( new_AGEMA_signal_12815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4795 ( .C ( clk ), .D ( new_AGEMA_signal_12822 ), .Q ( new_AGEMA_signal_12823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4803 ( .C ( clk ), .D ( new_AGEMA_signal_12830 ), .Q ( new_AGEMA_signal_12831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4811 ( .C ( clk ), .D ( new_AGEMA_signal_12838 ), .Q ( new_AGEMA_signal_12839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4819 ( .C ( clk ), .D ( new_AGEMA_signal_12846 ), .Q ( new_AGEMA_signal_12847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4827 ( .C ( clk ), .D ( new_AGEMA_signal_12854 ), .Q ( new_AGEMA_signal_12855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4835 ( .C ( clk ), .D ( new_AGEMA_signal_12862 ), .Q ( new_AGEMA_signal_12863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4843 ( .C ( clk ), .D ( new_AGEMA_signal_12870 ), .Q ( new_AGEMA_signal_12871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4851 ( .C ( clk ), .D ( new_AGEMA_signal_12878 ), .Q ( new_AGEMA_signal_12879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4859 ( .C ( clk ), .D ( new_AGEMA_signal_12886 ), .Q ( new_AGEMA_signal_12887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4867 ( .C ( clk ), .D ( new_AGEMA_signal_12894 ), .Q ( new_AGEMA_signal_12895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4875 ( .C ( clk ), .D ( new_AGEMA_signal_12902 ), .Q ( new_AGEMA_signal_12903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4883 ( .C ( clk ), .D ( new_AGEMA_signal_12910 ), .Q ( new_AGEMA_signal_12911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4891 ( .C ( clk ), .D ( new_AGEMA_signal_12918 ), .Q ( new_AGEMA_signal_12919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4899 ( .C ( clk ), .D ( new_AGEMA_signal_12926 ), .Q ( new_AGEMA_signal_12927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4905 ( .C ( clk ), .D ( new_AGEMA_signal_12932 ), .Q ( new_AGEMA_signal_12933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4911 ( .C ( clk ), .D ( new_AGEMA_signal_12938 ), .Q ( new_AGEMA_signal_12939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4917 ( .C ( clk ), .D ( new_AGEMA_signal_12944 ), .Q ( new_AGEMA_signal_12945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4923 ( .C ( clk ), .D ( new_AGEMA_signal_12950 ), .Q ( new_AGEMA_signal_12951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4933 ( .C ( clk ), .D ( new_AGEMA_signal_12960 ), .Q ( new_AGEMA_signal_12961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4943 ( .C ( clk ), .D ( new_AGEMA_signal_12970 ), .Q ( new_AGEMA_signal_12971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4953 ( .C ( clk ), .D ( new_AGEMA_signal_12980 ), .Q ( new_AGEMA_signal_12981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4963 ( .C ( clk ), .D ( new_AGEMA_signal_12990 ), .Q ( new_AGEMA_signal_12991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4971 ( .C ( clk ), .D ( new_AGEMA_signal_12998 ), .Q ( new_AGEMA_signal_12999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4979 ( .C ( clk ), .D ( new_AGEMA_signal_13006 ), .Q ( new_AGEMA_signal_13007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4987 ( .C ( clk ), .D ( new_AGEMA_signal_13014 ), .Q ( new_AGEMA_signal_13015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4995 ( .C ( clk ), .D ( new_AGEMA_signal_13022 ), .Q ( new_AGEMA_signal_13023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5003 ( .C ( clk ), .D ( new_AGEMA_signal_13030 ), .Q ( new_AGEMA_signal_13031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5011 ( .C ( clk ), .D ( new_AGEMA_signal_13038 ), .Q ( new_AGEMA_signal_13039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5019 ( .C ( clk ), .D ( new_AGEMA_signal_13046 ), .Q ( new_AGEMA_signal_13047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5027 ( .C ( clk ), .D ( new_AGEMA_signal_13054 ), .Q ( new_AGEMA_signal_13055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5035 ( .C ( clk ), .D ( new_AGEMA_signal_13062 ), .Q ( new_AGEMA_signal_13063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5043 ( .C ( clk ), .D ( new_AGEMA_signal_13070 ), .Q ( new_AGEMA_signal_13071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5051 ( .C ( clk ), .D ( new_AGEMA_signal_13078 ), .Q ( new_AGEMA_signal_13079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5059 ( .C ( clk ), .D ( new_AGEMA_signal_13086 ), .Q ( new_AGEMA_signal_13087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5071 ( .C ( clk ), .D ( new_AGEMA_signal_11750 ), .Q ( new_AGEMA_signal_13099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5075 ( .C ( clk ), .D ( new_AGEMA_signal_11754 ), .Q ( new_AGEMA_signal_13103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5079 ( .C ( clk ), .D ( new_AGEMA_signal_11758 ), .Q ( new_AGEMA_signal_13107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5083 ( .C ( clk ), .D ( new_AGEMA_signal_11762 ), .Q ( new_AGEMA_signal_13111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5089 ( .C ( clk ), .D ( new_AGEMA_signal_13116 ), .Q ( new_AGEMA_signal_13117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5095 ( .C ( clk ), .D ( new_AGEMA_signal_13122 ), .Q ( new_AGEMA_signal_13123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5101 ( .C ( clk ), .D ( new_AGEMA_signal_13128 ), .Q ( new_AGEMA_signal_13129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5107 ( .C ( clk ), .D ( new_AGEMA_signal_13134 ), .Q ( new_AGEMA_signal_13135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5111 ( .C ( clk ), .D ( new_AGEMA_signal_11304 ), .Q ( new_AGEMA_signal_13139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5115 ( .C ( clk ), .D ( new_AGEMA_signal_11310 ), .Q ( new_AGEMA_signal_13143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5119 ( .C ( clk ), .D ( new_AGEMA_signal_11316 ), .Q ( new_AGEMA_signal_13147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5123 ( .C ( clk ), .D ( new_AGEMA_signal_11322 ), .Q ( new_AGEMA_signal_13151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5133 ( .C ( clk ), .D ( new_AGEMA_signal_13160 ), .Q ( new_AGEMA_signal_13161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5143 ( .C ( clk ), .D ( new_AGEMA_signal_13170 ), .Q ( new_AGEMA_signal_13171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5153 ( .C ( clk ), .D ( new_AGEMA_signal_13180 ), .Q ( new_AGEMA_signal_13181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5163 ( .C ( clk ), .D ( new_AGEMA_signal_13190 ), .Q ( new_AGEMA_signal_13191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5171 ( .C ( clk ), .D ( new_AGEMA_signal_13198 ), .Q ( new_AGEMA_signal_13199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5179 ( .C ( clk ), .D ( new_AGEMA_signal_13206 ), .Q ( new_AGEMA_signal_13207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5187 ( .C ( clk ), .D ( new_AGEMA_signal_13214 ), .Q ( new_AGEMA_signal_13215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C ( clk ), .D ( new_AGEMA_signal_13222 ), .Q ( new_AGEMA_signal_13223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C ( clk ), .D ( n2478 ), .Q ( new_AGEMA_signal_13227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C ( clk ), .D ( new_AGEMA_signal_2775 ), .Q ( new_AGEMA_signal_13231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C ( clk ), .D ( new_AGEMA_signal_2776 ), .Q ( new_AGEMA_signal_13235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C ( clk ), .D ( new_AGEMA_signal_2777 ), .Q ( new_AGEMA_signal_13239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C ( clk ), .D ( new_AGEMA_signal_13254 ), .Q ( new_AGEMA_signal_13255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C ( clk ), .D ( new_AGEMA_signal_13262 ), .Q ( new_AGEMA_signal_13263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C ( clk ), .D ( new_AGEMA_signal_13270 ), .Q ( new_AGEMA_signal_13271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C ( clk ), .D ( new_AGEMA_signal_13278 ), .Q ( new_AGEMA_signal_13279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5259 ( .C ( clk ), .D ( new_AGEMA_signal_13286 ), .Q ( new_AGEMA_signal_13287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5267 ( .C ( clk ), .D ( new_AGEMA_signal_13294 ), .Q ( new_AGEMA_signal_13295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5275 ( .C ( clk ), .D ( new_AGEMA_signal_13302 ), .Q ( new_AGEMA_signal_13303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5283 ( .C ( clk ), .D ( new_AGEMA_signal_13310 ), .Q ( new_AGEMA_signal_13311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5289 ( .C ( clk ), .D ( new_AGEMA_signal_13316 ), .Q ( new_AGEMA_signal_13317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5295 ( .C ( clk ), .D ( new_AGEMA_signal_13322 ), .Q ( new_AGEMA_signal_13323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5301 ( .C ( clk ), .D ( new_AGEMA_signal_13328 ), .Q ( new_AGEMA_signal_13329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5307 ( .C ( clk ), .D ( new_AGEMA_signal_13334 ), .Q ( new_AGEMA_signal_13335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5311 ( .C ( clk ), .D ( n2660 ), .Q ( new_AGEMA_signal_13339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5315 ( .C ( clk ), .D ( new_AGEMA_signal_3075 ), .Q ( new_AGEMA_signal_13343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5319 ( .C ( clk ), .D ( new_AGEMA_signal_3076 ), .Q ( new_AGEMA_signal_13347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5323 ( .C ( clk ), .D ( new_AGEMA_signal_3077 ), .Q ( new_AGEMA_signal_13351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5331 ( .C ( clk ), .D ( new_AGEMA_signal_13358 ), .Q ( new_AGEMA_signal_13359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5339 ( .C ( clk ), .D ( new_AGEMA_signal_13366 ), .Q ( new_AGEMA_signal_13367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5347 ( .C ( clk ), .D ( new_AGEMA_signal_13374 ), .Q ( new_AGEMA_signal_13375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5355 ( .C ( clk ), .D ( new_AGEMA_signal_13382 ), .Q ( new_AGEMA_signal_13383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5367 ( .C ( clk ), .D ( n1940 ), .Q ( new_AGEMA_signal_13395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5373 ( .C ( clk ), .D ( new_AGEMA_signal_2877 ), .Q ( new_AGEMA_signal_13401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5379 ( .C ( clk ), .D ( new_AGEMA_signal_2878 ), .Q ( new_AGEMA_signal_13407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5385 ( .C ( clk ), .D ( new_AGEMA_signal_2879 ), .Q ( new_AGEMA_signal_13413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5391 ( .C ( clk ), .D ( n1961 ), .Q ( new_AGEMA_signal_13419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5397 ( .C ( clk ), .D ( new_AGEMA_signal_2880 ), .Q ( new_AGEMA_signal_13425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5403 ( .C ( clk ), .D ( new_AGEMA_signal_2881 ), .Q ( new_AGEMA_signal_13431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5409 ( .C ( clk ), .D ( new_AGEMA_signal_2882 ), .Q ( new_AGEMA_signal_13437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5415 ( .C ( clk ), .D ( n1987 ), .Q ( new_AGEMA_signal_13443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5421 ( .C ( clk ), .D ( new_AGEMA_signal_2571 ), .Q ( new_AGEMA_signal_13449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5427 ( .C ( clk ), .D ( new_AGEMA_signal_2572 ), .Q ( new_AGEMA_signal_13455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5433 ( .C ( clk ), .D ( new_AGEMA_signal_2573 ), .Q ( new_AGEMA_signal_13461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5457 ( .C ( clk ), .D ( new_AGEMA_signal_13484 ), .Q ( new_AGEMA_signal_13485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5465 ( .C ( clk ), .D ( new_AGEMA_signal_13492 ), .Q ( new_AGEMA_signal_13493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5473 ( .C ( clk ), .D ( new_AGEMA_signal_13500 ), .Q ( new_AGEMA_signal_13501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5481 ( .C ( clk ), .D ( new_AGEMA_signal_13508 ), .Q ( new_AGEMA_signal_13509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5487 ( .C ( clk ), .D ( n2054 ), .Q ( new_AGEMA_signal_13515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5493 ( .C ( clk ), .D ( new_AGEMA_signal_2910 ), .Q ( new_AGEMA_signal_13521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5499 ( .C ( clk ), .D ( new_AGEMA_signal_2911 ), .Q ( new_AGEMA_signal_13527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5505 ( .C ( clk ), .D ( new_AGEMA_signal_2912 ), .Q ( new_AGEMA_signal_13533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5529 ( .C ( clk ), .D ( new_AGEMA_signal_13556 ), .Q ( new_AGEMA_signal_13557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5537 ( .C ( clk ), .D ( new_AGEMA_signal_13564 ), .Q ( new_AGEMA_signal_13565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5545 ( .C ( clk ), .D ( new_AGEMA_signal_13572 ), .Q ( new_AGEMA_signal_13573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5553 ( .C ( clk ), .D ( new_AGEMA_signal_13580 ), .Q ( new_AGEMA_signal_13581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5561 ( .C ( clk ), .D ( new_AGEMA_signal_13588 ), .Q ( new_AGEMA_signal_13589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5569 ( .C ( clk ), .D ( new_AGEMA_signal_13596 ), .Q ( new_AGEMA_signal_13597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5577 ( .C ( clk ), .D ( new_AGEMA_signal_13604 ), .Q ( new_AGEMA_signal_13605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5585 ( .C ( clk ), .D ( new_AGEMA_signal_13612 ), .Q ( new_AGEMA_signal_13613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5595 ( .C ( clk ), .D ( new_AGEMA_signal_13622 ), .Q ( new_AGEMA_signal_13623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5605 ( .C ( clk ), .D ( new_AGEMA_signal_13632 ), .Q ( new_AGEMA_signal_13633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5615 ( .C ( clk ), .D ( new_AGEMA_signal_13642 ), .Q ( new_AGEMA_signal_13643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5625 ( .C ( clk ), .D ( new_AGEMA_signal_13652 ), .Q ( new_AGEMA_signal_13653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5633 ( .C ( clk ), .D ( new_AGEMA_signal_13660 ), .Q ( new_AGEMA_signal_13661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5641 ( .C ( clk ), .D ( new_AGEMA_signal_13668 ), .Q ( new_AGEMA_signal_13669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5649 ( .C ( clk ), .D ( new_AGEMA_signal_13676 ), .Q ( new_AGEMA_signal_13677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5657 ( .C ( clk ), .D ( new_AGEMA_signal_13684 ), .Q ( new_AGEMA_signal_13685 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5663 ( .C ( clk ), .D ( n2255 ), .Q ( new_AGEMA_signal_13691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5669 ( .C ( clk ), .D ( new_AGEMA_signal_2970 ), .Q ( new_AGEMA_signal_13697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5675 ( .C ( clk ), .D ( new_AGEMA_signal_2971 ), .Q ( new_AGEMA_signal_13703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5681 ( .C ( clk ), .D ( new_AGEMA_signal_2972 ), .Q ( new_AGEMA_signal_13709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5703 ( .C ( clk ), .D ( n2304 ), .Q ( new_AGEMA_signal_13731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5709 ( .C ( clk ), .D ( new_AGEMA_signal_2982 ), .Q ( new_AGEMA_signal_13737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5715 ( .C ( clk ), .D ( new_AGEMA_signal_2983 ), .Q ( new_AGEMA_signal_13743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5721 ( .C ( clk ), .D ( new_AGEMA_signal_2984 ), .Q ( new_AGEMA_signal_13749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5729 ( .C ( clk ), .D ( new_AGEMA_signal_13756 ), .Q ( new_AGEMA_signal_13757 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5737 ( .C ( clk ), .D ( new_AGEMA_signal_13764 ), .Q ( new_AGEMA_signal_13765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5745 ( .C ( clk ), .D ( new_AGEMA_signal_13772 ), .Q ( new_AGEMA_signal_13773 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5753 ( .C ( clk ), .D ( new_AGEMA_signal_13780 ), .Q ( new_AGEMA_signal_13781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5759 ( .C ( clk ), .D ( n2450 ), .Q ( new_AGEMA_signal_13787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5765 ( .C ( clk ), .D ( new_AGEMA_signal_3024 ), .Q ( new_AGEMA_signal_13793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5771 ( .C ( clk ), .D ( new_AGEMA_signal_3025 ), .Q ( new_AGEMA_signal_13799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5777 ( .C ( clk ), .D ( new_AGEMA_signal_3026 ), .Q ( new_AGEMA_signal_13805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5793 ( .C ( clk ), .D ( new_AGEMA_signal_13820 ), .Q ( new_AGEMA_signal_13821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5801 ( .C ( clk ), .D ( new_AGEMA_signal_13828 ), .Q ( new_AGEMA_signal_13829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5809 ( .C ( clk ), .D ( new_AGEMA_signal_13836 ), .Q ( new_AGEMA_signal_13837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5817 ( .C ( clk ), .D ( new_AGEMA_signal_13844 ), .Q ( new_AGEMA_signal_13845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5839 ( .C ( clk ), .D ( n2666 ), .Q ( new_AGEMA_signal_13867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5845 ( .C ( clk ), .D ( new_AGEMA_signal_3081 ), .Q ( new_AGEMA_signal_13873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5851 ( .C ( clk ), .D ( new_AGEMA_signal_3082 ), .Q ( new_AGEMA_signal_13879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5857 ( .C ( clk ), .D ( new_AGEMA_signal_3083 ), .Q ( new_AGEMA_signal_13885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5863 ( .C ( clk ), .D ( n2704 ), .Q ( new_AGEMA_signal_13891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5869 ( .C ( clk ), .D ( new_AGEMA_signal_3087 ), .Q ( new_AGEMA_signal_13897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5875 ( .C ( clk ), .D ( new_AGEMA_signal_3088 ), .Q ( new_AGEMA_signal_13903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5881 ( .C ( clk ), .D ( new_AGEMA_signal_3089 ), .Q ( new_AGEMA_signal_13909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5969 ( .C ( clk ), .D ( new_AGEMA_signal_13996 ), .Q ( new_AGEMA_signal_13997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5979 ( .C ( clk ), .D ( new_AGEMA_signal_14006 ), .Q ( new_AGEMA_signal_14007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5989 ( .C ( clk ), .D ( new_AGEMA_signal_14016 ), .Q ( new_AGEMA_signal_14017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5999 ( .C ( clk ), .D ( new_AGEMA_signal_14026 ), .Q ( new_AGEMA_signal_14027 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6087 ( .C ( clk ), .D ( n2280 ), .Q ( new_AGEMA_signal_14115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6095 ( .C ( clk ), .D ( new_AGEMA_signal_2694 ), .Q ( new_AGEMA_signal_14123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6103 ( .C ( clk ), .D ( new_AGEMA_signal_2695 ), .Q ( new_AGEMA_signal_14131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6111 ( .C ( clk ), .D ( new_AGEMA_signal_2696 ), .Q ( new_AGEMA_signal_14139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6143 ( .C ( clk ), .D ( new_AGEMA_signal_11292 ), .Q ( new_AGEMA_signal_14171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6151 ( .C ( clk ), .D ( new_AGEMA_signal_11294 ), .Q ( new_AGEMA_signal_14179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6159 ( .C ( clk ), .D ( new_AGEMA_signal_11296 ), .Q ( new_AGEMA_signal_14187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6167 ( .C ( clk ), .D ( new_AGEMA_signal_11298 ), .Q ( new_AGEMA_signal_14195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6175 ( .C ( clk ), .D ( n2456 ), .Q ( new_AGEMA_signal_14203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6183 ( .C ( clk ), .D ( new_AGEMA_signal_3027 ), .Q ( new_AGEMA_signal_14211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6191 ( .C ( clk ), .D ( new_AGEMA_signal_3028 ), .Q ( new_AGEMA_signal_14219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6199 ( .C ( clk ), .D ( new_AGEMA_signal_3029 ), .Q ( new_AGEMA_signal_14227 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6247 ( .C ( clk ), .D ( n2706 ), .Q ( new_AGEMA_signal_14275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6255 ( .C ( clk ), .D ( new_AGEMA_signal_3084 ), .Q ( new_AGEMA_signal_14283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6263 ( .C ( clk ), .D ( new_AGEMA_signal_3085 ), .Q ( new_AGEMA_signal_14291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6271 ( .C ( clk ), .D ( new_AGEMA_signal_3086 ), .Q ( new_AGEMA_signal_14299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6329 ( .C ( clk ), .D ( new_AGEMA_signal_14356 ), .Q ( new_AGEMA_signal_14357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6341 ( .C ( clk ), .D ( new_AGEMA_signal_14368 ), .Q ( new_AGEMA_signal_14369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6353 ( .C ( clk ), .D ( new_AGEMA_signal_14380 ), .Q ( new_AGEMA_signal_14381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6365 ( .C ( clk ), .D ( new_AGEMA_signal_14392 ), .Q ( new_AGEMA_signal_14393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6379 ( .C ( clk ), .D ( new_AGEMA_signal_14406 ), .Q ( new_AGEMA_signal_14407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6393 ( .C ( clk ), .D ( new_AGEMA_signal_14420 ), .Q ( new_AGEMA_signal_14421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6407 ( .C ( clk ), .D ( new_AGEMA_signal_14434 ), .Q ( new_AGEMA_signal_14435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6421 ( .C ( clk ), .D ( new_AGEMA_signal_14448 ), .Q ( new_AGEMA_signal_14449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6467 ( .C ( clk ), .D ( new_AGEMA_signal_14494 ), .Q ( new_AGEMA_signal_14495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6481 ( .C ( clk ), .D ( new_AGEMA_signal_14508 ), .Q ( new_AGEMA_signal_14509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6495 ( .C ( clk ), .D ( new_AGEMA_signal_14522 ), .Q ( new_AGEMA_signal_14523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6509 ( .C ( clk ), .D ( new_AGEMA_signal_14536 ), .Q ( new_AGEMA_signal_14537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6611 ( .C ( clk ), .D ( new_AGEMA_signal_14638 ), .Q ( new_AGEMA_signal_14639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6627 ( .C ( clk ), .D ( new_AGEMA_signal_14654 ), .Q ( new_AGEMA_signal_14655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6643 ( .C ( clk ), .D ( new_AGEMA_signal_14670 ), .Q ( new_AGEMA_signal_14671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6659 ( .C ( clk ), .D ( new_AGEMA_signal_14686 ), .Q ( new_AGEMA_signal_14687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6699 ( .C ( clk ), .D ( new_AGEMA_signal_14726 ), .Q ( new_AGEMA_signal_14727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6715 ( .C ( clk ), .D ( new_AGEMA_signal_14742 ), .Q ( new_AGEMA_signal_14743 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6731 ( .C ( clk ), .D ( new_AGEMA_signal_14758 ), .Q ( new_AGEMA_signal_14759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6747 ( .C ( clk ), .D ( new_AGEMA_signal_14774 ), .Q ( new_AGEMA_signal_14775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6897 ( .C ( clk ), .D ( new_AGEMA_signal_14924 ), .Q ( new_AGEMA_signal_14925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6913 ( .C ( clk ), .D ( new_AGEMA_signal_14940 ), .Q ( new_AGEMA_signal_14941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6929 ( .C ( clk ), .D ( new_AGEMA_signal_14956 ), .Q ( new_AGEMA_signal_14957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6945 ( .C ( clk ), .D ( new_AGEMA_signal_14972 ), .Q ( new_AGEMA_signal_14973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7003 ( .C ( clk ), .D ( new_AGEMA_signal_15030 ), .Q ( new_AGEMA_signal_15031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7021 ( .C ( clk ), .D ( new_AGEMA_signal_15048 ), .Q ( new_AGEMA_signal_15049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7039 ( .C ( clk ), .D ( new_AGEMA_signal_15066 ), .Q ( new_AGEMA_signal_15067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7057 ( .C ( clk ), .D ( new_AGEMA_signal_15084 ), .Q ( new_AGEMA_signal_15085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7203 ( .C ( clk ), .D ( new_AGEMA_signal_15230 ), .Q ( new_AGEMA_signal_15231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7223 ( .C ( clk ), .D ( new_AGEMA_signal_15250 ), .Q ( new_AGEMA_signal_15251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7243 ( .C ( clk ), .D ( new_AGEMA_signal_15270 ), .Q ( new_AGEMA_signal_15271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7263 ( .C ( clk ), .D ( new_AGEMA_signal_15290 ), .Q ( new_AGEMA_signal_15291 ) ) ;

    /* cells in depth 12 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2001 ( .a ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, n1932}), .b ({new_AGEMA_signal_11138, new_AGEMA_signal_11134, new_AGEMA_signal_11130, new_AGEMA_signal_11126}), .clk ( clk ), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, n1933}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2051 ( .a ({new_AGEMA_signal_11154, new_AGEMA_signal_11150, new_AGEMA_signal_11146, new_AGEMA_signal_11142}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, n1955}), .clk ( clk ), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, n1958}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2067 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, n1967}), .b ({new_AGEMA_signal_11186, new_AGEMA_signal_11178, new_AGEMA_signal_11170, new_AGEMA_signal_11162}), .clk ( clk ), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, n1990}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2104 ( .a ({new_AGEMA_signal_11194, new_AGEMA_signal_11192, new_AGEMA_signal_11190, new_AGEMA_signal_11188}), .b ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, n1977}), .clk ( clk ), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n1982}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2128 ( .a ({new_AGEMA_signal_11226, new_AGEMA_signal_11218, new_AGEMA_signal_11210, new_AGEMA_signal_11202}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, n1998}), .clk ( clk ), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, n1999}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2148 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, n2010}), .b ({new_AGEMA_signal_11250, new_AGEMA_signal_11244, new_AGEMA_signal_11238, new_AGEMA_signal_11232}), .clk ( clk ), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, new_AGEMA_signal_3132, n2011}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2165 ( .a ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, n2024}), .b ({new_AGEMA_signal_11266, new_AGEMA_signal_11262, new_AGEMA_signal_11258, new_AGEMA_signal_11254}), .clk ( clk ), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, n2025}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2179 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, n2035}), .b ({new_AGEMA_signal_11290, new_AGEMA_signal_11284, new_AGEMA_signal_11278, new_AGEMA_signal_11272}), .clk ( clk ), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2036}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2196 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, n2048}), .b ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, n2047}), .clk ( clk ), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, n2049}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2207 ( .a ({new_AGEMA_signal_11298, new_AGEMA_signal_11296, new_AGEMA_signal_11294, new_AGEMA_signal_11292}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, n2059}), .clk ( clk ), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({new_AGEMA_signal_3146, new_AGEMA_signal_3145, new_AGEMA_signal_3144, n2072}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2214 ( .a ({new_AGEMA_signal_11322, new_AGEMA_signal_11316, new_AGEMA_signal_11310, new_AGEMA_signal_11304}), .b ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, n2064}), .clk ( clk ), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, n2067}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2230 ( .a ({new_AGEMA_signal_11346, new_AGEMA_signal_11340, new_AGEMA_signal_11334, new_AGEMA_signal_11328}), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, n2077}), .clk ( clk ), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, n2078}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2250 ( .a ({new_AGEMA_signal_11354, new_AGEMA_signal_11352, new_AGEMA_signal_11350, new_AGEMA_signal_11348}), .b ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}), .clk ( clk ), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, n2097}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2257 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, n2095}), .b ({new_AGEMA_signal_11370, new_AGEMA_signal_11366, new_AGEMA_signal_11362, new_AGEMA_signal_11358}), .clk ( clk ), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, n2096}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2275 ( .a ({new_AGEMA_signal_11394, new_AGEMA_signal_11388, new_AGEMA_signal_11382, new_AGEMA_signal_11376}), .b ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, n2117}), .clk ( clk ), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, n2128}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2285 ( .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, n2123}), .b ({new_AGEMA_signal_11418, new_AGEMA_signal_11412, new_AGEMA_signal_11406, new_AGEMA_signal_11400}), .clk ( clk ), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2124}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2301 ( .a ({new_AGEMA_signal_11426, new_AGEMA_signal_11424, new_AGEMA_signal_11422, new_AGEMA_signal_11420}), .b ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, n2135}), .clk ( clk ), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, n2148}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2310 ( .a ({new_AGEMA_signal_11450, new_AGEMA_signal_11444, new_AGEMA_signal_11438, new_AGEMA_signal_11432}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, n2141}), .clk ( clk ), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, n2142}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2325 ( .a ({new_AGEMA_signal_11458, new_AGEMA_signal_11456, new_AGEMA_signal_11454, new_AGEMA_signal_11452}), .b ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, n2158}), .clk ( clk ), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, n2168}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2332 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, n2166}), .b ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, n2165}), .clk ( clk ), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, n2167}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2347 ( .a ({new_AGEMA_signal_11474, new_AGEMA_signal_11470, new_AGEMA_signal_11466, new_AGEMA_signal_11462}), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, n2180}), .clk ( clk ), .r ({Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080]}), .c ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2184}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2361 ( .a ({new_AGEMA_signal_11490, new_AGEMA_signal_11486, new_AGEMA_signal_11482, new_AGEMA_signal_11478}), .b ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, n2194}), .clk ( clk ), .r ({Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086]}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, n2197}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2373 ( .a ({new_AGEMA_signal_11498, new_AGEMA_signal_11496, new_AGEMA_signal_11494, new_AGEMA_signal_11492}), .b ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, n2204}), .clk ( clk ), .r ({Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092]}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, n2205}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2390 ( .a ({new_AGEMA_signal_11530, new_AGEMA_signal_11522, new_AGEMA_signal_11514, new_AGEMA_signal_11506}), .b ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, n2225}), .clk ( clk ), .r ({Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098]}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, n2232}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2395 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, n2230}), .b ({new_AGEMA_signal_11554, new_AGEMA_signal_11548, new_AGEMA_signal_11542, new_AGEMA_signal_11536}), .clk ( clk ), .r ({Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104]}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, n2231}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2401 ( .a ({new_AGEMA_signal_11570, new_AGEMA_signal_11566, new_AGEMA_signal_11562, new_AGEMA_signal_11558}), .b ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, n2236}), .clk ( clk ), .r ({Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110]}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, n2239}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2413 ( .a ({new_AGEMA_signal_11586, new_AGEMA_signal_11582, new_AGEMA_signal_11578, new_AGEMA_signal_11574}), .b ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, n2247}), .clk ( clk ), .r ({Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116]}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, n2250}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2428 ( .a ({new_AGEMA_signal_11298, new_AGEMA_signal_11296, new_AGEMA_signal_11294, new_AGEMA_signal_11292}), .b ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, n2264}), .clk ( clk ), .r ({Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122]}), .c ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, n2276}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2439 ( .a ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, n2271}), .b ({new_AGEMA_signal_11594, new_AGEMA_signal_11592, new_AGEMA_signal_11590, new_AGEMA_signal_11588}), .clk ( clk ), .r ({Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128]}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, n2272}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2454 ( .a ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, n2286}), .b ({new_AGEMA_signal_11602, new_AGEMA_signal_11600, new_AGEMA_signal_11598, new_AGEMA_signal_11596}), .clk ( clk ), .r ({Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134]}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, n2306}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2468 ( .a ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, n2295}), .b ({new_AGEMA_signal_11618, new_AGEMA_signal_11614, new_AGEMA_signal_11610, new_AGEMA_signal_11606}), .clk ( clk ), .r ({Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140]}), .c ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2296}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2489 ( .a ({new_AGEMA_signal_11634, new_AGEMA_signal_11630, new_AGEMA_signal_11626, new_AGEMA_signal_11622}), .b ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, n2322}), .clk ( clk ), .r ({Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, n2324}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2500 ( .a ({new_AGEMA_signal_11642, new_AGEMA_signal_11640, new_AGEMA_signal_11638, new_AGEMA_signal_11636}), .b ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, n2333}), .clk ( clk ), .r ({Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152]}), .c ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, n2337}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2511 ( .a ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, n2345}), .b ({new_AGEMA_signal_11666, new_AGEMA_signal_11660, new_AGEMA_signal_11654, new_AGEMA_signal_11648}), .clk ( clk ), .r ({Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158]}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, n2350}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2528 ( .a ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, n2361}), .b ({new_AGEMA_signal_11682, new_AGEMA_signal_11678, new_AGEMA_signal_11674, new_AGEMA_signal_11670}), .clk ( clk ), .r ({Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164]}), .c ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2362}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2550 ( .a ({new_AGEMA_signal_11690, new_AGEMA_signal_11688, new_AGEMA_signal_11686, new_AGEMA_signal_11684}), .b ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, n2388}), .clk ( clk ), .r ({Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170]}), .c ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, n2389}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2557 ( .a ({new_AGEMA_signal_11706, new_AGEMA_signal_11702, new_AGEMA_signal_11698, new_AGEMA_signal_11694}), .b ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, n2393}), .clk ( clk ), .r ({Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176]}), .c ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, n2397}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2568 ( .a ({new_AGEMA_signal_11722, new_AGEMA_signal_11718, new_AGEMA_signal_11714, new_AGEMA_signal_11710}), .b ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, n2405}), .clk ( clk ), .r ({Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182]}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, n2411}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2580 ( .a ({new_AGEMA_signal_11738, new_AGEMA_signal_11734, new_AGEMA_signal_11730, new_AGEMA_signal_11726}), .b ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, n2419}), .clk ( clk ), .r ({Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188]}), .c ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2420}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2593 ( .a ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, n2436}), .b ({new_AGEMA_signal_11746, new_AGEMA_signal_11744, new_AGEMA_signal_11742, new_AGEMA_signal_11740}), .clk ( clk ), .r ({Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, n2440}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2614 ( .a ({new_AGEMA_signal_11762, new_AGEMA_signal_11758, new_AGEMA_signal_11754, new_AGEMA_signal_11750}), .b ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, n2461}), .clk ( clk ), .r ({Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200]}), .c ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, n2516}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2621 ( .s ({new_AGEMA_signal_11770, new_AGEMA_signal_11768, new_AGEMA_signal_11766, new_AGEMA_signal_11764}), .b ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, n2469}), .a ({new_AGEMA_signal_11794, new_AGEMA_signal_11788, new_AGEMA_signal_11782, new_AGEMA_signal_11776}), .clk ( clk ), .r ({Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206]}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, n2471}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2636 ( .a ({new_AGEMA_signal_11818, new_AGEMA_signal_11812, new_AGEMA_signal_11806, new_AGEMA_signal_11800}), .b ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, n2484}), .clk ( clk ), .r ({Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212]}), .c ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2485}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2644 ( .a ({new_AGEMA_signal_11322, new_AGEMA_signal_11316, new_AGEMA_signal_11310, new_AGEMA_signal_11304}), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, n2491}), .clk ( clk ), .r ({Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218]}), .c ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, n2502}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2651 ( .a ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, n2500}), .b ({new_AGEMA_signal_11834, new_AGEMA_signal_11830, new_AGEMA_signal_11826, new_AGEMA_signal_11822}), .clk ( clk ), .r ({Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, n2501}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2657 ( .a ({new_AGEMA_signal_11738, new_AGEMA_signal_11734, new_AGEMA_signal_11730, new_AGEMA_signal_11726}), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, n2508}), .clk ( clk ), .r ({Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230]}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, n2509}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2671 ( .a ({new_AGEMA_signal_11842, new_AGEMA_signal_11840, new_AGEMA_signal_11838, new_AGEMA_signal_11836}), .b ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, n2526}), .clk ( clk ), .r ({Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236]}), .c ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, n2527}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2680 ( .a ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, n2539}), .b ({new_AGEMA_signal_11874, new_AGEMA_signal_11866, new_AGEMA_signal_11858, new_AGEMA_signal_11850}), .clk ( clk ), .r ({Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242]}), .c ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2550}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2685 ( .a ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, n2548}), .b ({new_AGEMA_signal_11882, new_AGEMA_signal_11880, new_AGEMA_signal_11878, new_AGEMA_signal_11876}), .clk ( clk ), .r ({Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, n2549}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2701 ( .a ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, n2568}), .b ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, n2567}), .clk ( clk ), .r ({Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254]}), .c ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, n2569}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2712 ( .a ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, n2583}), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11894, new_AGEMA_signal_11890, new_AGEMA_signal_11886}), .clk ( clk ), .r ({Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, n2584}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2729 ( .a ({new_AGEMA_signal_11914, new_AGEMA_signal_11910, new_AGEMA_signal_11906, new_AGEMA_signal_11902}), .b ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, n2604}), .clk ( clk ), .r ({Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266]}), .c ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n2606}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2740 ( .a ({new_AGEMA_signal_11322, new_AGEMA_signal_11316, new_AGEMA_signal_11310, new_AGEMA_signal_11304}), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, n2621}), .clk ( clk ), .r ({Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, n2622}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2747 ( .a ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, n2633}), .b ({new_AGEMA_signal_11930, new_AGEMA_signal_11926, new_AGEMA_signal_11922, new_AGEMA_signal_11918}), .clk ( clk ), .r ({Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278]}), .c ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, n2634}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2761 ( .a ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, n2656}), .b ({new_AGEMA_signal_11946, new_AGEMA_signal_11942, new_AGEMA_signal_11938, new_AGEMA_signal_11934}), .clk ( clk ), .r ({Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, n2657}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2783 ( .a ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, n2696}), .b ({new_AGEMA_signal_11962, new_AGEMA_signal_11958, new_AGEMA_signal_11954, new_AGEMA_signal_11950}), .clk ( clk ), .r ({Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290]}), .c ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2697}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2795 ( .a ({new_AGEMA_signal_11298, new_AGEMA_signal_11296, new_AGEMA_signal_11294, new_AGEMA_signal_11292}), .b ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, n2718}), .clk ( clk ), .r ({Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, n2808}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2802 ( .a ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, n2730}), .b ({new_AGEMA_signal_11994, new_AGEMA_signal_11986, new_AGEMA_signal_11978, new_AGEMA_signal_11970}), .clk ( clk ), .r ({Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302]}), .c ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, n2747}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2810 ( .a ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, n2745}), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, n2744}), .clk ( clk ), .r ({Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, n2746}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2818 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, n2759}), .b ({new_AGEMA_signal_12002, new_AGEMA_signal_12000, new_AGEMA_signal_11998, new_AGEMA_signal_11996}), .clk ( clk ), .r ({Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314]}), .c ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, n2804}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2824 ( .a ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, n2771}), .b ({new_AGEMA_signal_12018, new_AGEMA_signal_12014, new_AGEMA_signal_12010, new_AGEMA_signal_12006}), .clk ( clk ), .r ({Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, n2802}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2838 ( .a ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, n2798}), .b ({new_AGEMA_signal_12026, new_AGEMA_signal_12024, new_AGEMA_signal_12022, new_AGEMA_signal_12020}), .clk ( clk ), .r ({Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, n2799}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2852 ( .a ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, n2826}), .b ({new_AGEMA_signal_12050, new_AGEMA_signal_12044, new_AGEMA_signal_12038, new_AGEMA_signal_12032}), .clk ( clk ), .r ({Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332]}), .c ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, n2827}) ) ;
    buf_clk new_AGEMA_reg_buffer_4024 ( .C ( clk ), .D ( new_AGEMA_signal_12051 ), .Q ( new_AGEMA_signal_12052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4026 ( .C ( clk ), .D ( new_AGEMA_signal_12053 ), .Q ( new_AGEMA_signal_12054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4028 ( .C ( clk ), .D ( new_AGEMA_signal_12055 ), .Q ( new_AGEMA_signal_12056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4030 ( .C ( clk ), .D ( new_AGEMA_signal_12057 ), .Q ( new_AGEMA_signal_12058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4038 ( .C ( clk ), .D ( new_AGEMA_signal_12065 ), .Q ( new_AGEMA_signal_12066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4046 ( .C ( clk ), .D ( new_AGEMA_signal_12073 ), .Q ( new_AGEMA_signal_12074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4054 ( .C ( clk ), .D ( new_AGEMA_signal_12081 ), .Q ( new_AGEMA_signal_12082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4062 ( .C ( clk ), .D ( new_AGEMA_signal_12089 ), .Q ( new_AGEMA_signal_12090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4064 ( .C ( clk ), .D ( new_AGEMA_signal_12091 ), .Q ( new_AGEMA_signal_12092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4066 ( .C ( clk ), .D ( new_AGEMA_signal_12093 ), .Q ( new_AGEMA_signal_12094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4068 ( .C ( clk ), .D ( new_AGEMA_signal_12095 ), .Q ( new_AGEMA_signal_12096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4070 ( .C ( clk ), .D ( new_AGEMA_signal_12097 ), .Q ( new_AGEMA_signal_12098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4074 ( .C ( clk ), .D ( new_AGEMA_signal_12101 ), .Q ( new_AGEMA_signal_12102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4078 ( .C ( clk ), .D ( new_AGEMA_signal_12105 ), .Q ( new_AGEMA_signal_12106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4082 ( .C ( clk ), .D ( new_AGEMA_signal_12109 ), .Q ( new_AGEMA_signal_12110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4086 ( .C ( clk ), .D ( new_AGEMA_signal_12113 ), .Q ( new_AGEMA_signal_12114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4094 ( .C ( clk ), .D ( new_AGEMA_signal_12121 ), .Q ( new_AGEMA_signal_12122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4102 ( .C ( clk ), .D ( new_AGEMA_signal_12129 ), .Q ( new_AGEMA_signal_12130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4110 ( .C ( clk ), .D ( new_AGEMA_signal_12137 ), .Q ( new_AGEMA_signal_12138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4118 ( .C ( clk ), .D ( new_AGEMA_signal_12145 ), .Q ( new_AGEMA_signal_12146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4120 ( .C ( clk ), .D ( new_AGEMA_signal_12147 ), .Q ( new_AGEMA_signal_12148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4122 ( .C ( clk ), .D ( new_AGEMA_signal_12149 ), .Q ( new_AGEMA_signal_12150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4124 ( .C ( clk ), .D ( new_AGEMA_signal_12151 ), .Q ( new_AGEMA_signal_12152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4126 ( .C ( clk ), .D ( new_AGEMA_signal_12153 ), .Q ( new_AGEMA_signal_12154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4132 ( .C ( clk ), .D ( new_AGEMA_signal_12159 ), .Q ( new_AGEMA_signal_12160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4138 ( .C ( clk ), .D ( new_AGEMA_signal_12165 ), .Q ( new_AGEMA_signal_12166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4144 ( .C ( clk ), .D ( new_AGEMA_signal_12171 ), .Q ( new_AGEMA_signal_12172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4150 ( .C ( clk ), .D ( new_AGEMA_signal_12177 ), .Q ( new_AGEMA_signal_12178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4154 ( .C ( clk ), .D ( new_AGEMA_signal_12181 ), .Q ( new_AGEMA_signal_12182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4158 ( .C ( clk ), .D ( new_AGEMA_signal_12185 ), .Q ( new_AGEMA_signal_12186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4162 ( .C ( clk ), .D ( new_AGEMA_signal_12189 ), .Q ( new_AGEMA_signal_12190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4166 ( .C ( clk ), .D ( new_AGEMA_signal_12193 ), .Q ( new_AGEMA_signal_12194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4174 ( .C ( clk ), .D ( new_AGEMA_signal_12201 ), .Q ( new_AGEMA_signal_12202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4182 ( .C ( clk ), .D ( new_AGEMA_signal_12209 ), .Q ( new_AGEMA_signal_12210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4190 ( .C ( clk ), .D ( new_AGEMA_signal_12217 ), .Q ( new_AGEMA_signal_12218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4198 ( .C ( clk ), .D ( new_AGEMA_signal_12225 ), .Q ( new_AGEMA_signal_12226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4202 ( .C ( clk ), .D ( new_AGEMA_signal_12229 ), .Q ( new_AGEMA_signal_12230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4206 ( .C ( clk ), .D ( new_AGEMA_signal_12233 ), .Q ( new_AGEMA_signal_12234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4210 ( .C ( clk ), .D ( new_AGEMA_signal_12237 ), .Q ( new_AGEMA_signal_12238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4214 ( .C ( clk ), .D ( new_AGEMA_signal_12241 ), .Q ( new_AGEMA_signal_12242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4220 ( .C ( clk ), .D ( new_AGEMA_signal_12247 ), .Q ( new_AGEMA_signal_12248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4226 ( .C ( clk ), .D ( new_AGEMA_signal_12253 ), .Q ( new_AGEMA_signal_12254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4232 ( .C ( clk ), .D ( new_AGEMA_signal_12259 ), .Q ( new_AGEMA_signal_12260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4238 ( .C ( clk ), .D ( new_AGEMA_signal_12265 ), .Q ( new_AGEMA_signal_12266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4244 ( .C ( clk ), .D ( new_AGEMA_signal_12271 ), .Q ( new_AGEMA_signal_12272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4250 ( .C ( clk ), .D ( new_AGEMA_signal_12277 ), .Q ( new_AGEMA_signal_12278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4256 ( .C ( clk ), .D ( new_AGEMA_signal_12283 ), .Q ( new_AGEMA_signal_12284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4262 ( .C ( clk ), .D ( new_AGEMA_signal_12289 ), .Q ( new_AGEMA_signal_12290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4268 ( .C ( clk ), .D ( new_AGEMA_signal_12295 ), .Q ( new_AGEMA_signal_12296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4274 ( .C ( clk ), .D ( new_AGEMA_signal_12301 ), .Q ( new_AGEMA_signal_12302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4280 ( .C ( clk ), .D ( new_AGEMA_signal_12307 ), .Q ( new_AGEMA_signal_12308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4286 ( .C ( clk ), .D ( new_AGEMA_signal_12313 ), .Q ( new_AGEMA_signal_12314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4292 ( .C ( clk ), .D ( new_AGEMA_signal_12319 ), .Q ( new_AGEMA_signal_12320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4298 ( .C ( clk ), .D ( new_AGEMA_signal_12325 ), .Q ( new_AGEMA_signal_12326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4304 ( .C ( clk ), .D ( new_AGEMA_signal_12331 ), .Q ( new_AGEMA_signal_12332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4310 ( .C ( clk ), .D ( new_AGEMA_signal_12337 ), .Q ( new_AGEMA_signal_12338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4316 ( .C ( clk ), .D ( new_AGEMA_signal_12343 ), .Q ( new_AGEMA_signal_12344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4322 ( .C ( clk ), .D ( new_AGEMA_signal_12349 ), .Q ( new_AGEMA_signal_12350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4328 ( .C ( clk ), .D ( new_AGEMA_signal_12355 ), .Q ( new_AGEMA_signal_12356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4334 ( .C ( clk ), .D ( new_AGEMA_signal_12361 ), .Q ( new_AGEMA_signal_12362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4338 ( .C ( clk ), .D ( new_AGEMA_signal_12365 ), .Q ( new_AGEMA_signal_12366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4342 ( .C ( clk ), .D ( new_AGEMA_signal_12369 ), .Q ( new_AGEMA_signal_12370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4346 ( .C ( clk ), .D ( new_AGEMA_signal_12373 ), .Q ( new_AGEMA_signal_12374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4350 ( .C ( clk ), .D ( new_AGEMA_signal_12377 ), .Q ( new_AGEMA_signal_12378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4358 ( .C ( clk ), .D ( new_AGEMA_signal_12385 ), .Q ( new_AGEMA_signal_12386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4366 ( .C ( clk ), .D ( new_AGEMA_signal_12393 ), .Q ( new_AGEMA_signal_12394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4374 ( .C ( clk ), .D ( new_AGEMA_signal_12401 ), .Q ( new_AGEMA_signal_12402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4382 ( .C ( clk ), .D ( new_AGEMA_signal_12409 ), .Q ( new_AGEMA_signal_12410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4386 ( .C ( clk ), .D ( new_AGEMA_signal_12413 ), .Q ( new_AGEMA_signal_12414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4390 ( .C ( clk ), .D ( new_AGEMA_signal_12417 ), .Q ( new_AGEMA_signal_12418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4394 ( .C ( clk ), .D ( new_AGEMA_signal_12421 ), .Q ( new_AGEMA_signal_12422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4398 ( .C ( clk ), .D ( new_AGEMA_signal_12425 ), .Q ( new_AGEMA_signal_12426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4404 ( .C ( clk ), .D ( new_AGEMA_signal_12431 ), .Q ( new_AGEMA_signal_12432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4410 ( .C ( clk ), .D ( new_AGEMA_signal_12437 ), .Q ( new_AGEMA_signal_12438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4416 ( .C ( clk ), .D ( new_AGEMA_signal_12443 ), .Q ( new_AGEMA_signal_12444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4422 ( .C ( clk ), .D ( new_AGEMA_signal_12449 ), .Q ( new_AGEMA_signal_12450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4430 ( .C ( clk ), .D ( new_AGEMA_signal_12457 ), .Q ( new_AGEMA_signal_12458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4438 ( .C ( clk ), .D ( new_AGEMA_signal_12465 ), .Q ( new_AGEMA_signal_12466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4446 ( .C ( clk ), .D ( new_AGEMA_signal_12473 ), .Q ( new_AGEMA_signal_12474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4454 ( .C ( clk ), .D ( new_AGEMA_signal_12481 ), .Q ( new_AGEMA_signal_12482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4456 ( .C ( clk ), .D ( new_AGEMA_signal_12483 ), .Q ( new_AGEMA_signal_12484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4458 ( .C ( clk ), .D ( new_AGEMA_signal_12485 ), .Q ( new_AGEMA_signal_12486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4460 ( .C ( clk ), .D ( new_AGEMA_signal_12487 ), .Q ( new_AGEMA_signal_12488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4462 ( .C ( clk ), .D ( new_AGEMA_signal_12489 ), .Q ( new_AGEMA_signal_12490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4468 ( .C ( clk ), .D ( new_AGEMA_signal_12495 ), .Q ( new_AGEMA_signal_12496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4474 ( .C ( clk ), .D ( new_AGEMA_signal_12501 ), .Q ( new_AGEMA_signal_12502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4480 ( .C ( clk ), .D ( new_AGEMA_signal_12507 ), .Q ( new_AGEMA_signal_12508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4486 ( .C ( clk ), .D ( new_AGEMA_signal_12513 ), .Q ( new_AGEMA_signal_12514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4488 ( .C ( clk ), .D ( new_AGEMA_signal_12515 ), .Q ( new_AGEMA_signal_12516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4490 ( .C ( clk ), .D ( new_AGEMA_signal_12517 ), .Q ( new_AGEMA_signal_12518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4492 ( .C ( clk ), .D ( new_AGEMA_signal_12519 ), .Q ( new_AGEMA_signal_12520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4494 ( .C ( clk ), .D ( new_AGEMA_signal_12521 ), .Q ( new_AGEMA_signal_12522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4496 ( .C ( clk ), .D ( new_AGEMA_signal_12523 ), .Q ( new_AGEMA_signal_12524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4498 ( .C ( clk ), .D ( new_AGEMA_signal_12525 ), .Q ( new_AGEMA_signal_12526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4500 ( .C ( clk ), .D ( new_AGEMA_signal_12527 ), .Q ( new_AGEMA_signal_12528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4502 ( .C ( clk ), .D ( new_AGEMA_signal_12529 ), .Q ( new_AGEMA_signal_12530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4508 ( .C ( clk ), .D ( new_AGEMA_signal_12535 ), .Q ( new_AGEMA_signal_12536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4514 ( .C ( clk ), .D ( new_AGEMA_signal_12541 ), .Q ( new_AGEMA_signal_12542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4520 ( .C ( clk ), .D ( new_AGEMA_signal_12547 ), .Q ( new_AGEMA_signal_12548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4526 ( .C ( clk ), .D ( new_AGEMA_signal_12553 ), .Q ( new_AGEMA_signal_12554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4532 ( .C ( clk ), .D ( new_AGEMA_signal_12559 ), .Q ( new_AGEMA_signal_12560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4538 ( .C ( clk ), .D ( new_AGEMA_signal_12565 ), .Q ( new_AGEMA_signal_12566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4544 ( .C ( clk ), .D ( new_AGEMA_signal_12571 ), .Q ( new_AGEMA_signal_12572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4550 ( .C ( clk ), .D ( new_AGEMA_signal_12577 ), .Q ( new_AGEMA_signal_12578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4558 ( .C ( clk ), .D ( new_AGEMA_signal_12585 ), .Q ( new_AGEMA_signal_12586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4566 ( .C ( clk ), .D ( new_AGEMA_signal_12593 ), .Q ( new_AGEMA_signal_12594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4574 ( .C ( clk ), .D ( new_AGEMA_signal_12601 ), .Q ( new_AGEMA_signal_12602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4582 ( .C ( clk ), .D ( new_AGEMA_signal_12609 ), .Q ( new_AGEMA_signal_12610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4590 ( .C ( clk ), .D ( new_AGEMA_signal_12617 ), .Q ( new_AGEMA_signal_12618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4598 ( .C ( clk ), .D ( new_AGEMA_signal_12625 ), .Q ( new_AGEMA_signal_12626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4606 ( .C ( clk ), .D ( new_AGEMA_signal_12633 ), .Q ( new_AGEMA_signal_12634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4614 ( .C ( clk ), .D ( new_AGEMA_signal_12641 ), .Q ( new_AGEMA_signal_12642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4620 ( .C ( clk ), .D ( new_AGEMA_signal_12647 ), .Q ( new_AGEMA_signal_12648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4626 ( .C ( clk ), .D ( new_AGEMA_signal_12653 ), .Q ( new_AGEMA_signal_12654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4632 ( .C ( clk ), .D ( new_AGEMA_signal_12659 ), .Q ( new_AGEMA_signal_12660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4638 ( .C ( clk ), .D ( new_AGEMA_signal_12665 ), .Q ( new_AGEMA_signal_12666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4644 ( .C ( clk ), .D ( new_AGEMA_signal_12671 ), .Q ( new_AGEMA_signal_12672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4650 ( .C ( clk ), .D ( new_AGEMA_signal_12677 ), .Q ( new_AGEMA_signal_12678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4656 ( .C ( clk ), .D ( new_AGEMA_signal_12683 ), .Q ( new_AGEMA_signal_12684 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4662 ( .C ( clk ), .D ( new_AGEMA_signal_12689 ), .Q ( new_AGEMA_signal_12690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4664 ( .C ( clk ), .D ( new_AGEMA_signal_12691 ), .Q ( new_AGEMA_signal_12692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4666 ( .C ( clk ), .D ( new_AGEMA_signal_12693 ), .Q ( new_AGEMA_signal_12694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4668 ( .C ( clk ), .D ( new_AGEMA_signal_12695 ), .Q ( new_AGEMA_signal_12696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4670 ( .C ( clk ), .D ( new_AGEMA_signal_12697 ), .Q ( new_AGEMA_signal_12698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4674 ( .C ( clk ), .D ( new_AGEMA_signal_12701 ), .Q ( new_AGEMA_signal_12702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4678 ( .C ( clk ), .D ( new_AGEMA_signal_12705 ), .Q ( new_AGEMA_signal_12706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4682 ( .C ( clk ), .D ( new_AGEMA_signal_12709 ), .Q ( new_AGEMA_signal_12710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4686 ( .C ( clk ), .D ( new_AGEMA_signal_12713 ), .Q ( new_AGEMA_signal_12714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4690 ( .C ( clk ), .D ( new_AGEMA_signal_12717 ), .Q ( new_AGEMA_signal_12718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4694 ( .C ( clk ), .D ( new_AGEMA_signal_12721 ), .Q ( new_AGEMA_signal_12722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4698 ( .C ( clk ), .D ( new_AGEMA_signal_12725 ), .Q ( new_AGEMA_signal_12726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4702 ( .C ( clk ), .D ( new_AGEMA_signal_12729 ), .Q ( new_AGEMA_signal_12730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4706 ( .C ( clk ), .D ( new_AGEMA_signal_12733 ), .Q ( new_AGEMA_signal_12734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4710 ( .C ( clk ), .D ( new_AGEMA_signal_12737 ), .Q ( new_AGEMA_signal_12738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4714 ( .C ( clk ), .D ( new_AGEMA_signal_12741 ), .Q ( new_AGEMA_signal_12742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4718 ( .C ( clk ), .D ( new_AGEMA_signal_12745 ), .Q ( new_AGEMA_signal_12746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4720 ( .C ( clk ), .D ( new_AGEMA_signal_12747 ), .Q ( new_AGEMA_signal_12748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4722 ( .C ( clk ), .D ( new_AGEMA_signal_12749 ), .Q ( new_AGEMA_signal_12750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4724 ( .C ( clk ), .D ( new_AGEMA_signal_12751 ), .Q ( new_AGEMA_signal_12752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4726 ( .C ( clk ), .D ( new_AGEMA_signal_12753 ), .Q ( new_AGEMA_signal_12754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4730 ( .C ( clk ), .D ( new_AGEMA_signal_12757 ), .Q ( new_AGEMA_signal_12758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4736 ( .C ( clk ), .D ( new_AGEMA_signal_12763 ), .Q ( new_AGEMA_signal_12764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4742 ( .C ( clk ), .D ( new_AGEMA_signal_12769 ), .Q ( new_AGEMA_signal_12770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4748 ( .C ( clk ), .D ( new_AGEMA_signal_12775 ), .Q ( new_AGEMA_signal_12776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4760 ( .C ( clk ), .D ( new_AGEMA_signal_12787 ), .Q ( new_AGEMA_signal_12788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4764 ( .C ( clk ), .D ( new_AGEMA_signal_12791 ), .Q ( new_AGEMA_signal_12792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4768 ( .C ( clk ), .D ( new_AGEMA_signal_12795 ), .Q ( new_AGEMA_signal_12796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4772 ( .C ( clk ), .D ( new_AGEMA_signal_12799 ), .Q ( new_AGEMA_signal_12800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4780 ( .C ( clk ), .D ( new_AGEMA_signal_12807 ), .Q ( new_AGEMA_signal_12808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4788 ( .C ( clk ), .D ( new_AGEMA_signal_12815 ), .Q ( new_AGEMA_signal_12816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4796 ( .C ( clk ), .D ( new_AGEMA_signal_12823 ), .Q ( new_AGEMA_signal_12824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4804 ( .C ( clk ), .D ( new_AGEMA_signal_12831 ), .Q ( new_AGEMA_signal_12832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4812 ( .C ( clk ), .D ( new_AGEMA_signal_12839 ), .Q ( new_AGEMA_signal_12840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4820 ( .C ( clk ), .D ( new_AGEMA_signal_12847 ), .Q ( new_AGEMA_signal_12848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4828 ( .C ( clk ), .D ( new_AGEMA_signal_12855 ), .Q ( new_AGEMA_signal_12856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4836 ( .C ( clk ), .D ( new_AGEMA_signal_12863 ), .Q ( new_AGEMA_signal_12864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4844 ( .C ( clk ), .D ( new_AGEMA_signal_12871 ), .Q ( new_AGEMA_signal_12872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4852 ( .C ( clk ), .D ( new_AGEMA_signal_12879 ), .Q ( new_AGEMA_signal_12880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4860 ( .C ( clk ), .D ( new_AGEMA_signal_12887 ), .Q ( new_AGEMA_signal_12888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4868 ( .C ( clk ), .D ( new_AGEMA_signal_12895 ), .Q ( new_AGEMA_signal_12896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4876 ( .C ( clk ), .D ( new_AGEMA_signal_12903 ), .Q ( new_AGEMA_signal_12904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4884 ( .C ( clk ), .D ( new_AGEMA_signal_12911 ), .Q ( new_AGEMA_signal_12912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4892 ( .C ( clk ), .D ( new_AGEMA_signal_12919 ), .Q ( new_AGEMA_signal_12920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4900 ( .C ( clk ), .D ( new_AGEMA_signal_12927 ), .Q ( new_AGEMA_signal_12928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4906 ( .C ( clk ), .D ( new_AGEMA_signal_12933 ), .Q ( new_AGEMA_signal_12934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4912 ( .C ( clk ), .D ( new_AGEMA_signal_12939 ), .Q ( new_AGEMA_signal_12940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4918 ( .C ( clk ), .D ( new_AGEMA_signal_12945 ), .Q ( new_AGEMA_signal_12946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4924 ( .C ( clk ), .D ( new_AGEMA_signal_12951 ), .Q ( new_AGEMA_signal_12952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4934 ( .C ( clk ), .D ( new_AGEMA_signal_12961 ), .Q ( new_AGEMA_signal_12962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4944 ( .C ( clk ), .D ( new_AGEMA_signal_12971 ), .Q ( new_AGEMA_signal_12972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4954 ( .C ( clk ), .D ( new_AGEMA_signal_12981 ), .Q ( new_AGEMA_signal_12982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4964 ( .C ( clk ), .D ( new_AGEMA_signal_12991 ), .Q ( new_AGEMA_signal_12992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4972 ( .C ( clk ), .D ( new_AGEMA_signal_12999 ), .Q ( new_AGEMA_signal_13000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4980 ( .C ( clk ), .D ( new_AGEMA_signal_13007 ), .Q ( new_AGEMA_signal_13008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4988 ( .C ( clk ), .D ( new_AGEMA_signal_13015 ), .Q ( new_AGEMA_signal_13016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4996 ( .C ( clk ), .D ( new_AGEMA_signal_13023 ), .Q ( new_AGEMA_signal_13024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5004 ( .C ( clk ), .D ( new_AGEMA_signal_13031 ), .Q ( new_AGEMA_signal_13032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5012 ( .C ( clk ), .D ( new_AGEMA_signal_13039 ), .Q ( new_AGEMA_signal_13040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5020 ( .C ( clk ), .D ( new_AGEMA_signal_13047 ), .Q ( new_AGEMA_signal_13048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5028 ( .C ( clk ), .D ( new_AGEMA_signal_13055 ), .Q ( new_AGEMA_signal_13056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5036 ( .C ( clk ), .D ( new_AGEMA_signal_13063 ), .Q ( new_AGEMA_signal_13064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5044 ( .C ( clk ), .D ( new_AGEMA_signal_13071 ), .Q ( new_AGEMA_signal_13072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5052 ( .C ( clk ), .D ( new_AGEMA_signal_13079 ), .Q ( new_AGEMA_signal_13080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5060 ( .C ( clk ), .D ( new_AGEMA_signal_13087 ), .Q ( new_AGEMA_signal_13088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5072 ( .C ( clk ), .D ( new_AGEMA_signal_13099 ), .Q ( new_AGEMA_signal_13100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5076 ( .C ( clk ), .D ( new_AGEMA_signal_13103 ), .Q ( new_AGEMA_signal_13104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5080 ( .C ( clk ), .D ( new_AGEMA_signal_13107 ), .Q ( new_AGEMA_signal_13108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5084 ( .C ( clk ), .D ( new_AGEMA_signal_13111 ), .Q ( new_AGEMA_signal_13112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5090 ( .C ( clk ), .D ( new_AGEMA_signal_13117 ), .Q ( new_AGEMA_signal_13118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5096 ( .C ( clk ), .D ( new_AGEMA_signal_13123 ), .Q ( new_AGEMA_signal_13124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5102 ( .C ( clk ), .D ( new_AGEMA_signal_13129 ), .Q ( new_AGEMA_signal_13130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5108 ( .C ( clk ), .D ( new_AGEMA_signal_13135 ), .Q ( new_AGEMA_signal_13136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5112 ( .C ( clk ), .D ( new_AGEMA_signal_13139 ), .Q ( new_AGEMA_signal_13140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5116 ( .C ( clk ), .D ( new_AGEMA_signal_13143 ), .Q ( new_AGEMA_signal_13144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5120 ( .C ( clk ), .D ( new_AGEMA_signal_13147 ), .Q ( new_AGEMA_signal_13148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5124 ( .C ( clk ), .D ( new_AGEMA_signal_13151 ), .Q ( new_AGEMA_signal_13152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5134 ( .C ( clk ), .D ( new_AGEMA_signal_13161 ), .Q ( new_AGEMA_signal_13162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5144 ( .C ( clk ), .D ( new_AGEMA_signal_13171 ), .Q ( new_AGEMA_signal_13172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5154 ( .C ( clk ), .D ( new_AGEMA_signal_13181 ), .Q ( new_AGEMA_signal_13182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5164 ( .C ( clk ), .D ( new_AGEMA_signal_13191 ), .Q ( new_AGEMA_signal_13192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5172 ( .C ( clk ), .D ( new_AGEMA_signal_13199 ), .Q ( new_AGEMA_signal_13200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5180 ( .C ( clk ), .D ( new_AGEMA_signal_13207 ), .Q ( new_AGEMA_signal_13208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5188 ( .C ( clk ), .D ( new_AGEMA_signal_13215 ), .Q ( new_AGEMA_signal_13216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C ( clk ), .D ( new_AGEMA_signal_13223 ), .Q ( new_AGEMA_signal_13224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C ( clk ), .D ( new_AGEMA_signal_13227 ), .Q ( new_AGEMA_signal_13228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C ( clk ), .D ( new_AGEMA_signal_13231 ), .Q ( new_AGEMA_signal_13232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C ( clk ), .D ( new_AGEMA_signal_13235 ), .Q ( new_AGEMA_signal_13236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C ( clk ), .D ( new_AGEMA_signal_13239 ), .Q ( new_AGEMA_signal_13240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C ( clk ), .D ( new_AGEMA_signal_13255 ), .Q ( new_AGEMA_signal_13256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C ( clk ), .D ( new_AGEMA_signal_13263 ), .Q ( new_AGEMA_signal_13264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C ( clk ), .D ( new_AGEMA_signal_13271 ), .Q ( new_AGEMA_signal_13272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C ( clk ), .D ( new_AGEMA_signal_13279 ), .Q ( new_AGEMA_signal_13280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5260 ( .C ( clk ), .D ( new_AGEMA_signal_13287 ), .Q ( new_AGEMA_signal_13288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5268 ( .C ( clk ), .D ( new_AGEMA_signal_13295 ), .Q ( new_AGEMA_signal_13296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5276 ( .C ( clk ), .D ( new_AGEMA_signal_13303 ), .Q ( new_AGEMA_signal_13304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5284 ( .C ( clk ), .D ( new_AGEMA_signal_13311 ), .Q ( new_AGEMA_signal_13312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5290 ( .C ( clk ), .D ( new_AGEMA_signal_13317 ), .Q ( new_AGEMA_signal_13318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5296 ( .C ( clk ), .D ( new_AGEMA_signal_13323 ), .Q ( new_AGEMA_signal_13324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5302 ( .C ( clk ), .D ( new_AGEMA_signal_13329 ), .Q ( new_AGEMA_signal_13330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5308 ( .C ( clk ), .D ( new_AGEMA_signal_13335 ), .Q ( new_AGEMA_signal_13336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5312 ( .C ( clk ), .D ( new_AGEMA_signal_13339 ), .Q ( new_AGEMA_signal_13340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5316 ( .C ( clk ), .D ( new_AGEMA_signal_13343 ), .Q ( new_AGEMA_signal_13344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5320 ( .C ( clk ), .D ( new_AGEMA_signal_13347 ), .Q ( new_AGEMA_signal_13348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5324 ( .C ( clk ), .D ( new_AGEMA_signal_13351 ), .Q ( new_AGEMA_signal_13352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5332 ( .C ( clk ), .D ( new_AGEMA_signal_13359 ), .Q ( new_AGEMA_signal_13360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5340 ( .C ( clk ), .D ( new_AGEMA_signal_13367 ), .Q ( new_AGEMA_signal_13368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5348 ( .C ( clk ), .D ( new_AGEMA_signal_13375 ), .Q ( new_AGEMA_signal_13376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5356 ( .C ( clk ), .D ( new_AGEMA_signal_13383 ), .Q ( new_AGEMA_signal_13384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5368 ( .C ( clk ), .D ( new_AGEMA_signal_13395 ), .Q ( new_AGEMA_signal_13396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5374 ( .C ( clk ), .D ( new_AGEMA_signal_13401 ), .Q ( new_AGEMA_signal_13402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5380 ( .C ( clk ), .D ( new_AGEMA_signal_13407 ), .Q ( new_AGEMA_signal_13408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5386 ( .C ( clk ), .D ( new_AGEMA_signal_13413 ), .Q ( new_AGEMA_signal_13414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5392 ( .C ( clk ), .D ( new_AGEMA_signal_13419 ), .Q ( new_AGEMA_signal_13420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5398 ( .C ( clk ), .D ( new_AGEMA_signal_13425 ), .Q ( new_AGEMA_signal_13426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5404 ( .C ( clk ), .D ( new_AGEMA_signal_13431 ), .Q ( new_AGEMA_signal_13432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5410 ( .C ( clk ), .D ( new_AGEMA_signal_13437 ), .Q ( new_AGEMA_signal_13438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5416 ( .C ( clk ), .D ( new_AGEMA_signal_13443 ), .Q ( new_AGEMA_signal_13444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5422 ( .C ( clk ), .D ( new_AGEMA_signal_13449 ), .Q ( new_AGEMA_signal_13450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5428 ( .C ( clk ), .D ( new_AGEMA_signal_13455 ), .Q ( new_AGEMA_signal_13456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5434 ( .C ( clk ), .D ( new_AGEMA_signal_13461 ), .Q ( new_AGEMA_signal_13462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5458 ( .C ( clk ), .D ( new_AGEMA_signal_13485 ), .Q ( new_AGEMA_signal_13486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5466 ( .C ( clk ), .D ( new_AGEMA_signal_13493 ), .Q ( new_AGEMA_signal_13494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5474 ( .C ( clk ), .D ( new_AGEMA_signal_13501 ), .Q ( new_AGEMA_signal_13502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5482 ( .C ( clk ), .D ( new_AGEMA_signal_13509 ), .Q ( new_AGEMA_signal_13510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5488 ( .C ( clk ), .D ( new_AGEMA_signal_13515 ), .Q ( new_AGEMA_signal_13516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5494 ( .C ( clk ), .D ( new_AGEMA_signal_13521 ), .Q ( new_AGEMA_signal_13522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5500 ( .C ( clk ), .D ( new_AGEMA_signal_13527 ), .Q ( new_AGEMA_signal_13528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5506 ( .C ( clk ), .D ( new_AGEMA_signal_13533 ), .Q ( new_AGEMA_signal_13534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5530 ( .C ( clk ), .D ( new_AGEMA_signal_13557 ), .Q ( new_AGEMA_signal_13558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5538 ( .C ( clk ), .D ( new_AGEMA_signal_13565 ), .Q ( new_AGEMA_signal_13566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5546 ( .C ( clk ), .D ( new_AGEMA_signal_13573 ), .Q ( new_AGEMA_signal_13574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5554 ( .C ( clk ), .D ( new_AGEMA_signal_13581 ), .Q ( new_AGEMA_signal_13582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5562 ( .C ( clk ), .D ( new_AGEMA_signal_13589 ), .Q ( new_AGEMA_signal_13590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5570 ( .C ( clk ), .D ( new_AGEMA_signal_13597 ), .Q ( new_AGEMA_signal_13598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5578 ( .C ( clk ), .D ( new_AGEMA_signal_13605 ), .Q ( new_AGEMA_signal_13606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5586 ( .C ( clk ), .D ( new_AGEMA_signal_13613 ), .Q ( new_AGEMA_signal_13614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5596 ( .C ( clk ), .D ( new_AGEMA_signal_13623 ), .Q ( new_AGEMA_signal_13624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5606 ( .C ( clk ), .D ( new_AGEMA_signal_13633 ), .Q ( new_AGEMA_signal_13634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5616 ( .C ( clk ), .D ( new_AGEMA_signal_13643 ), .Q ( new_AGEMA_signal_13644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5626 ( .C ( clk ), .D ( new_AGEMA_signal_13653 ), .Q ( new_AGEMA_signal_13654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5634 ( .C ( clk ), .D ( new_AGEMA_signal_13661 ), .Q ( new_AGEMA_signal_13662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5642 ( .C ( clk ), .D ( new_AGEMA_signal_13669 ), .Q ( new_AGEMA_signal_13670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5650 ( .C ( clk ), .D ( new_AGEMA_signal_13677 ), .Q ( new_AGEMA_signal_13678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5658 ( .C ( clk ), .D ( new_AGEMA_signal_13685 ), .Q ( new_AGEMA_signal_13686 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5664 ( .C ( clk ), .D ( new_AGEMA_signal_13691 ), .Q ( new_AGEMA_signal_13692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5670 ( .C ( clk ), .D ( new_AGEMA_signal_13697 ), .Q ( new_AGEMA_signal_13698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5676 ( .C ( clk ), .D ( new_AGEMA_signal_13703 ), .Q ( new_AGEMA_signal_13704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5682 ( .C ( clk ), .D ( new_AGEMA_signal_13709 ), .Q ( new_AGEMA_signal_13710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5704 ( .C ( clk ), .D ( new_AGEMA_signal_13731 ), .Q ( new_AGEMA_signal_13732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5710 ( .C ( clk ), .D ( new_AGEMA_signal_13737 ), .Q ( new_AGEMA_signal_13738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5716 ( .C ( clk ), .D ( new_AGEMA_signal_13743 ), .Q ( new_AGEMA_signal_13744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5722 ( .C ( clk ), .D ( new_AGEMA_signal_13749 ), .Q ( new_AGEMA_signal_13750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5730 ( .C ( clk ), .D ( new_AGEMA_signal_13757 ), .Q ( new_AGEMA_signal_13758 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5738 ( .C ( clk ), .D ( new_AGEMA_signal_13765 ), .Q ( new_AGEMA_signal_13766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5746 ( .C ( clk ), .D ( new_AGEMA_signal_13773 ), .Q ( new_AGEMA_signal_13774 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5754 ( .C ( clk ), .D ( new_AGEMA_signal_13781 ), .Q ( new_AGEMA_signal_13782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5760 ( .C ( clk ), .D ( new_AGEMA_signal_13787 ), .Q ( new_AGEMA_signal_13788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5766 ( .C ( clk ), .D ( new_AGEMA_signal_13793 ), .Q ( new_AGEMA_signal_13794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5772 ( .C ( clk ), .D ( new_AGEMA_signal_13799 ), .Q ( new_AGEMA_signal_13800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5778 ( .C ( clk ), .D ( new_AGEMA_signal_13805 ), .Q ( new_AGEMA_signal_13806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5794 ( .C ( clk ), .D ( new_AGEMA_signal_13821 ), .Q ( new_AGEMA_signal_13822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5802 ( .C ( clk ), .D ( new_AGEMA_signal_13829 ), .Q ( new_AGEMA_signal_13830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5810 ( .C ( clk ), .D ( new_AGEMA_signal_13837 ), .Q ( new_AGEMA_signal_13838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5818 ( .C ( clk ), .D ( new_AGEMA_signal_13845 ), .Q ( new_AGEMA_signal_13846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5840 ( .C ( clk ), .D ( new_AGEMA_signal_13867 ), .Q ( new_AGEMA_signal_13868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5846 ( .C ( clk ), .D ( new_AGEMA_signal_13873 ), .Q ( new_AGEMA_signal_13874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5852 ( .C ( clk ), .D ( new_AGEMA_signal_13879 ), .Q ( new_AGEMA_signal_13880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5858 ( .C ( clk ), .D ( new_AGEMA_signal_13885 ), .Q ( new_AGEMA_signal_13886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5864 ( .C ( clk ), .D ( new_AGEMA_signal_13891 ), .Q ( new_AGEMA_signal_13892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5870 ( .C ( clk ), .D ( new_AGEMA_signal_13897 ), .Q ( new_AGEMA_signal_13898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5876 ( .C ( clk ), .D ( new_AGEMA_signal_13903 ), .Q ( new_AGEMA_signal_13904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5882 ( .C ( clk ), .D ( new_AGEMA_signal_13909 ), .Q ( new_AGEMA_signal_13910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5970 ( .C ( clk ), .D ( new_AGEMA_signal_13997 ), .Q ( new_AGEMA_signal_13998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5980 ( .C ( clk ), .D ( new_AGEMA_signal_14007 ), .Q ( new_AGEMA_signal_14008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5990 ( .C ( clk ), .D ( new_AGEMA_signal_14017 ), .Q ( new_AGEMA_signal_14018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6000 ( .C ( clk ), .D ( new_AGEMA_signal_14027 ), .Q ( new_AGEMA_signal_14028 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6088 ( .C ( clk ), .D ( new_AGEMA_signal_14115 ), .Q ( new_AGEMA_signal_14116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6096 ( .C ( clk ), .D ( new_AGEMA_signal_14123 ), .Q ( new_AGEMA_signal_14124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6104 ( .C ( clk ), .D ( new_AGEMA_signal_14131 ), .Q ( new_AGEMA_signal_14132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6112 ( .C ( clk ), .D ( new_AGEMA_signal_14139 ), .Q ( new_AGEMA_signal_14140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6144 ( .C ( clk ), .D ( new_AGEMA_signal_14171 ), .Q ( new_AGEMA_signal_14172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6152 ( .C ( clk ), .D ( new_AGEMA_signal_14179 ), .Q ( new_AGEMA_signal_14180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6160 ( .C ( clk ), .D ( new_AGEMA_signal_14187 ), .Q ( new_AGEMA_signal_14188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6168 ( .C ( clk ), .D ( new_AGEMA_signal_14195 ), .Q ( new_AGEMA_signal_14196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6176 ( .C ( clk ), .D ( new_AGEMA_signal_14203 ), .Q ( new_AGEMA_signal_14204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6184 ( .C ( clk ), .D ( new_AGEMA_signal_14211 ), .Q ( new_AGEMA_signal_14212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6192 ( .C ( clk ), .D ( new_AGEMA_signal_14219 ), .Q ( new_AGEMA_signal_14220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6200 ( .C ( clk ), .D ( new_AGEMA_signal_14227 ), .Q ( new_AGEMA_signal_14228 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6248 ( .C ( clk ), .D ( new_AGEMA_signal_14275 ), .Q ( new_AGEMA_signal_14276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6256 ( .C ( clk ), .D ( new_AGEMA_signal_14283 ), .Q ( new_AGEMA_signal_14284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6264 ( .C ( clk ), .D ( new_AGEMA_signal_14291 ), .Q ( new_AGEMA_signal_14292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6272 ( .C ( clk ), .D ( new_AGEMA_signal_14299 ), .Q ( new_AGEMA_signal_14300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6330 ( .C ( clk ), .D ( new_AGEMA_signal_14357 ), .Q ( new_AGEMA_signal_14358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6342 ( .C ( clk ), .D ( new_AGEMA_signal_14369 ), .Q ( new_AGEMA_signal_14370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6354 ( .C ( clk ), .D ( new_AGEMA_signal_14381 ), .Q ( new_AGEMA_signal_14382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6366 ( .C ( clk ), .D ( new_AGEMA_signal_14393 ), .Q ( new_AGEMA_signal_14394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6380 ( .C ( clk ), .D ( new_AGEMA_signal_14407 ), .Q ( new_AGEMA_signal_14408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6394 ( .C ( clk ), .D ( new_AGEMA_signal_14421 ), .Q ( new_AGEMA_signal_14422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6408 ( .C ( clk ), .D ( new_AGEMA_signal_14435 ), .Q ( new_AGEMA_signal_14436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6422 ( .C ( clk ), .D ( new_AGEMA_signal_14449 ), .Q ( new_AGEMA_signal_14450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6468 ( .C ( clk ), .D ( new_AGEMA_signal_14495 ), .Q ( new_AGEMA_signal_14496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6482 ( .C ( clk ), .D ( new_AGEMA_signal_14509 ), .Q ( new_AGEMA_signal_14510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6496 ( .C ( clk ), .D ( new_AGEMA_signal_14523 ), .Q ( new_AGEMA_signal_14524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6510 ( .C ( clk ), .D ( new_AGEMA_signal_14537 ), .Q ( new_AGEMA_signal_14538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6612 ( .C ( clk ), .D ( new_AGEMA_signal_14639 ), .Q ( new_AGEMA_signal_14640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6628 ( .C ( clk ), .D ( new_AGEMA_signal_14655 ), .Q ( new_AGEMA_signal_14656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6644 ( .C ( clk ), .D ( new_AGEMA_signal_14671 ), .Q ( new_AGEMA_signal_14672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6660 ( .C ( clk ), .D ( new_AGEMA_signal_14687 ), .Q ( new_AGEMA_signal_14688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6700 ( .C ( clk ), .D ( new_AGEMA_signal_14727 ), .Q ( new_AGEMA_signal_14728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6716 ( .C ( clk ), .D ( new_AGEMA_signal_14743 ), .Q ( new_AGEMA_signal_14744 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6732 ( .C ( clk ), .D ( new_AGEMA_signal_14759 ), .Q ( new_AGEMA_signal_14760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6748 ( .C ( clk ), .D ( new_AGEMA_signal_14775 ), .Q ( new_AGEMA_signal_14776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6898 ( .C ( clk ), .D ( new_AGEMA_signal_14925 ), .Q ( new_AGEMA_signal_14926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6914 ( .C ( clk ), .D ( new_AGEMA_signal_14941 ), .Q ( new_AGEMA_signal_14942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6930 ( .C ( clk ), .D ( new_AGEMA_signal_14957 ), .Q ( new_AGEMA_signal_14958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6946 ( .C ( clk ), .D ( new_AGEMA_signal_14973 ), .Q ( new_AGEMA_signal_14974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7004 ( .C ( clk ), .D ( new_AGEMA_signal_15031 ), .Q ( new_AGEMA_signal_15032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7022 ( .C ( clk ), .D ( new_AGEMA_signal_15049 ), .Q ( new_AGEMA_signal_15050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7040 ( .C ( clk ), .D ( new_AGEMA_signal_15067 ), .Q ( new_AGEMA_signal_15068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7058 ( .C ( clk ), .D ( new_AGEMA_signal_15085 ), .Q ( new_AGEMA_signal_15086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7204 ( .C ( clk ), .D ( new_AGEMA_signal_15231 ), .Q ( new_AGEMA_signal_15232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7224 ( .C ( clk ), .D ( new_AGEMA_signal_15251 ), .Q ( new_AGEMA_signal_15252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7244 ( .C ( clk ), .D ( new_AGEMA_signal_15271 ), .Q ( new_AGEMA_signal_15272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7264 ( .C ( clk ), .D ( new_AGEMA_signal_15291 ), .Q ( new_AGEMA_signal_15292 ) ) ;

    /* cells in depth 13 */
    buf_clk new_AGEMA_reg_buffer_4731 ( .C ( clk ), .D ( new_AGEMA_signal_12758 ), .Q ( new_AGEMA_signal_12759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4737 ( .C ( clk ), .D ( new_AGEMA_signal_12764 ), .Q ( new_AGEMA_signal_12765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4743 ( .C ( clk ), .D ( new_AGEMA_signal_12770 ), .Q ( new_AGEMA_signal_12771 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4749 ( .C ( clk ), .D ( new_AGEMA_signal_12776 ), .Q ( new_AGEMA_signal_12777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4751 ( .C ( clk ), .D ( new_AGEMA_signal_12702 ), .Q ( new_AGEMA_signal_12779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4753 ( .C ( clk ), .D ( new_AGEMA_signal_12706 ), .Q ( new_AGEMA_signal_12781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4755 ( .C ( clk ), .D ( new_AGEMA_signal_12710 ), .Q ( new_AGEMA_signal_12783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4757 ( .C ( clk ), .D ( new_AGEMA_signal_12714 ), .Q ( new_AGEMA_signal_12785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4761 ( .C ( clk ), .D ( new_AGEMA_signal_12788 ), .Q ( new_AGEMA_signal_12789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4765 ( .C ( clk ), .D ( new_AGEMA_signal_12792 ), .Q ( new_AGEMA_signal_12793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4769 ( .C ( clk ), .D ( new_AGEMA_signal_12796 ), .Q ( new_AGEMA_signal_12797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4773 ( .C ( clk ), .D ( new_AGEMA_signal_12800 ), .Q ( new_AGEMA_signal_12801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4781 ( .C ( clk ), .D ( new_AGEMA_signal_12808 ), .Q ( new_AGEMA_signal_12809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4789 ( .C ( clk ), .D ( new_AGEMA_signal_12816 ), .Q ( new_AGEMA_signal_12817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4797 ( .C ( clk ), .D ( new_AGEMA_signal_12824 ), .Q ( new_AGEMA_signal_12825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4805 ( .C ( clk ), .D ( new_AGEMA_signal_12832 ), .Q ( new_AGEMA_signal_12833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4813 ( .C ( clk ), .D ( new_AGEMA_signal_12840 ), .Q ( new_AGEMA_signal_12841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4821 ( .C ( clk ), .D ( new_AGEMA_signal_12848 ), .Q ( new_AGEMA_signal_12849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4829 ( .C ( clk ), .D ( new_AGEMA_signal_12856 ), .Q ( new_AGEMA_signal_12857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4837 ( .C ( clk ), .D ( new_AGEMA_signal_12864 ), .Q ( new_AGEMA_signal_12865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4845 ( .C ( clk ), .D ( new_AGEMA_signal_12872 ), .Q ( new_AGEMA_signal_12873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4853 ( .C ( clk ), .D ( new_AGEMA_signal_12880 ), .Q ( new_AGEMA_signal_12881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4861 ( .C ( clk ), .D ( new_AGEMA_signal_12888 ), .Q ( new_AGEMA_signal_12889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4869 ( .C ( clk ), .D ( new_AGEMA_signal_12896 ), .Q ( new_AGEMA_signal_12897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4877 ( .C ( clk ), .D ( new_AGEMA_signal_12904 ), .Q ( new_AGEMA_signal_12905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4885 ( .C ( clk ), .D ( new_AGEMA_signal_12912 ), .Q ( new_AGEMA_signal_12913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4893 ( .C ( clk ), .D ( new_AGEMA_signal_12920 ), .Q ( new_AGEMA_signal_12921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4901 ( .C ( clk ), .D ( new_AGEMA_signal_12928 ), .Q ( new_AGEMA_signal_12929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4907 ( .C ( clk ), .D ( new_AGEMA_signal_12934 ), .Q ( new_AGEMA_signal_12935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4913 ( .C ( clk ), .D ( new_AGEMA_signal_12940 ), .Q ( new_AGEMA_signal_12941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4919 ( .C ( clk ), .D ( new_AGEMA_signal_12946 ), .Q ( new_AGEMA_signal_12947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4925 ( .C ( clk ), .D ( new_AGEMA_signal_12952 ), .Q ( new_AGEMA_signal_12953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4935 ( .C ( clk ), .D ( new_AGEMA_signal_12962 ), .Q ( new_AGEMA_signal_12963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4945 ( .C ( clk ), .D ( new_AGEMA_signal_12972 ), .Q ( new_AGEMA_signal_12973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4955 ( .C ( clk ), .D ( new_AGEMA_signal_12982 ), .Q ( new_AGEMA_signal_12983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4965 ( .C ( clk ), .D ( new_AGEMA_signal_12992 ), .Q ( new_AGEMA_signal_12993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4973 ( .C ( clk ), .D ( new_AGEMA_signal_13000 ), .Q ( new_AGEMA_signal_13001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4981 ( .C ( clk ), .D ( new_AGEMA_signal_13008 ), .Q ( new_AGEMA_signal_13009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4989 ( .C ( clk ), .D ( new_AGEMA_signal_13016 ), .Q ( new_AGEMA_signal_13017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4997 ( .C ( clk ), .D ( new_AGEMA_signal_13024 ), .Q ( new_AGEMA_signal_13025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5005 ( .C ( clk ), .D ( new_AGEMA_signal_13032 ), .Q ( new_AGEMA_signal_13033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5013 ( .C ( clk ), .D ( new_AGEMA_signal_13040 ), .Q ( new_AGEMA_signal_13041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5021 ( .C ( clk ), .D ( new_AGEMA_signal_13048 ), .Q ( new_AGEMA_signal_13049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5029 ( .C ( clk ), .D ( new_AGEMA_signal_13056 ), .Q ( new_AGEMA_signal_13057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5037 ( .C ( clk ), .D ( new_AGEMA_signal_13064 ), .Q ( new_AGEMA_signal_13065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5045 ( .C ( clk ), .D ( new_AGEMA_signal_13072 ), .Q ( new_AGEMA_signal_13073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5053 ( .C ( clk ), .D ( new_AGEMA_signal_13080 ), .Q ( new_AGEMA_signal_13081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5061 ( .C ( clk ), .D ( new_AGEMA_signal_13088 ), .Q ( new_AGEMA_signal_13089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5063 ( .C ( clk ), .D ( new_AGEMA_signal_12148 ), .Q ( new_AGEMA_signal_13091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5065 ( .C ( clk ), .D ( new_AGEMA_signal_12150 ), .Q ( new_AGEMA_signal_13093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5067 ( .C ( clk ), .D ( new_AGEMA_signal_12152 ), .Q ( new_AGEMA_signal_13095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5069 ( .C ( clk ), .D ( new_AGEMA_signal_12154 ), .Q ( new_AGEMA_signal_13097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5073 ( .C ( clk ), .D ( new_AGEMA_signal_13100 ), .Q ( new_AGEMA_signal_13101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5077 ( .C ( clk ), .D ( new_AGEMA_signal_13104 ), .Q ( new_AGEMA_signal_13105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5081 ( .C ( clk ), .D ( new_AGEMA_signal_13108 ), .Q ( new_AGEMA_signal_13109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5085 ( .C ( clk ), .D ( new_AGEMA_signal_13112 ), .Q ( new_AGEMA_signal_13113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5091 ( .C ( clk ), .D ( new_AGEMA_signal_13118 ), .Q ( new_AGEMA_signal_13119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5097 ( .C ( clk ), .D ( new_AGEMA_signal_13124 ), .Q ( new_AGEMA_signal_13125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5103 ( .C ( clk ), .D ( new_AGEMA_signal_13130 ), .Q ( new_AGEMA_signal_13131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5109 ( .C ( clk ), .D ( new_AGEMA_signal_13136 ), .Q ( new_AGEMA_signal_13137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5113 ( .C ( clk ), .D ( new_AGEMA_signal_13140 ), .Q ( new_AGEMA_signal_13141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5117 ( .C ( clk ), .D ( new_AGEMA_signal_13144 ), .Q ( new_AGEMA_signal_13145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5121 ( .C ( clk ), .D ( new_AGEMA_signal_13148 ), .Q ( new_AGEMA_signal_13149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5125 ( .C ( clk ), .D ( new_AGEMA_signal_13152 ), .Q ( new_AGEMA_signal_13153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5135 ( .C ( clk ), .D ( new_AGEMA_signal_13162 ), .Q ( new_AGEMA_signal_13163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5145 ( .C ( clk ), .D ( new_AGEMA_signal_13172 ), .Q ( new_AGEMA_signal_13173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5155 ( .C ( clk ), .D ( new_AGEMA_signal_13182 ), .Q ( new_AGEMA_signal_13183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5165 ( .C ( clk ), .D ( new_AGEMA_signal_13192 ), .Q ( new_AGEMA_signal_13193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5173 ( .C ( clk ), .D ( new_AGEMA_signal_13200 ), .Q ( new_AGEMA_signal_13201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5181 ( .C ( clk ), .D ( new_AGEMA_signal_13208 ), .Q ( new_AGEMA_signal_13209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5189 ( .C ( clk ), .D ( new_AGEMA_signal_13216 ), .Q ( new_AGEMA_signal_13217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C ( clk ), .D ( new_AGEMA_signal_13224 ), .Q ( new_AGEMA_signal_13225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C ( clk ), .D ( new_AGEMA_signal_13228 ), .Q ( new_AGEMA_signal_13229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C ( clk ), .D ( new_AGEMA_signal_13232 ), .Q ( new_AGEMA_signal_13233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C ( clk ), .D ( new_AGEMA_signal_13236 ), .Q ( new_AGEMA_signal_13237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C ( clk ), .D ( new_AGEMA_signal_13240 ), .Q ( new_AGEMA_signal_13241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C ( clk ), .D ( n2509 ), .Q ( new_AGEMA_signal_13243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C ( clk ), .D ( new_AGEMA_signal_3387 ), .Q ( new_AGEMA_signal_13245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C ( clk ), .D ( new_AGEMA_signal_3388 ), .Q ( new_AGEMA_signal_13247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C ( clk ), .D ( new_AGEMA_signal_3389 ), .Q ( new_AGEMA_signal_13249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C ( clk ), .D ( new_AGEMA_signal_13256 ), .Q ( new_AGEMA_signal_13257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C ( clk ), .D ( new_AGEMA_signal_13264 ), .Q ( new_AGEMA_signal_13265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C ( clk ), .D ( new_AGEMA_signal_13272 ), .Q ( new_AGEMA_signal_13273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5253 ( .C ( clk ), .D ( new_AGEMA_signal_13280 ), .Q ( new_AGEMA_signal_13281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5261 ( .C ( clk ), .D ( new_AGEMA_signal_13288 ), .Q ( new_AGEMA_signal_13289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5269 ( .C ( clk ), .D ( new_AGEMA_signal_13296 ), .Q ( new_AGEMA_signal_13297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5277 ( .C ( clk ), .D ( new_AGEMA_signal_13304 ), .Q ( new_AGEMA_signal_13305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5285 ( .C ( clk ), .D ( new_AGEMA_signal_13312 ), .Q ( new_AGEMA_signal_13313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5291 ( .C ( clk ), .D ( new_AGEMA_signal_13318 ), .Q ( new_AGEMA_signal_13319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5297 ( .C ( clk ), .D ( new_AGEMA_signal_13324 ), .Q ( new_AGEMA_signal_13325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5303 ( .C ( clk ), .D ( new_AGEMA_signal_13330 ), .Q ( new_AGEMA_signal_13331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5309 ( .C ( clk ), .D ( new_AGEMA_signal_13336 ), .Q ( new_AGEMA_signal_13337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5313 ( .C ( clk ), .D ( new_AGEMA_signal_13340 ), .Q ( new_AGEMA_signal_13341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5317 ( .C ( clk ), .D ( new_AGEMA_signal_13344 ), .Q ( new_AGEMA_signal_13345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5321 ( .C ( clk ), .D ( new_AGEMA_signal_13348 ), .Q ( new_AGEMA_signal_13349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5325 ( .C ( clk ), .D ( new_AGEMA_signal_13352 ), .Q ( new_AGEMA_signal_13353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5333 ( .C ( clk ), .D ( new_AGEMA_signal_13360 ), .Q ( new_AGEMA_signal_13361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5341 ( .C ( clk ), .D ( new_AGEMA_signal_13368 ), .Q ( new_AGEMA_signal_13369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5349 ( .C ( clk ), .D ( new_AGEMA_signal_13376 ), .Q ( new_AGEMA_signal_13377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5357 ( .C ( clk ), .D ( new_AGEMA_signal_13384 ), .Q ( new_AGEMA_signal_13385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5359 ( .C ( clk ), .D ( n2802 ), .Q ( new_AGEMA_signal_13387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5361 ( .C ( clk ), .D ( new_AGEMA_signal_3285 ), .Q ( new_AGEMA_signal_13389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5363 ( .C ( clk ), .D ( new_AGEMA_signal_3286 ), .Q ( new_AGEMA_signal_13391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5365 ( .C ( clk ), .D ( new_AGEMA_signal_3287 ), .Q ( new_AGEMA_signal_13393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5369 ( .C ( clk ), .D ( new_AGEMA_signal_13396 ), .Q ( new_AGEMA_signal_13397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5375 ( .C ( clk ), .D ( new_AGEMA_signal_13402 ), .Q ( new_AGEMA_signal_13403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5381 ( .C ( clk ), .D ( new_AGEMA_signal_13408 ), .Q ( new_AGEMA_signal_13409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5387 ( .C ( clk ), .D ( new_AGEMA_signal_13414 ), .Q ( new_AGEMA_signal_13415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5393 ( .C ( clk ), .D ( new_AGEMA_signal_13420 ), .Q ( new_AGEMA_signal_13421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5399 ( .C ( clk ), .D ( new_AGEMA_signal_13426 ), .Q ( new_AGEMA_signal_13427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5405 ( .C ( clk ), .D ( new_AGEMA_signal_13432 ), .Q ( new_AGEMA_signal_13433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5411 ( .C ( clk ), .D ( new_AGEMA_signal_13438 ), .Q ( new_AGEMA_signal_13439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5417 ( .C ( clk ), .D ( new_AGEMA_signal_13444 ), .Q ( new_AGEMA_signal_13445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5423 ( .C ( clk ), .D ( new_AGEMA_signal_13450 ), .Q ( new_AGEMA_signal_13451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5429 ( .C ( clk ), .D ( new_AGEMA_signal_13456 ), .Q ( new_AGEMA_signal_13457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5435 ( .C ( clk ), .D ( new_AGEMA_signal_13462 ), .Q ( new_AGEMA_signal_13463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5439 ( .C ( clk ), .D ( new_AGEMA_signal_12748 ), .Q ( new_AGEMA_signal_13467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5443 ( .C ( clk ), .D ( new_AGEMA_signal_12750 ), .Q ( new_AGEMA_signal_13471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5447 ( .C ( clk ), .D ( new_AGEMA_signal_12752 ), .Q ( new_AGEMA_signal_13475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5451 ( .C ( clk ), .D ( new_AGEMA_signal_12754 ), .Q ( new_AGEMA_signal_13479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5459 ( .C ( clk ), .D ( new_AGEMA_signal_13486 ), .Q ( new_AGEMA_signal_13487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5467 ( .C ( clk ), .D ( new_AGEMA_signal_13494 ), .Q ( new_AGEMA_signal_13495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5475 ( .C ( clk ), .D ( new_AGEMA_signal_13502 ), .Q ( new_AGEMA_signal_13503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5483 ( .C ( clk ), .D ( new_AGEMA_signal_13510 ), .Q ( new_AGEMA_signal_13511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5489 ( .C ( clk ), .D ( new_AGEMA_signal_13516 ), .Q ( new_AGEMA_signal_13517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5495 ( .C ( clk ), .D ( new_AGEMA_signal_13522 ), .Q ( new_AGEMA_signal_13523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5501 ( .C ( clk ), .D ( new_AGEMA_signal_13528 ), .Q ( new_AGEMA_signal_13529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5507 ( .C ( clk ), .D ( new_AGEMA_signal_13534 ), .Q ( new_AGEMA_signal_13535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5511 ( .C ( clk ), .D ( n2072 ), .Q ( new_AGEMA_signal_13539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5515 ( .C ( clk ), .D ( new_AGEMA_signal_3144 ), .Q ( new_AGEMA_signal_13543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5519 ( .C ( clk ), .D ( new_AGEMA_signal_3145 ), .Q ( new_AGEMA_signal_13547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5523 ( .C ( clk ), .D ( new_AGEMA_signal_3146 ), .Q ( new_AGEMA_signal_13551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5531 ( .C ( clk ), .D ( new_AGEMA_signal_13558 ), .Q ( new_AGEMA_signal_13559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5539 ( .C ( clk ), .D ( new_AGEMA_signal_13566 ), .Q ( new_AGEMA_signal_13567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5547 ( .C ( clk ), .D ( new_AGEMA_signal_13574 ), .Q ( new_AGEMA_signal_13575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5555 ( .C ( clk ), .D ( new_AGEMA_signal_13582 ), .Q ( new_AGEMA_signal_13583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5563 ( .C ( clk ), .D ( new_AGEMA_signal_13590 ), .Q ( new_AGEMA_signal_13591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5571 ( .C ( clk ), .D ( new_AGEMA_signal_13598 ), .Q ( new_AGEMA_signal_13599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5579 ( .C ( clk ), .D ( new_AGEMA_signal_13606 ), .Q ( new_AGEMA_signal_13607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5587 ( .C ( clk ), .D ( new_AGEMA_signal_13614 ), .Q ( new_AGEMA_signal_13615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5597 ( .C ( clk ), .D ( new_AGEMA_signal_13624 ), .Q ( new_AGEMA_signal_13625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5607 ( .C ( clk ), .D ( new_AGEMA_signal_13634 ), .Q ( new_AGEMA_signal_13635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5617 ( .C ( clk ), .D ( new_AGEMA_signal_13644 ), .Q ( new_AGEMA_signal_13645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5627 ( .C ( clk ), .D ( new_AGEMA_signal_13654 ), .Q ( new_AGEMA_signal_13655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5635 ( .C ( clk ), .D ( new_AGEMA_signal_13662 ), .Q ( new_AGEMA_signal_13663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5643 ( .C ( clk ), .D ( new_AGEMA_signal_13670 ), .Q ( new_AGEMA_signal_13671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5651 ( .C ( clk ), .D ( new_AGEMA_signal_13678 ), .Q ( new_AGEMA_signal_13679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5659 ( .C ( clk ), .D ( new_AGEMA_signal_13686 ), .Q ( new_AGEMA_signal_13687 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5665 ( .C ( clk ), .D ( new_AGEMA_signal_13692 ), .Q ( new_AGEMA_signal_13693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5671 ( .C ( clk ), .D ( new_AGEMA_signal_13698 ), .Q ( new_AGEMA_signal_13699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5677 ( .C ( clk ), .D ( new_AGEMA_signal_13704 ), .Q ( new_AGEMA_signal_13705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5683 ( .C ( clk ), .D ( new_AGEMA_signal_13710 ), .Q ( new_AGEMA_signal_13711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5687 ( .C ( clk ), .D ( n2276 ), .Q ( new_AGEMA_signal_13715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5691 ( .C ( clk ), .D ( new_AGEMA_signal_3192 ), .Q ( new_AGEMA_signal_13719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5695 ( .C ( clk ), .D ( new_AGEMA_signal_3193 ), .Q ( new_AGEMA_signal_13723 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5699 ( .C ( clk ), .D ( new_AGEMA_signal_3194 ), .Q ( new_AGEMA_signal_13727 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5705 ( .C ( clk ), .D ( new_AGEMA_signal_13732 ), .Q ( new_AGEMA_signal_13733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5711 ( .C ( clk ), .D ( new_AGEMA_signal_13738 ), .Q ( new_AGEMA_signal_13739 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5717 ( .C ( clk ), .D ( new_AGEMA_signal_13744 ), .Q ( new_AGEMA_signal_13745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5723 ( .C ( clk ), .D ( new_AGEMA_signal_13750 ), .Q ( new_AGEMA_signal_13751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5731 ( .C ( clk ), .D ( new_AGEMA_signal_13758 ), .Q ( new_AGEMA_signal_13759 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5739 ( .C ( clk ), .D ( new_AGEMA_signal_13766 ), .Q ( new_AGEMA_signal_13767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5747 ( .C ( clk ), .D ( new_AGEMA_signal_13774 ), .Q ( new_AGEMA_signal_13775 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5755 ( .C ( clk ), .D ( new_AGEMA_signal_13782 ), .Q ( new_AGEMA_signal_13783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5761 ( .C ( clk ), .D ( new_AGEMA_signal_13788 ), .Q ( new_AGEMA_signal_13789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5767 ( .C ( clk ), .D ( new_AGEMA_signal_13794 ), .Q ( new_AGEMA_signal_13795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5773 ( .C ( clk ), .D ( new_AGEMA_signal_13800 ), .Q ( new_AGEMA_signal_13801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5779 ( .C ( clk ), .D ( new_AGEMA_signal_13806 ), .Q ( new_AGEMA_signal_13807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5795 ( .C ( clk ), .D ( new_AGEMA_signal_13822 ), .Q ( new_AGEMA_signal_13823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5803 ( .C ( clk ), .D ( new_AGEMA_signal_13830 ), .Q ( new_AGEMA_signal_13831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5811 ( .C ( clk ), .D ( new_AGEMA_signal_13838 ), .Q ( new_AGEMA_signal_13839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5819 ( .C ( clk ), .D ( new_AGEMA_signal_13846 ), .Q ( new_AGEMA_signal_13847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5823 ( .C ( clk ), .D ( n2622 ), .Q ( new_AGEMA_signal_13851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5827 ( .C ( clk ), .D ( new_AGEMA_signal_3261 ), .Q ( new_AGEMA_signal_13855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5831 ( .C ( clk ), .D ( new_AGEMA_signal_3262 ), .Q ( new_AGEMA_signal_13859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5835 ( .C ( clk ), .D ( new_AGEMA_signal_3263 ), .Q ( new_AGEMA_signal_13863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5841 ( .C ( clk ), .D ( new_AGEMA_signal_13868 ), .Q ( new_AGEMA_signal_13869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5847 ( .C ( clk ), .D ( new_AGEMA_signal_13874 ), .Q ( new_AGEMA_signal_13875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5853 ( .C ( clk ), .D ( new_AGEMA_signal_13880 ), .Q ( new_AGEMA_signal_13881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5859 ( .C ( clk ), .D ( new_AGEMA_signal_13886 ), .Q ( new_AGEMA_signal_13887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5865 ( .C ( clk ), .D ( new_AGEMA_signal_13892 ), .Q ( new_AGEMA_signal_13893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5871 ( .C ( clk ), .D ( new_AGEMA_signal_13898 ), .Q ( new_AGEMA_signal_13899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5877 ( .C ( clk ), .D ( new_AGEMA_signal_13904 ), .Q ( new_AGEMA_signal_13905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5883 ( .C ( clk ), .D ( new_AGEMA_signal_13910 ), .Q ( new_AGEMA_signal_13911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5887 ( .C ( clk ), .D ( n2804 ), .Q ( new_AGEMA_signal_13915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5891 ( .C ( clk ), .D ( new_AGEMA_signal_3282 ), .Q ( new_AGEMA_signal_13919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5895 ( .C ( clk ), .D ( new_AGEMA_signal_3283 ), .Q ( new_AGEMA_signal_13923 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5899 ( .C ( clk ), .D ( new_AGEMA_signal_3284 ), .Q ( new_AGEMA_signal_13927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5903 ( .C ( clk ), .D ( n1990 ), .Q ( new_AGEMA_signal_13931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5909 ( .C ( clk ), .D ( new_AGEMA_signal_2886 ), .Q ( new_AGEMA_signal_13937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5915 ( .C ( clk ), .D ( new_AGEMA_signal_2887 ), .Q ( new_AGEMA_signal_13943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5921 ( .C ( clk ), .D ( new_AGEMA_signal_2888 ), .Q ( new_AGEMA_signal_13949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5943 ( .C ( clk ), .D ( n2078 ), .Q ( new_AGEMA_signal_13971 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5949 ( .C ( clk ), .D ( new_AGEMA_signal_3150 ), .Q ( new_AGEMA_signal_13977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5955 ( .C ( clk ), .D ( new_AGEMA_signal_3151 ), .Q ( new_AGEMA_signal_13983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5961 ( .C ( clk ), .D ( new_AGEMA_signal_3152 ), .Q ( new_AGEMA_signal_13989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5971 ( .C ( clk ), .D ( new_AGEMA_signal_13998 ), .Q ( new_AGEMA_signal_13999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5981 ( .C ( clk ), .D ( new_AGEMA_signal_14008 ), .Q ( new_AGEMA_signal_14009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5991 ( .C ( clk ), .D ( new_AGEMA_signal_14018 ), .Q ( new_AGEMA_signal_14019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6001 ( .C ( clk ), .D ( new_AGEMA_signal_14028 ), .Q ( new_AGEMA_signal_14029 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6007 ( .C ( clk ), .D ( n2128 ), .Q ( new_AGEMA_signal_14035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6013 ( .C ( clk ), .D ( new_AGEMA_signal_3321 ), .Q ( new_AGEMA_signal_14041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6019 ( .C ( clk ), .D ( new_AGEMA_signal_3322 ), .Q ( new_AGEMA_signal_14047 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C ( clk ), .D ( new_AGEMA_signal_3323 ), .Q ( new_AGEMA_signal_14053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C ( clk ), .D ( n2148 ), .Q ( new_AGEMA_signal_14059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C ( clk ), .D ( new_AGEMA_signal_2940 ), .Q ( new_AGEMA_signal_14065 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C ( clk ), .D ( new_AGEMA_signal_2941 ), .Q ( new_AGEMA_signal_14071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6049 ( .C ( clk ), .D ( new_AGEMA_signal_2942 ), .Q ( new_AGEMA_signal_14077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6089 ( .C ( clk ), .D ( new_AGEMA_signal_14116 ), .Q ( new_AGEMA_signal_14117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6097 ( .C ( clk ), .D ( new_AGEMA_signal_14124 ), .Q ( new_AGEMA_signal_14125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6105 ( .C ( clk ), .D ( new_AGEMA_signal_14132 ), .Q ( new_AGEMA_signal_14133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6113 ( .C ( clk ), .D ( new_AGEMA_signal_14140 ), .Q ( new_AGEMA_signal_14141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6119 ( .C ( clk ), .D ( n2306 ), .Q ( new_AGEMA_signal_14147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6125 ( .C ( clk ), .D ( new_AGEMA_signal_2979 ), .Q ( new_AGEMA_signal_14153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6131 ( .C ( clk ), .D ( new_AGEMA_signal_2980 ), .Q ( new_AGEMA_signal_14159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6137 ( .C ( clk ), .D ( new_AGEMA_signal_2981 ), .Q ( new_AGEMA_signal_14165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6145 ( .C ( clk ), .D ( new_AGEMA_signal_14172 ), .Q ( new_AGEMA_signal_14173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6153 ( .C ( clk ), .D ( new_AGEMA_signal_14180 ), .Q ( new_AGEMA_signal_14181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6161 ( .C ( clk ), .D ( new_AGEMA_signal_14188 ), .Q ( new_AGEMA_signal_14189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6169 ( .C ( clk ), .D ( new_AGEMA_signal_14196 ), .Q ( new_AGEMA_signal_14197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6177 ( .C ( clk ), .D ( new_AGEMA_signal_14204 ), .Q ( new_AGEMA_signal_14205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6185 ( .C ( clk ), .D ( new_AGEMA_signal_14212 ), .Q ( new_AGEMA_signal_14213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6193 ( .C ( clk ), .D ( new_AGEMA_signal_14220 ), .Q ( new_AGEMA_signal_14221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6201 ( .C ( clk ), .D ( new_AGEMA_signal_14228 ), .Q ( new_AGEMA_signal_14229 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6249 ( .C ( clk ), .D ( new_AGEMA_signal_14276 ), .Q ( new_AGEMA_signal_14277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6257 ( .C ( clk ), .D ( new_AGEMA_signal_14284 ), .Q ( new_AGEMA_signal_14285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6265 ( .C ( clk ), .D ( new_AGEMA_signal_14292 ), .Q ( new_AGEMA_signal_14293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6273 ( .C ( clk ), .D ( new_AGEMA_signal_14300 ), .Q ( new_AGEMA_signal_14301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6295 ( .C ( clk ), .D ( n1999 ), .Q ( new_AGEMA_signal_14323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6303 ( .C ( clk ), .D ( new_AGEMA_signal_3129 ), .Q ( new_AGEMA_signal_14331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6311 ( .C ( clk ), .D ( new_AGEMA_signal_3130 ), .Q ( new_AGEMA_signal_14339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6319 ( .C ( clk ), .D ( new_AGEMA_signal_3131 ), .Q ( new_AGEMA_signal_14347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6331 ( .C ( clk ), .D ( new_AGEMA_signal_14358 ), .Q ( new_AGEMA_signal_14359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6343 ( .C ( clk ), .D ( new_AGEMA_signal_14370 ), .Q ( new_AGEMA_signal_14371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6355 ( .C ( clk ), .D ( new_AGEMA_signal_14382 ), .Q ( new_AGEMA_signal_14383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6367 ( .C ( clk ), .D ( new_AGEMA_signal_14394 ), .Q ( new_AGEMA_signal_14395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6381 ( .C ( clk ), .D ( new_AGEMA_signal_14408 ), .Q ( new_AGEMA_signal_14409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6395 ( .C ( clk ), .D ( new_AGEMA_signal_14422 ), .Q ( new_AGEMA_signal_14423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6409 ( .C ( clk ), .D ( new_AGEMA_signal_14436 ), .Q ( new_AGEMA_signal_14437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6423 ( .C ( clk ), .D ( new_AGEMA_signal_14450 ), .Q ( new_AGEMA_signal_14451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6431 ( .C ( clk ), .D ( n2205 ), .Q ( new_AGEMA_signal_14459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6439 ( .C ( clk ), .D ( new_AGEMA_signal_3339 ), .Q ( new_AGEMA_signal_14467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6447 ( .C ( clk ), .D ( new_AGEMA_signal_3340 ), .Q ( new_AGEMA_signal_14475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6455 ( .C ( clk ), .D ( new_AGEMA_signal_3341 ), .Q ( new_AGEMA_signal_14483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6469 ( .C ( clk ), .D ( new_AGEMA_signal_14496 ), .Q ( new_AGEMA_signal_14497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6483 ( .C ( clk ), .D ( new_AGEMA_signal_14510 ), .Q ( new_AGEMA_signal_14511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6497 ( .C ( clk ), .D ( new_AGEMA_signal_14524 ), .Q ( new_AGEMA_signal_14525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6511 ( .C ( clk ), .D ( new_AGEMA_signal_14538 ), .Q ( new_AGEMA_signal_14539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6519 ( .C ( clk ), .D ( n2516 ), .Q ( new_AGEMA_signal_14547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6527 ( .C ( clk ), .D ( new_AGEMA_signal_3228 ), .Q ( new_AGEMA_signal_14555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6535 ( .C ( clk ), .D ( new_AGEMA_signal_3229 ), .Q ( new_AGEMA_signal_14563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6543 ( .C ( clk ), .D ( new_AGEMA_signal_3230 ), .Q ( new_AGEMA_signal_14571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6551 ( .C ( clk ), .D ( n2808 ), .Q ( new_AGEMA_signal_14579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6559 ( .C ( clk ), .D ( new_AGEMA_signal_3273 ), .Q ( new_AGEMA_signal_14587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6567 ( .C ( clk ), .D ( new_AGEMA_signal_3274 ), .Q ( new_AGEMA_signal_14595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6575 ( .C ( clk ), .D ( new_AGEMA_signal_3275 ), .Q ( new_AGEMA_signal_14603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6613 ( .C ( clk ), .D ( new_AGEMA_signal_14640 ), .Q ( new_AGEMA_signal_14641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6629 ( .C ( clk ), .D ( new_AGEMA_signal_14656 ), .Q ( new_AGEMA_signal_14657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6645 ( .C ( clk ), .D ( new_AGEMA_signal_14672 ), .Q ( new_AGEMA_signal_14673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6661 ( .C ( clk ), .D ( new_AGEMA_signal_14688 ), .Q ( new_AGEMA_signal_14689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6701 ( .C ( clk ), .D ( new_AGEMA_signal_14728 ), .Q ( new_AGEMA_signal_14729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6717 ( .C ( clk ), .D ( new_AGEMA_signal_14744 ), .Q ( new_AGEMA_signal_14745 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6733 ( .C ( clk ), .D ( new_AGEMA_signal_14760 ), .Q ( new_AGEMA_signal_14761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6749 ( .C ( clk ), .D ( new_AGEMA_signal_14776 ), .Q ( new_AGEMA_signal_14777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6759 ( .C ( clk ), .D ( n2527 ), .Q ( new_AGEMA_signal_14787 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6769 ( .C ( clk ), .D ( new_AGEMA_signal_3390 ), .Q ( new_AGEMA_signal_14797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6779 ( .C ( clk ), .D ( new_AGEMA_signal_3391 ), .Q ( new_AGEMA_signal_14807 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6789 ( .C ( clk ), .D ( new_AGEMA_signal_3392 ), .Q ( new_AGEMA_signal_14817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6899 ( .C ( clk ), .D ( new_AGEMA_signal_14926 ), .Q ( new_AGEMA_signal_14927 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6915 ( .C ( clk ), .D ( new_AGEMA_signal_14942 ), .Q ( new_AGEMA_signal_14943 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6931 ( .C ( clk ), .D ( new_AGEMA_signal_14958 ), .Q ( new_AGEMA_signal_14959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6947 ( .C ( clk ), .D ( new_AGEMA_signal_14974 ), .Q ( new_AGEMA_signal_14975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7005 ( .C ( clk ), .D ( new_AGEMA_signal_15032 ), .Q ( new_AGEMA_signal_15033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7023 ( .C ( clk ), .D ( new_AGEMA_signal_15050 ), .Q ( new_AGEMA_signal_15051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7041 ( .C ( clk ), .D ( new_AGEMA_signal_15068 ), .Q ( new_AGEMA_signal_15069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7059 ( .C ( clk ), .D ( new_AGEMA_signal_15086 ), .Q ( new_AGEMA_signal_15087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7205 ( .C ( clk ), .D ( new_AGEMA_signal_15232 ), .Q ( new_AGEMA_signal_15233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7225 ( .C ( clk ), .D ( new_AGEMA_signal_15252 ), .Q ( new_AGEMA_signal_15253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7245 ( .C ( clk ), .D ( new_AGEMA_signal_15272 ), .Q ( new_AGEMA_signal_15273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7265 ( .C ( clk ), .D ( new_AGEMA_signal_15292 ), .Q ( new_AGEMA_signal_15293 ) ) ;

    /* cells in depth 14 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2002 ( .a ({new_AGEMA_signal_12058, new_AGEMA_signal_12056, new_AGEMA_signal_12054, new_AGEMA_signal_12052}), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, n1933}), .clk ( clk ), .r ({Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338]}), .c ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n1935}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2054 ( .a ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, n1958}), .b ({new_AGEMA_signal_12090, new_AGEMA_signal_12082, new_AGEMA_signal_12074, new_AGEMA_signal_12066}), .clk ( clk ), .r ({Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344]}), .c ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, new_AGEMA_signal_3297, n1959}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2109 ( .a ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, n1982}), .b ({new_AGEMA_signal_12098, new_AGEMA_signal_12096, new_AGEMA_signal_12094, new_AGEMA_signal_12092}), .clk ( clk ), .r ({Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350]}), .c ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, n1983}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2149 ( .a ({new_AGEMA_signal_12114, new_AGEMA_signal_12110, new_AGEMA_signal_12106, new_AGEMA_signal_12102}), .b ({new_AGEMA_signal_3134, new_AGEMA_signal_3133, new_AGEMA_signal_3132, n2011}), .clk ( clk ), .r ({Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356]}), .c ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, n2014}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2166 ( .a ({new_AGEMA_signal_12146, new_AGEMA_signal_12138, new_AGEMA_signal_12130, new_AGEMA_signal_12122}), .b ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, n2025}), .clk ( clk ), .r ({Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, n2029}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2180 ( .a ({new_AGEMA_signal_12154, new_AGEMA_signal_12152, new_AGEMA_signal_12150, new_AGEMA_signal_12148}), .b ({new_AGEMA_signal_3140, new_AGEMA_signal_3139, new_AGEMA_signal_3138, n2036}), .clk ( clk ), .r ({Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368]}), .c ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, n2037}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2197 ( .a ({new_AGEMA_signal_12178, new_AGEMA_signal_12172, new_AGEMA_signal_12166, new_AGEMA_signal_12160}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, n2049}), .clk ( clk ), .r ({Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374]}), .c ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, n2052}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2219 ( .a ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, n2067}), .b ({new_AGEMA_signal_12194, new_AGEMA_signal_12190, new_AGEMA_signal_12186, new_AGEMA_signal_12182}), .clk ( clk ), .r ({Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, n2070}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2258 ( .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, n2097}), .b ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, n2096}), .clk ( clk ), .r ({Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386]}), .c ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2098}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2287 ( .a ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, n2124}), .b ({new_AGEMA_signal_12226, new_AGEMA_signal_12218, new_AGEMA_signal_12210, new_AGEMA_signal_12202}), .clk ( clk ), .r ({Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392]}), .c ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, n2125}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2311 ( .a ({new_AGEMA_signal_12242, new_AGEMA_signal_12238, new_AGEMA_signal_12234, new_AGEMA_signal_12230}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, n2142}), .clk ( clk ), .r ({Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398]}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, n2145}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2333 ( .a ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, n2168}), .b ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, n2167}), .clk ( clk ), .r ({Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404]}), .c ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2169}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2350 ( .a ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, n2184}), .b ({new_AGEMA_signal_12266, new_AGEMA_signal_12260, new_AGEMA_signal_12254, new_AGEMA_signal_12248}), .clk ( clk ), .r ({Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410]}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, n2185}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2365 ( .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, n2197}), .b ({new_AGEMA_signal_12290, new_AGEMA_signal_12284, new_AGEMA_signal_12278, new_AGEMA_signal_12272}), .clk ( clk ), .r ({Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416]}), .c ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, n2198}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2396 ( .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, n2232}), .b ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, n2231}), .clk ( clk ), .r ({Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422]}), .c ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, n2312}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2404 ( .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, n2239}), .b ({new_AGEMA_signal_12314, new_AGEMA_signal_12308, new_AGEMA_signal_12302, new_AGEMA_signal_12296}), .clk ( clk ), .r ({Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, new_AGEMA_signal_3459, n2258}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2415 ( .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, n2250}), .b ({new_AGEMA_signal_12338, new_AGEMA_signal_12332, new_AGEMA_signal_12326, new_AGEMA_signal_12320}), .clk ( clk ), .r ({Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434]}), .c ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, n2251}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2440 ( .a ({new_AGEMA_signal_12362, new_AGEMA_signal_12356, new_AGEMA_signal_12350, new_AGEMA_signal_12344}), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, n2272}), .clk ( clk ), .r ({Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440]}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, n2274}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2469 ( .a ({new_AGEMA_signal_12378, new_AGEMA_signal_12374, new_AGEMA_signal_12370, new_AGEMA_signal_12366}), .b ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, n2296}), .clk ( clk ), .r ({Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446]}), .c ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2302}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2490 ( .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, n2324}), .b ({new_AGEMA_signal_12410, new_AGEMA_signal_12402, new_AGEMA_signal_12394, new_AGEMA_signal_12386}), .clk ( clk ), .r ({Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452]}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, n2339}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2503 ( .a ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, n2337}), .b ({new_AGEMA_signal_12426, new_AGEMA_signal_12422, new_AGEMA_signal_12418, new_AGEMA_signal_12414}), .clk ( clk ), .r ({Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458]}), .c ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, n2338}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2515 ( .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, n2350}), .b ({new_AGEMA_signal_12450, new_AGEMA_signal_12444, new_AGEMA_signal_12438, new_AGEMA_signal_12432}), .clk ( clk ), .r ({Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, n2351}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2529 ( .a ({new_AGEMA_signal_12482, new_AGEMA_signal_12474, new_AGEMA_signal_12466, new_AGEMA_signal_12458}), .b ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, n2362}), .clk ( clk ), .r ({Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470]}), .c ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2365}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2551 ( .a ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, n2389}), .b ({new_AGEMA_signal_12490, new_AGEMA_signal_12488, new_AGEMA_signal_12486, new_AGEMA_signal_12484}), .clk ( clk ), .r ({Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, n2399}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2560 ( .a ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, n2397}), .b ({new_AGEMA_signal_12514, new_AGEMA_signal_12508, new_AGEMA_signal_12502, new_AGEMA_signal_12496}), .clk ( clk ), .r ({Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482]}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, n2398}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2572 ( .a ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, n2411}), .b ({new_AGEMA_signal_12522, new_AGEMA_signal_12520, new_AGEMA_signal_12518, new_AGEMA_signal_12516}), .clk ( clk ), .r ({Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, n2423}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2581 ( .a ({new_AGEMA_signal_12530, new_AGEMA_signal_12528, new_AGEMA_signal_12526, new_AGEMA_signal_12524}), .b ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, n2420}), .clk ( clk ), .r ({Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494]}), .c ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2422}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2596 ( .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, n2440}), .b ({new_AGEMA_signal_12554, new_AGEMA_signal_12548, new_AGEMA_signal_12542, new_AGEMA_signal_12536}), .clk ( clk ), .r ({Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500]}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, n2441}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2623 ( .a ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, n2471}), .b ({new_AGEMA_signal_12578, new_AGEMA_signal_12572, new_AGEMA_signal_12566, new_AGEMA_signal_12560}), .clk ( clk ), .r ({Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, n2479}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2637 ( .a ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, n2485}), .b ({new_AGEMA_signal_12610, new_AGEMA_signal_12602, new_AGEMA_signal_12594, new_AGEMA_signal_12586}), .clk ( clk ), .r ({Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512]}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, n2512}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2652 ( .a ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, n2502}), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, n2501}), .clk ( clk ), .r ({Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518]}), .c ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, n2510}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2686 ( .a ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, n2550}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, n2549}), .clk ( clk ), .r ({Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524]}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, n2552}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2702 ( .a ({new_AGEMA_signal_12642, new_AGEMA_signal_12634, new_AGEMA_signal_12626, new_AGEMA_signal_12618}), .b ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, n2569}), .clk ( clk ), .r ({Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530]}), .c ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, n2593}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2713 ( .a ({new_AGEMA_signal_12666, new_AGEMA_signal_12660, new_AGEMA_signal_12654, new_AGEMA_signal_12648}), .b ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, n2584}), .clk ( clk ), .r ({Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, n2589}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2730 ( .a ({new_AGEMA_signal_12690, new_AGEMA_signal_12684, new_AGEMA_signal_12678, new_AGEMA_signal_12672}), .b ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, n2606}), .clk ( clk ), .r ({Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542]}), .c ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2608}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2748 ( .a ({new_AGEMA_signal_12698, new_AGEMA_signal_12696, new_AGEMA_signal_12694, new_AGEMA_signal_12692}), .b ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, n2634}), .clk ( clk ), .r ({Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548]}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, n2636}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2762 ( .a ({new_AGEMA_signal_12714, new_AGEMA_signal_12710, new_AGEMA_signal_12706, new_AGEMA_signal_12702}), .b ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, n2657}), .clk ( clk ), .r ({Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554]}), .c ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, n2659}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2784 ( .a ({new_AGEMA_signal_12730, new_AGEMA_signal_12726, new_AGEMA_signal_12722, new_AGEMA_signal_12718}), .b ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, n2697}), .clk ( clk ), .r ({Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560]}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, n2702}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2811 ( .a ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, n2747}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, n2746}), .clk ( clk ), .r ({Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566]}), .c ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, n2806}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2839 ( .a ({new_AGEMA_signal_12746, new_AGEMA_signal_12742, new_AGEMA_signal_12738, new_AGEMA_signal_12734}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, n2799}), .clk ( clk ), .r ({Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572]}), .c ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, n2801}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2853 ( .a ({new_AGEMA_signal_12754, new_AGEMA_signal_12752, new_AGEMA_signal_12750, new_AGEMA_signal_12748}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, new_AGEMA_signal_3291, n2827}), .clk ( clk ), .r ({Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578]}), .c ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, n2829}) ) ;
    buf_clk new_AGEMA_reg_buffer_4732 ( .C ( clk ), .D ( new_AGEMA_signal_12759 ), .Q ( new_AGEMA_signal_12760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4738 ( .C ( clk ), .D ( new_AGEMA_signal_12765 ), .Q ( new_AGEMA_signal_12766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4744 ( .C ( clk ), .D ( new_AGEMA_signal_12771 ), .Q ( new_AGEMA_signal_12772 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4750 ( .C ( clk ), .D ( new_AGEMA_signal_12777 ), .Q ( new_AGEMA_signal_12778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4752 ( .C ( clk ), .D ( new_AGEMA_signal_12779 ), .Q ( new_AGEMA_signal_12780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4754 ( .C ( clk ), .D ( new_AGEMA_signal_12781 ), .Q ( new_AGEMA_signal_12782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4756 ( .C ( clk ), .D ( new_AGEMA_signal_12783 ), .Q ( new_AGEMA_signal_12784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4758 ( .C ( clk ), .D ( new_AGEMA_signal_12785 ), .Q ( new_AGEMA_signal_12786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4762 ( .C ( clk ), .D ( new_AGEMA_signal_12789 ), .Q ( new_AGEMA_signal_12790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4766 ( .C ( clk ), .D ( new_AGEMA_signal_12793 ), .Q ( new_AGEMA_signal_12794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4770 ( .C ( clk ), .D ( new_AGEMA_signal_12797 ), .Q ( new_AGEMA_signal_12798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4774 ( .C ( clk ), .D ( new_AGEMA_signal_12801 ), .Q ( new_AGEMA_signal_12802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4782 ( .C ( clk ), .D ( new_AGEMA_signal_12809 ), .Q ( new_AGEMA_signal_12810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4790 ( .C ( clk ), .D ( new_AGEMA_signal_12817 ), .Q ( new_AGEMA_signal_12818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4798 ( .C ( clk ), .D ( new_AGEMA_signal_12825 ), .Q ( new_AGEMA_signal_12826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4806 ( .C ( clk ), .D ( new_AGEMA_signal_12833 ), .Q ( new_AGEMA_signal_12834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4814 ( .C ( clk ), .D ( new_AGEMA_signal_12841 ), .Q ( new_AGEMA_signal_12842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4822 ( .C ( clk ), .D ( new_AGEMA_signal_12849 ), .Q ( new_AGEMA_signal_12850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4830 ( .C ( clk ), .D ( new_AGEMA_signal_12857 ), .Q ( new_AGEMA_signal_12858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4838 ( .C ( clk ), .D ( new_AGEMA_signal_12865 ), .Q ( new_AGEMA_signal_12866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4846 ( .C ( clk ), .D ( new_AGEMA_signal_12873 ), .Q ( new_AGEMA_signal_12874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4854 ( .C ( clk ), .D ( new_AGEMA_signal_12881 ), .Q ( new_AGEMA_signal_12882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4862 ( .C ( clk ), .D ( new_AGEMA_signal_12889 ), .Q ( new_AGEMA_signal_12890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4870 ( .C ( clk ), .D ( new_AGEMA_signal_12897 ), .Q ( new_AGEMA_signal_12898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4878 ( .C ( clk ), .D ( new_AGEMA_signal_12905 ), .Q ( new_AGEMA_signal_12906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4886 ( .C ( clk ), .D ( new_AGEMA_signal_12913 ), .Q ( new_AGEMA_signal_12914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4894 ( .C ( clk ), .D ( new_AGEMA_signal_12921 ), .Q ( new_AGEMA_signal_12922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4902 ( .C ( clk ), .D ( new_AGEMA_signal_12929 ), .Q ( new_AGEMA_signal_12930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4908 ( .C ( clk ), .D ( new_AGEMA_signal_12935 ), .Q ( new_AGEMA_signal_12936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4914 ( .C ( clk ), .D ( new_AGEMA_signal_12941 ), .Q ( new_AGEMA_signal_12942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4920 ( .C ( clk ), .D ( new_AGEMA_signal_12947 ), .Q ( new_AGEMA_signal_12948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4926 ( .C ( clk ), .D ( new_AGEMA_signal_12953 ), .Q ( new_AGEMA_signal_12954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4936 ( .C ( clk ), .D ( new_AGEMA_signal_12963 ), .Q ( new_AGEMA_signal_12964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4946 ( .C ( clk ), .D ( new_AGEMA_signal_12973 ), .Q ( new_AGEMA_signal_12974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4956 ( .C ( clk ), .D ( new_AGEMA_signal_12983 ), .Q ( new_AGEMA_signal_12984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4966 ( .C ( clk ), .D ( new_AGEMA_signal_12993 ), .Q ( new_AGEMA_signal_12994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4974 ( .C ( clk ), .D ( new_AGEMA_signal_13001 ), .Q ( new_AGEMA_signal_13002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4982 ( .C ( clk ), .D ( new_AGEMA_signal_13009 ), .Q ( new_AGEMA_signal_13010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4990 ( .C ( clk ), .D ( new_AGEMA_signal_13017 ), .Q ( new_AGEMA_signal_13018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_4998 ( .C ( clk ), .D ( new_AGEMA_signal_13025 ), .Q ( new_AGEMA_signal_13026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5006 ( .C ( clk ), .D ( new_AGEMA_signal_13033 ), .Q ( new_AGEMA_signal_13034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5014 ( .C ( clk ), .D ( new_AGEMA_signal_13041 ), .Q ( new_AGEMA_signal_13042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5022 ( .C ( clk ), .D ( new_AGEMA_signal_13049 ), .Q ( new_AGEMA_signal_13050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5030 ( .C ( clk ), .D ( new_AGEMA_signal_13057 ), .Q ( new_AGEMA_signal_13058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5038 ( .C ( clk ), .D ( new_AGEMA_signal_13065 ), .Q ( new_AGEMA_signal_13066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5046 ( .C ( clk ), .D ( new_AGEMA_signal_13073 ), .Q ( new_AGEMA_signal_13074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5054 ( .C ( clk ), .D ( new_AGEMA_signal_13081 ), .Q ( new_AGEMA_signal_13082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5062 ( .C ( clk ), .D ( new_AGEMA_signal_13089 ), .Q ( new_AGEMA_signal_13090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5064 ( .C ( clk ), .D ( new_AGEMA_signal_13091 ), .Q ( new_AGEMA_signal_13092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5066 ( .C ( clk ), .D ( new_AGEMA_signal_13093 ), .Q ( new_AGEMA_signal_13094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5068 ( .C ( clk ), .D ( new_AGEMA_signal_13095 ), .Q ( new_AGEMA_signal_13096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5070 ( .C ( clk ), .D ( new_AGEMA_signal_13097 ), .Q ( new_AGEMA_signal_13098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5074 ( .C ( clk ), .D ( new_AGEMA_signal_13101 ), .Q ( new_AGEMA_signal_13102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5078 ( .C ( clk ), .D ( new_AGEMA_signal_13105 ), .Q ( new_AGEMA_signal_13106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5082 ( .C ( clk ), .D ( new_AGEMA_signal_13109 ), .Q ( new_AGEMA_signal_13110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5086 ( .C ( clk ), .D ( new_AGEMA_signal_13113 ), .Q ( new_AGEMA_signal_13114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5092 ( .C ( clk ), .D ( new_AGEMA_signal_13119 ), .Q ( new_AGEMA_signal_13120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5098 ( .C ( clk ), .D ( new_AGEMA_signal_13125 ), .Q ( new_AGEMA_signal_13126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5104 ( .C ( clk ), .D ( new_AGEMA_signal_13131 ), .Q ( new_AGEMA_signal_13132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5110 ( .C ( clk ), .D ( new_AGEMA_signal_13137 ), .Q ( new_AGEMA_signal_13138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5114 ( .C ( clk ), .D ( new_AGEMA_signal_13141 ), .Q ( new_AGEMA_signal_13142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5118 ( .C ( clk ), .D ( new_AGEMA_signal_13145 ), .Q ( new_AGEMA_signal_13146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5122 ( .C ( clk ), .D ( new_AGEMA_signal_13149 ), .Q ( new_AGEMA_signal_13150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5126 ( .C ( clk ), .D ( new_AGEMA_signal_13153 ), .Q ( new_AGEMA_signal_13154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5136 ( .C ( clk ), .D ( new_AGEMA_signal_13163 ), .Q ( new_AGEMA_signal_13164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5146 ( .C ( clk ), .D ( new_AGEMA_signal_13173 ), .Q ( new_AGEMA_signal_13174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5156 ( .C ( clk ), .D ( new_AGEMA_signal_13183 ), .Q ( new_AGEMA_signal_13184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5166 ( .C ( clk ), .D ( new_AGEMA_signal_13193 ), .Q ( new_AGEMA_signal_13194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5174 ( .C ( clk ), .D ( new_AGEMA_signal_13201 ), .Q ( new_AGEMA_signal_13202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5182 ( .C ( clk ), .D ( new_AGEMA_signal_13209 ), .Q ( new_AGEMA_signal_13210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5190 ( .C ( clk ), .D ( new_AGEMA_signal_13217 ), .Q ( new_AGEMA_signal_13218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C ( clk ), .D ( new_AGEMA_signal_13225 ), .Q ( new_AGEMA_signal_13226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C ( clk ), .D ( new_AGEMA_signal_13229 ), .Q ( new_AGEMA_signal_13230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C ( clk ), .D ( new_AGEMA_signal_13233 ), .Q ( new_AGEMA_signal_13234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C ( clk ), .D ( new_AGEMA_signal_13237 ), .Q ( new_AGEMA_signal_13238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C ( clk ), .D ( new_AGEMA_signal_13241 ), .Q ( new_AGEMA_signal_13242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C ( clk ), .D ( new_AGEMA_signal_13243 ), .Q ( new_AGEMA_signal_13244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C ( clk ), .D ( new_AGEMA_signal_13245 ), .Q ( new_AGEMA_signal_13246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C ( clk ), .D ( new_AGEMA_signal_13247 ), .Q ( new_AGEMA_signal_13248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C ( clk ), .D ( new_AGEMA_signal_13249 ), .Q ( new_AGEMA_signal_13250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C ( clk ), .D ( new_AGEMA_signal_13257 ), .Q ( new_AGEMA_signal_13258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C ( clk ), .D ( new_AGEMA_signal_13265 ), .Q ( new_AGEMA_signal_13266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C ( clk ), .D ( new_AGEMA_signal_13273 ), .Q ( new_AGEMA_signal_13274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5254 ( .C ( clk ), .D ( new_AGEMA_signal_13281 ), .Q ( new_AGEMA_signal_13282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5262 ( .C ( clk ), .D ( new_AGEMA_signal_13289 ), .Q ( new_AGEMA_signal_13290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5270 ( .C ( clk ), .D ( new_AGEMA_signal_13297 ), .Q ( new_AGEMA_signal_13298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5278 ( .C ( clk ), .D ( new_AGEMA_signal_13305 ), .Q ( new_AGEMA_signal_13306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5286 ( .C ( clk ), .D ( new_AGEMA_signal_13313 ), .Q ( new_AGEMA_signal_13314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5292 ( .C ( clk ), .D ( new_AGEMA_signal_13319 ), .Q ( new_AGEMA_signal_13320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5298 ( .C ( clk ), .D ( new_AGEMA_signal_13325 ), .Q ( new_AGEMA_signal_13326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5304 ( .C ( clk ), .D ( new_AGEMA_signal_13331 ), .Q ( new_AGEMA_signal_13332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5310 ( .C ( clk ), .D ( new_AGEMA_signal_13337 ), .Q ( new_AGEMA_signal_13338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5314 ( .C ( clk ), .D ( new_AGEMA_signal_13341 ), .Q ( new_AGEMA_signal_13342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5318 ( .C ( clk ), .D ( new_AGEMA_signal_13345 ), .Q ( new_AGEMA_signal_13346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5322 ( .C ( clk ), .D ( new_AGEMA_signal_13349 ), .Q ( new_AGEMA_signal_13350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5326 ( .C ( clk ), .D ( new_AGEMA_signal_13353 ), .Q ( new_AGEMA_signal_13354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5334 ( .C ( clk ), .D ( new_AGEMA_signal_13361 ), .Q ( new_AGEMA_signal_13362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5342 ( .C ( clk ), .D ( new_AGEMA_signal_13369 ), .Q ( new_AGEMA_signal_13370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5350 ( .C ( clk ), .D ( new_AGEMA_signal_13377 ), .Q ( new_AGEMA_signal_13378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5358 ( .C ( clk ), .D ( new_AGEMA_signal_13385 ), .Q ( new_AGEMA_signal_13386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5360 ( .C ( clk ), .D ( new_AGEMA_signal_13387 ), .Q ( new_AGEMA_signal_13388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5362 ( .C ( clk ), .D ( new_AGEMA_signal_13389 ), .Q ( new_AGEMA_signal_13390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5364 ( .C ( clk ), .D ( new_AGEMA_signal_13391 ), .Q ( new_AGEMA_signal_13392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5366 ( .C ( clk ), .D ( new_AGEMA_signal_13393 ), .Q ( new_AGEMA_signal_13394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5370 ( .C ( clk ), .D ( new_AGEMA_signal_13397 ), .Q ( new_AGEMA_signal_13398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5376 ( .C ( clk ), .D ( new_AGEMA_signal_13403 ), .Q ( new_AGEMA_signal_13404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5382 ( .C ( clk ), .D ( new_AGEMA_signal_13409 ), .Q ( new_AGEMA_signal_13410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5388 ( .C ( clk ), .D ( new_AGEMA_signal_13415 ), .Q ( new_AGEMA_signal_13416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5394 ( .C ( clk ), .D ( new_AGEMA_signal_13421 ), .Q ( new_AGEMA_signal_13422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5400 ( .C ( clk ), .D ( new_AGEMA_signal_13427 ), .Q ( new_AGEMA_signal_13428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5406 ( .C ( clk ), .D ( new_AGEMA_signal_13433 ), .Q ( new_AGEMA_signal_13434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5412 ( .C ( clk ), .D ( new_AGEMA_signal_13439 ), .Q ( new_AGEMA_signal_13440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5418 ( .C ( clk ), .D ( new_AGEMA_signal_13445 ), .Q ( new_AGEMA_signal_13446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5424 ( .C ( clk ), .D ( new_AGEMA_signal_13451 ), .Q ( new_AGEMA_signal_13452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5430 ( .C ( clk ), .D ( new_AGEMA_signal_13457 ), .Q ( new_AGEMA_signal_13458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5436 ( .C ( clk ), .D ( new_AGEMA_signal_13463 ), .Q ( new_AGEMA_signal_13464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5440 ( .C ( clk ), .D ( new_AGEMA_signal_13467 ), .Q ( new_AGEMA_signal_13468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5444 ( .C ( clk ), .D ( new_AGEMA_signal_13471 ), .Q ( new_AGEMA_signal_13472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5448 ( .C ( clk ), .D ( new_AGEMA_signal_13475 ), .Q ( new_AGEMA_signal_13476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5452 ( .C ( clk ), .D ( new_AGEMA_signal_13479 ), .Q ( new_AGEMA_signal_13480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5460 ( .C ( clk ), .D ( new_AGEMA_signal_13487 ), .Q ( new_AGEMA_signal_13488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5468 ( .C ( clk ), .D ( new_AGEMA_signal_13495 ), .Q ( new_AGEMA_signal_13496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5476 ( .C ( clk ), .D ( new_AGEMA_signal_13503 ), .Q ( new_AGEMA_signal_13504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5484 ( .C ( clk ), .D ( new_AGEMA_signal_13511 ), .Q ( new_AGEMA_signal_13512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5490 ( .C ( clk ), .D ( new_AGEMA_signal_13517 ), .Q ( new_AGEMA_signal_13518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5496 ( .C ( clk ), .D ( new_AGEMA_signal_13523 ), .Q ( new_AGEMA_signal_13524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5502 ( .C ( clk ), .D ( new_AGEMA_signal_13529 ), .Q ( new_AGEMA_signal_13530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5508 ( .C ( clk ), .D ( new_AGEMA_signal_13535 ), .Q ( new_AGEMA_signal_13536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5512 ( .C ( clk ), .D ( new_AGEMA_signal_13539 ), .Q ( new_AGEMA_signal_13540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5516 ( .C ( clk ), .D ( new_AGEMA_signal_13543 ), .Q ( new_AGEMA_signal_13544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5520 ( .C ( clk ), .D ( new_AGEMA_signal_13547 ), .Q ( new_AGEMA_signal_13548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5524 ( .C ( clk ), .D ( new_AGEMA_signal_13551 ), .Q ( new_AGEMA_signal_13552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5532 ( .C ( clk ), .D ( new_AGEMA_signal_13559 ), .Q ( new_AGEMA_signal_13560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5540 ( .C ( clk ), .D ( new_AGEMA_signal_13567 ), .Q ( new_AGEMA_signal_13568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5548 ( .C ( clk ), .D ( new_AGEMA_signal_13575 ), .Q ( new_AGEMA_signal_13576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5556 ( .C ( clk ), .D ( new_AGEMA_signal_13583 ), .Q ( new_AGEMA_signal_13584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5564 ( .C ( clk ), .D ( new_AGEMA_signal_13591 ), .Q ( new_AGEMA_signal_13592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5572 ( .C ( clk ), .D ( new_AGEMA_signal_13599 ), .Q ( new_AGEMA_signal_13600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5580 ( .C ( clk ), .D ( new_AGEMA_signal_13607 ), .Q ( new_AGEMA_signal_13608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5588 ( .C ( clk ), .D ( new_AGEMA_signal_13615 ), .Q ( new_AGEMA_signal_13616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5598 ( .C ( clk ), .D ( new_AGEMA_signal_13625 ), .Q ( new_AGEMA_signal_13626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5608 ( .C ( clk ), .D ( new_AGEMA_signal_13635 ), .Q ( new_AGEMA_signal_13636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5618 ( .C ( clk ), .D ( new_AGEMA_signal_13645 ), .Q ( new_AGEMA_signal_13646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5628 ( .C ( clk ), .D ( new_AGEMA_signal_13655 ), .Q ( new_AGEMA_signal_13656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5636 ( .C ( clk ), .D ( new_AGEMA_signal_13663 ), .Q ( new_AGEMA_signal_13664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5644 ( .C ( clk ), .D ( new_AGEMA_signal_13671 ), .Q ( new_AGEMA_signal_13672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5652 ( .C ( clk ), .D ( new_AGEMA_signal_13679 ), .Q ( new_AGEMA_signal_13680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5660 ( .C ( clk ), .D ( new_AGEMA_signal_13687 ), .Q ( new_AGEMA_signal_13688 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5666 ( .C ( clk ), .D ( new_AGEMA_signal_13693 ), .Q ( new_AGEMA_signal_13694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5672 ( .C ( clk ), .D ( new_AGEMA_signal_13699 ), .Q ( new_AGEMA_signal_13700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5678 ( .C ( clk ), .D ( new_AGEMA_signal_13705 ), .Q ( new_AGEMA_signal_13706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5684 ( .C ( clk ), .D ( new_AGEMA_signal_13711 ), .Q ( new_AGEMA_signal_13712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5688 ( .C ( clk ), .D ( new_AGEMA_signal_13715 ), .Q ( new_AGEMA_signal_13716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5692 ( .C ( clk ), .D ( new_AGEMA_signal_13719 ), .Q ( new_AGEMA_signal_13720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5696 ( .C ( clk ), .D ( new_AGEMA_signal_13723 ), .Q ( new_AGEMA_signal_13724 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5700 ( .C ( clk ), .D ( new_AGEMA_signal_13727 ), .Q ( new_AGEMA_signal_13728 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5706 ( .C ( clk ), .D ( new_AGEMA_signal_13733 ), .Q ( new_AGEMA_signal_13734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5712 ( .C ( clk ), .D ( new_AGEMA_signal_13739 ), .Q ( new_AGEMA_signal_13740 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5718 ( .C ( clk ), .D ( new_AGEMA_signal_13745 ), .Q ( new_AGEMA_signal_13746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5724 ( .C ( clk ), .D ( new_AGEMA_signal_13751 ), .Q ( new_AGEMA_signal_13752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5732 ( .C ( clk ), .D ( new_AGEMA_signal_13759 ), .Q ( new_AGEMA_signal_13760 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5740 ( .C ( clk ), .D ( new_AGEMA_signal_13767 ), .Q ( new_AGEMA_signal_13768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5748 ( .C ( clk ), .D ( new_AGEMA_signal_13775 ), .Q ( new_AGEMA_signal_13776 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5756 ( .C ( clk ), .D ( new_AGEMA_signal_13783 ), .Q ( new_AGEMA_signal_13784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5762 ( .C ( clk ), .D ( new_AGEMA_signal_13789 ), .Q ( new_AGEMA_signal_13790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5768 ( .C ( clk ), .D ( new_AGEMA_signal_13795 ), .Q ( new_AGEMA_signal_13796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5774 ( .C ( clk ), .D ( new_AGEMA_signal_13801 ), .Q ( new_AGEMA_signal_13802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5780 ( .C ( clk ), .D ( new_AGEMA_signal_13807 ), .Q ( new_AGEMA_signal_13808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5796 ( .C ( clk ), .D ( new_AGEMA_signal_13823 ), .Q ( new_AGEMA_signal_13824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5804 ( .C ( clk ), .D ( new_AGEMA_signal_13831 ), .Q ( new_AGEMA_signal_13832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5812 ( .C ( clk ), .D ( new_AGEMA_signal_13839 ), .Q ( new_AGEMA_signal_13840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5820 ( .C ( clk ), .D ( new_AGEMA_signal_13847 ), .Q ( new_AGEMA_signal_13848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5824 ( .C ( clk ), .D ( new_AGEMA_signal_13851 ), .Q ( new_AGEMA_signal_13852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5828 ( .C ( clk ), .D ( new_AGEMA_signal_13855 ), .Q ( new_AGEMA_signal_13856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5832 ( .C ( clk ), .D ( new_AGEMA_signal_13859 ), .Q ( new_AGEMA_signal_13860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5836 ( .C ( clk ), .D ( new_AGEMA_signal_13863 ), .Q ( new_AGEMA_signal_13864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5842 ( .C ( clk ), .D ( new_AGEMA_signal_13869 ), .Q ( new_AGEMA_signal_13870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5848 ( .C ( clk ), .D ( new_AGEMA_signal_13875 ), .Q ( new_AGEMA_signal_13876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5854 ( .C ( clk ), .D ( new_AGEMA_signal_13881 ), .Q ( new_AGEMA_signal_13882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5860 ( .C ( clk ), .D ( new_AGEMA_signal_13887 ), .Q ( new_AGEMA_signal_13888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5866 ( .C ( clk ), .D ( new_AGEMA_signal_13893 ), .Q ( new_AGEMA_signal_13894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5872 ( .C ( clk ), .D ( new_AGEMA_signal_13899 ), .Q ( new_AGEMA_signal_13900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5878 ( .C ( clk ), .D ( new_AGEMA_signal_13905 ), .Q ( new_AGEMA_signal_13906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5884 ( .C ( clk ), .D ( new_AGEMA_signal_13911 ), .Q ( new_AGEMA_signal_13912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5888 ( .C ( clk ), .D ( new_AGEMA_signal_13915 ), .Q ( new_AGEMA_signal_13916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5892 ( .C ( clk ), .D ( new_AGEMA_signal_13919 ), .Q ( new_AGEMA_signal_13920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5896 ( .C ( clk ), .D ( new_AGEMA_signal_13923 ), .Q ( new_AGEMA_signal_13924 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5900 ( .C ( clk ), .D ( new_AGEMA_signal_13927 ), .Q ( new_AGEMA_signal_13928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5904 ( .C ( clk ), .D ( new_AGEMA_signal_13931 ), .Q ( new_AGEMA_signal_13932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5910 ( .C ( clk ), .D ( new_AGEMA_signal_13937 ), .Q ( new_AGEMA_signal_13938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5916 ( .C ( clk ), .D ( new_AGEMA_signal_13943 ), .Q ( new_AGEMA_signal_13944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5922 ( .C ( clk ), .D ( new_AGEMA_signal_13949 ), .Q ( new_AGEMA_signal_13950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5944 ( .C ( clk ), .D ( new_AGEMA_signal_13971 ), .Q ( new_AGEMA_signal_13972 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5950 ( .C ( clk ), .D ( new_AGEMA_signal_13977 ), .Q ( new_AGEMA_signal_13978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5956 ( .C ( clk ), .D ( new_AGEMA_signal_13983 ), .Q ( new_AGEMA_signal_13984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5962 ( .C ( clk ), .D ( new_AGEMA_signal_13989 ), .Q ( new_AGEMA_signal_13990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5972 ( .C ( clk ), .D ( new_AGEMA_signal_13999 ), .Q ( new_AGEMA_signal_14000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5982 ( .C ( clk ), .D ( new_AGEMA_signal_14009 ), .Q ( new_AGEMA_signal_14010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5992 ( .C ( clk ), .D ( new_AGEMA_signal_14019 ), .Q ( new_AGEMA_signal_14020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6002 ( .C ( clk ), .D ( new_AGEMA_signal_14029 ), .Q ( new_AGEMA_signal_14030 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6008 ( .C ( clk ), .D ( new_AGEMA_signal_14035 ), .Q ( new_AGEMA_signal_14036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6014 ( .C ( clk ), .D ( new_AGEMA_signal_14041 ), .Q ( new_AGEMA_signal_14042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6020 ( .C ( clk ), .D ( new_AGEMA_signal_14047 ), .Q ( new_AGEMA_signal_14048 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C ( clk ), .D ( new_AGEMA_signal_14053 ), .Q ( new_AGEMA_signal_14054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C ( clk ), .D ( new_AGEMA_signal_14059 ), .Q ( new_AGEMA_signal_14060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C ( clk ), .D ( new_AGEMA_signal_14065 ), .Q ( new_AGEMA_signal_14066 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C ( clk ), .D ( new_AGEMA_signal_14071 ), .Q ( new_AGEMA_signal_14072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6050 ( .C ( clk ), .D ( new_AGEMA_signal_14077 ), .Q ( new_AGEMA_signal_14078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6090 ( .C ( clk ), .D ( new_AGEMA_signal_14117 ), .Q ( new_AGEMA_signal_14118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6098 ( .C ( clk ), .D ( new_AGEMA_signal_14125 ), .Q ( new_AGEMA_signal_14126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6106 ( .C ( clk ), .D ( new_AGEMA_signal_14133 ), .Q ( new_AGEMA_signal_14134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6114 ( .C ( clk ), .D ( new_AGEMA_signal_14141 ), .Q ( new_AGEMA_signal_14142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6120 ( .C ( clk ), .D ( new_AGEMA_signal_14147 ), .Q ( new_AGEMA_signal_14148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6126 ( .C ( clk ), .D ( new_AGEMA_signal_14153 ), .Q ( new_AGEMA_signal_14154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6132 ( .C ( clk ), .D ( new_AGEMA_signal_14159 ), .Q ( new_AGEMA_signal_14160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6138 ( .C ( clk ), .D ( new_AGEMA_signal_14165 ), .Q ( new_AGEMA_signal_14166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6146 ( .C ( clk ), .D ( new_AGEMA_signal_14173 ), .Q ( new_AGEMA_signal_14174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6154 ( .C ( clk ), .D ( new_AGEMA_signal_14181 ), .Q ( new_AGEMA_signal_14182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6162 ( .C ( clk ), .D ( new_AGEMA_signal_14189 ), .Q ( new_AGEMA_signal_14190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6170 ( .C ( clk ), .D ( new_AGEMA_signal_14197 ), .Q ( new_AGEMA_signal_14198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6178 ( .C ( clk ), .D ( new_AGEMA_signal_14205 ), .Q ( new_AGEMA_signal_14206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6186 ( .C ( clk ), .D ( new_AGEMA_signal_14213 ), .Q ( new_AGEMA_signal_14214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6194 ( .C ( clk ), .D ( new_AGEMA_signal_14221 ), .Q ( new_AGEMA_signal_14222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6202 ( .C ( clk ), .D ( new_AGEMA_signal_14229 ), .Q ( new_AGEMA_signal_14230 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6250 ( .C ( clk ), .D ( new_AGEMA_signal_14277 ), .Q ( new_AGEMA_signal_14278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6258 ( .C ( clk ), .D ( new_AGEMA_signal_14285 ), .Q ( new_AGEMA_signal_14286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6266 ( .C ( clk ), .D ( new_AGEMA_signal_14293 ), .Q ( new_AGEMA_signal_14294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6274 ( .C ( clk ), .D ( new_AGEMA_signal_14301 ), .Q ( new_AGEMA_signal_14302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6296 ( .C ( clk ), .D ( new_AGEMA_signal_14323 ), .Q ( new_AGEMA_signal_14324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6304 ( .C ( clk ), .D ( new_AGEMA_signal_14331 ), .Q ( new_AGEMA_signal_14332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6312 ( .C ( clk ), .D ( new_AGEMA_signal_14339 ), .Q ( new_AGEMA_signal_14340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6320 ( .C ( clk ), .D ( new_AGEMA_signal_14347 ), .Q ( new_AGEMA_signal_14348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6332 ( .C ( clk ), .D ( new_AGEMA_signal_14359 ), .Q ( new_AGEMA_signal_14360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6344 ( .C ( clk ), .D ( new_AGEMA_signal_14371 ), .Q ( new_AGEMA_signal_14372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6356 ( .C ( clk ), .D ( new_AGEMA_signal_14383 ), .Q ( new_AGEMA_signal_14384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6368 ( .C ( clk ), .D ( new_AGEMA_signal_14395 ), .Q ( new_AGEMA_signal_14396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6382 ( .C ( clk ), .D ( new_AGEMA_signal_14409 ), .Q ( new_AGEMA_signal_14410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6396 ( .C ( clk ), .D ( new_AGEMA_signal_14423 ), .Q ( new_AGEMA_signal_14424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6410 ( .C ( clk ), .D ( new_AGEMA_signal_14437 ), .Q ( new_AGEMA_signal_14438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6424 ( .C ( clk ), .D ( new_AGEMA_signal_14451 ), .Q ( new_AGEMA_signal_14452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6432 ( .C ( clk ), .D ( new_AGEMA_signal_14459 ), .Q ( new_AGEMA_signal_14460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6440 ( .C ( clk ), .D ( new_AGEMA_signal_14467 ), .Q ( new_AGEMA_signal_14468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6448 ( .C ( clk ), .D ( new_AGEMA_signal_14475 ), .Q ( new_AGEMA_signal_14476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6456 ( .C ( clk ), .D ( new_AGEMA_signal_14483 ), .Q ( new_AGEMA_signal_14484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6470 ( .C ( clk ), .D ( new_AGEMA_signal_14497 ), .Q ( new_AGEMA_signal_14498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6484 ( .C ( clk ), .D ( new_AGEMA_signal_14511 ), .Q ( new_AGEMA_signal_14512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6498 ( .C ( clk ), .D ( new_AGEMA_signal_14525 ), .Q ( new_AGEMA_signal_14526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6512 ( .C ( clk ), .D ( new_AGEMA_signal_14539 ), .Q ( new_AGEMA_signal_14540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6520 ( .C ( clk ), .D ( new_AGEMA_signal_14547 ), .Q ( new_AGEMA_signal_14548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6528 ( .C ( clk ), .D ( new_AGEMA_signal_14555 ), .Q ( new_AGEMA_signal_14556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6536 ( .C ( clk ), .D ( new_AGEMA_signal_14563 ), .Q ( new_AGEMA_signal_14564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6544 ( .C ( clk ), .D ( new_AGEMA_signal_14571 ), .Q ( new_AGEMA_signal_14572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6552 ( .C ( clk ), .D ( new_AGEMA_signal_14579 ), .Q ( new_AGEMA_signal_14580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6560 ( .C ( clk ), .D ( new_AGEMA_signal_14587 ), .Q ( new_AGEMA_signal_14588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6568 ( .C ( clk ), .D ( new_AGEMA_signal_14595 ), .Q ( new_AGEMA_signal_14596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6576 ( .C ( clk ), .D ( new_AGEMA_signal_14603 ), .Q ( new_AGEMA_signal_14604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6614 ( .C ( clk ), .D ( new_AGEMA_signal_14641 ), .Q ( new_AGEMA_signal_14642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6630 ( .C ( clk ), .D ( new_AGEMA_signal_14657 ), .Q ( new_AGEMA_signal_14658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6646 ( .C ( clk ), .D ( new_AGEMA_signal_14673 ), .Q ( new_AGEMA_signal_14674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6662 ( .C ( clk ), .D ( new_AGEMA_signal_14689 ), .Q ( new_AGEMA_signal_14690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6702 ( .C ( clk ), .D ( new_AGEMA_signal_14729 ), .Q ( new_AGEMA_signal_14730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6718 ( .C ( clk ), .D ( new_AGEMA_signal_14745 ), .Q ( new_AGEMA_signal_14746 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6734 ( .C ( clk ), .D ( new_AGEMA_signal_14761 ), .Q ( new_AGEMA_signal_14762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6750 ( .C ( clk ), .D ( new_AGEMA_signal_14777 ), .Q ( new_AGEMA_signal_14778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6760 ( .C ( clk ), .D ( new_AGEMA_signal_14787 ), .Q ( new_AGEMA_signal_14788 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6770 ( .C ( clk ), .D ( new_AGEMA_signal_14797 ), .Q ( new_AGEMA_signal_14798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6780 ( .C ( clk ), .D ( new_AGEMA_signal_14807 ), .Q ( new_AGEMA_signal_14808 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6790 ( .C ( clk ), .D ( new_AGEMA_signal_14817 ), .Q ( new_AGEMA_signal_14818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6900 ( .C ( clk ), .D ( new_AGEMA_signal_14927 ), .Q ( new_AGEMA_signal_14928 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6916 ( .C ( clk ), .D ( new_AGEMA_signal_14943 ), .Q ( new_AGEMA_signal_14944 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6932 ( .C ( clk ), .D ( new_AGEMA_signal_14959 ), .Q ( new_AGEMA_signal_14960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6948 ( .C ( clk ), .D ( new_AGEMA_signal_14975 ), .Q ( new_AGEMA_signal_14976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7006 ( .C ( clk ), .D ( new_AGEMA_signal_15033 ), .Q ( new_AGEMA_signal_15034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7024 ( .C ( clk ), .D ( new_AGEMA_signal_15051 ), .Q ( new_AGEMA_signal_15052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7042 ( .C ( clk ), .D ( new_AGEMA_signal_15069 ), .Q ( new_AGEMA_signal_15070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7060 ( .C ( clk ), .D ( new_AGEMA_signal_15087 ), .Q ( new_AGEMA_signal_15088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7206 ( .C ( clk ), .D ( new_AGEMA_signal_15233 ), .Q ( new_AGEMA_signal_15234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7226 ( .C ( clk ), .D ( new_AGEMA_signal_15253 ), .Q ( new_AGEMA_signal_15254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7246 ( .C ( clk ), .D ( new_AGEMA_signal_15273 ), .Q ( new_AGEMA_signal_15274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7266 ( .C ( clk ), .D ( new_AGEMA_signal_15293 ), .Q ( new_AGEMA_signal_15294 ) ) ;

    /* cells in depth 15 */
    buf_clk new_AGEMA_reg_buffer_5371 ( .C ( clk ), .D ( new_AGEMA_signal_13398 ), .Q ( new_AGEMA_signal_13399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5377 ( .C ( clk ), .D ( new_AGEMA_signal_13404 ), .Q ( new_AGEMA_signal_13405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5383 ( .C ( clk ), .D ( new_AGEMA_signal_13410 ), .Q ( new_AGEMA_signal_13411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5389 ( .C ( clk ), .D ( new_AGEMA_signal_13416 ), .Q ( new_AGEMA_signal_13417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5395 ( .C ( clk ), .D ( new_AGEMA_signal_13422 ), .Q ( new_AGEMA_signal_13423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5401 ( .C ( clk ), .D ( new_AGEMA_signal_13428 ), .Q ( new_AGEMA_signal_13429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5407 ( .C ( clk ), .D ( new_AGEMA_signal_13434 ), .Q ( new_AGEMA_signal_13435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5413 ( .C ( clk ), .D ( new_AGEMA_signal_13440 ), .Q ( new_AGEMA_signal_13441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5419 ( .C ( clk ), .D ( new_AGEMA_signal_13446 ), .Q ( new_AGEMA_signal_13447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5425 ( .C ( clk ), .D ( new_AGEMA_signal_13452 ), .Q ( new_AGEMA_signal_13453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5431 ( .C ( clk ), .D ( new_AGEMA_signal_13458 ), .Q ( new_AGEMA_signal_13459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5437 ( .C ( clk ), .D ( new_AGEMA_signal_13464 ), .Q ( new_AGEMA_signal_13465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5441 ( .C ( clk ), .D ( new_AGEMA_signal_13468 ), .Q ( new_AGEMA_signal_13469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5445 ( .C ( clk ), .D ( new_AGEMA_signal_13472 ), .Q ( new_AGEMA_signal_13473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5449 ( .C ( clk ), .D ( new_AGEMA_signal_13476 ), .Q ( new_AGEMA_signal_13477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5453 ( .C ( clk ), .D ( new_AGEMA_signal_13480 ), .Q ( new_AGEMA_signal_13481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5461 ( .C ( clk ), .D ( new_AGEMA_signal_13488 ), .Q ( new_AGEMA_signal_13489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5469 ( .C ( clk ), .D ( new_AGEMA_signal_13496 ), .Q ( new_AGEMA_signal_13497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5477 ( .C ( clk ), .D ( new_AGEMA_signal_13504 ), .Q ( new_AGEMA_signal_13505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5485 ( .C ( clk ), .D ( new_AGEMA_signal_13512 ), .Q ( new_AGEMA_signal_13513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5491 ( .C ( clk ), .D ( new_AGEMA_signal_13518 ), .Q ( new_AGEMA_signal_13519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5497 ( .C ( clk ), .D ( new_AGEMA_signal_13524 ), .Q ( new_AGEMA_signal_13525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5503 ( .C ( clk ), .D ( new_AGEMA_signal_13530 ), .Q ( new_AGEMA_signal_13531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5509 ( .C ( clk ), .D ( new_AGEMA_signal_13536 ), .Q ( new_AGEMA_signal_13537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5513 ( .C ( clk ), .D ( new_AGEMA_signal_13540 ), .Q ( new_AGEMA_signal_13541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5517 ( .C ( clk ), .D ( new_AGEMA_signal_13544 ), .Q ( new_AGEMA_signal_13545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5521 ( .C ( clk ), .D ( new_AGEMA_signal_13548 ), .Q ( new_AGEMA_signal_13549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5525 ( .C ( clk ), .D ( new_AGEMA_signal_13552 ), .Q ( new_AGEMA_signal_13553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5533 ( .C ( clk ), .D ( new_AGEMA_signal_13560 ), .Q ( new_AGEMA_signal_13561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5541 ( .C ( clk ), .D ( new_AGEMA_signal_13568 ), .Q ( new_AGEMA_signal_13569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5549 ( .C ( clk ), .D ( new_AGEMA_signal_13576 ), .Q ( new_AGEMA_signal_13577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5557 ( .C ( clk ), .D ( new_AGEMA_signal_13584 ), .Q ( new_AGEMA_signal_13585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5565 ( .C ( clk ), .D ( new_AGEMA_signal_13592 ), .Q ( new_AGEMA_signal_13593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5573 ( .C ( clk ), .D ( new_AGEMA_signal_13600 ), .Q ( new_AGEMA_signal_13601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5581 ( .C ( clk ), .D ( new_AGEMA_signal_13608 ), .Q ( new_AGEMA_signal_13609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5589 ( .C ( clk ), .D ( new_AGEMA_signal_13616 ), .Q ( new_AGEMA_signal_13617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5599 ( .C ( clk ), .D ( new_AGEMA_signal_13626 ), .Q ( new_AGEMA_signal_13627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5609 ( .C ( clk ), .D ( new_AGEMA_signal_13636 ), .Q ( new_AGEMA_signal_13637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5619 ( .C ( clk ), .D ( new_AGEMA_signal_13646 ), .Q ( new_AGEMA_signal_13647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5629 ( .C ( clk ), .D ( new_AGEMA_signal_13656 ), .Q ( new_AGEMA_signal_13657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5637 ( .C ( clk ), .D ( new_AGEMA_signal_13664 ), .Q ( new_AGEMA_signal_13665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5645 ( .C ( clk ), .D ( new_AGEMA_signal_13672 ), .Q ( new_AGEMA_signal_13673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5653 ( .C ( clk ), .D ( new_AGEMA_signal_13680 ), .Q ( new_AGEMA_signal_13681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5661 ( .C ( clk ), .D ( new_AGEMA_signal_13688 ), .Q ( new_AGEMA_signal_13689 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5667 ( .C ( clk ), .D ( new_AGEMA_signal_13694 ), .Q ( new_AGEMA_signal_13695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5673 ( .C ( clk ), .D ( new_AGEMA_signal_13700 ), .Q ( new_AGEMA_signal_13701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5679 ( .C ( clk ), .D ( new_AGEMA_signal_13706 ), .Q ( new_AGEMA_signal_13707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5685 ( .C ( clk ), .D ( new_AGEMA_signal_13712 ), .Q ( new_AGEMA_signal_13713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5689 ( .C ( clk ), .D ( new_AGEMA_signal_13716 ), .Q ( new_AGEMA_signal_13717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5693 ( .C ( clk ), .D ( new_AGEMA_signal_13720 ), .Q ( new_AGEMA_signal_13721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5697 ( .C ( clk ), .D ( new_AGEMA_signal_13724 ), .Q ( new_AGEMA_signal_13725 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5701 ( .C ( clk ), .D ( new_AGEMA_signal_13728 ), .Q ( new_AGEMA_signal_13729 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5707 ( .C ( clk ), .D ( new_AGEMA_signal_13734 ), .Q ( new_AGEMA_signal_13735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5713 ( .C ( clk ), .D ( new_AGEMA_signal_13740 ), .Q ( new_AGEMA_signal_13741 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5719 ( .C ( clk ), .D ( new_AGEMA_signal_13746 ), .Q ( new_AGEMA_signal_13747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5725 ( .C ( clk ), .D ( new_AGEMA_signal_13752 ), .Q ( new_AGEMA_signal_13753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5733 ( .C ( clk ), .D ( new_AGEMA_signal_13760 ), .Q ( new_AGEMA_signal_13761 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5741 ( .C ( clk ), .D ( new_AGEMA_signal_13768 ), .Q ( new_AGEMA_signal_13769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5749 ( .C ( clk ), .D ( new_AGEMA_signal_13776 ), .Q ( new_AGEMA_signal_13777 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5757 ( .C ( clk ), .D ( new_AGEMA_signal_13784 ), .Q ( new_AGEMA_signal_13785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5763 ( .C ( clk ), .D ( new_AGEMA_signal_13790 ), .Q ( new_AGEMA_signal_13791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5769 ( .C ( clk ), .D ( new_AGEMA_signal_13796 ), .Q ( new_AGEMA_signal_13797 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5775 ( .C ( clk ), .D ( new_AGEMA_signal_13802 ), .Q ( new_AGEMA_signal_13803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5781 ( .C ( clk ), .D ( new_AGEMA_signal_13808 ), .Q ( new_AGEMA_signal_13809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5783 ( .C ( clk ), .D ( n2512 ), .Q ( new_AGEMA_signal_13811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5785 ( .C ( clk ), .D ( new_AGEMA_signal_3381 ), .Q ( new_AGEMA_signal_13813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5787 ( .C ( clk ), .D ( new_AGEMA_signal_3382 ), .Q ( new_AGEMA_signal_13815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5789 ( .C ( clk ), .D ( new_AGEMA_signal_3383 ), .Q ( new_AGEMA_signal_13817 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5797 ( .C ( clk ), .D ( new_AGEMA_signal_13824 ), .Q ( new_AGEMA_signal_13825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5805 ( .C ( clk ), .D ( new_AGEMA_signal_13832 ), .Q ( new_AGEMA_signal_13833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5813 ( .C ( clk ), .D ( new_AGEMA_signal_13840 ), .Q ( new_AGEMA_signal_13841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5821 ( .C ( clk ), .D ( new_AGEMA_signal_13848 ), .Q ( new_AGEMA_signal_13849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5825 ( .C ( clk ), .D ( new_AGEMA_signal_13852 ), .Q ( new_AGEMA_signal_13853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5829 ( .C ( clk ), .D ( new_AGEMA_signal_13856 ), .Q ( new_AGEMA_signal_13857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5833 ( .C ( clk ), .D ( new_AGEMA_signal_13860 ), .Q ( new_AGEMA_signal_13861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5837 ( .C ( clk ), .D ( new_AGEMA_signal_13864 ), .Q ( new_AGEMA_signal_13865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5843 ( .C ( clk ), .D ( new_AGEMA_signal_13870 ), .Q ( new_AGEMA_signal_13871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5849 ( .C ( clk ), .D ( new_AGEMA_signal_13876 ), .Q ( new_AGEMA_signal_13877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5855 ( .C ( clk ), .D ( new_AGEMA_signal_13882 ), .Q ( new_AGEMA_signal_13883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5861 ( .C ( clk ), .D ( new_AGEMA_signal_13888 ), .Q ( new_AGEMA_signal_13889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5867 ( .C ( clk ), .D ( new_AGEMA_signal_13894 ), .Q ( new_AGEMA_signal_13895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5873 ( .C ( clk ), .D ( new_AGEMA_signal_13900 ), .Q ( new_AGEMA_signal_13901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5879 ( .C ( clk ), .D ( new_AGEMA_signal_13906 ), .Q ( new_AGEMA_signal_13907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5885 ( .C ( clk ), .D ( new_AGEMA_signal_13912 ), .Q ( new_AGEMA_signal_13913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5889 ( .C ( clk ), .D ( new_AGEMA_signal_13916 ), .Q ( new_AGEMA_signal_13917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5893 ( .C ( clk ), .D ( new_AGEMA_signal_13920 ), .Q ( new_AGEMA_signal_13921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5897 ( .C ( clk ), .D ( new_AGEMA_signal_13924 ), .Q ( new_AGEMA_signal_13925 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5901 ( .C ( clk ), .D ( new_AGEMA_signal_13928 ), .Q ( new_AGEMA_signal_13929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5905 ( .C ( clk ), .D ( new_AGEMA_signal_13932 ), .Q ( new_AGEMA_signal_13933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5911 ( .C ( clk ), .D ( new_AGEMA_signal_13938 ), .Q ( new_AGEMA_signal_13939 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5917 ( .C ( clk ), .D ( new_AGEMA_signal_13944 ), .Q ( new_AGEMA_signal_13945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5923 ( .C ( clk ), .D ( new_AGEMA_signal_13950 ), .Q ( new_AGEMA_signal_13951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5927 ( .C ( clk ), .D ( n2037 ), .Q ( new_AGEMA_signal_13955 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5931 ( .C ( clk ), .D ( new_AGEMA_signal_3309 ), .Q ( new_AGEMA_signal_13959 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5935 ( .C ( clk ), .D ( new_AGEMA_signal_3310 ), .Q ( new_AGEMA_signal_13963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5939 ( .C ( clk ), .D ( new_AGEMA_signal_3311 ), .Q ( new_AGEMA_signal_13967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5945 ( .C ( clk ), .D ( new_AGEMA_signal_13972 ), .Q ( new_AGEMA_signal_13973 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5951 ( .C ( clk ), .D ( new_AGEMA_signal_13978 ), .Q ( new_AGEMA_signal_13979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5957 ( .C ( clk ), .D ( new_AGEMA_signal_13984 ), .Q ( new_AGEMA_signal_13985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5963 ( .C ( clk ), .D ( new_AGEMA_signal_13990 ), .Q ( new_AGEMA_signal_13991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5973 ( .C ( clk ), .D ( new_AGEMA_signal_14000 ), .Q ( new_AGEMA_signal_14001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5983 ( .C ( clk ), .D ( new_AGEMA_signal_14010 ), .Q ( new_AGEMA_signal_14011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5993 ( .C ( clk ), .D ( new_AGEMA_signal_14020 ), .Q ( new_AGEMA_signal_14021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6003 ( .C ( clk ), .D ( new_AGEMA_signal_14030 ), .Q ( new_AGEMA_signal_14031 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6009 ( .C ( clk ), .D ( new_AGEMA_signal_14036 ), .Q ( new_AGEMA_signal_14037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6015 ( .C ( clk ), .D ( new_AGEMA_signal_14042 ), .Q ( new_AGEMA_signal_14043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C ( clk ), .D ( new_AGEMA_signal_14048 ), .Q ( new_AGEMA_signal_14049 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C ( clk ), .D ( new_AGEMA_signal_14054 ), .Q ( new_AGEMA_signal_14055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C ( clk ), .D ( new_AGEMA_signal_14060 ), .Q ( new_AGEMA_signal_14061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C ( clk ), .D ( new_AGEMA_signal_14066 ), .Q ( new_AGEMA_signal_14067 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C ( clk ), .D ( new_AGEMA_signal_14072 ), .Q ( new_AGEMA_signal_14073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6051 ( .C ( clk ), .D ( new_AGEMA_signal_14078 ), .Q ( new_AGEMA_signal_14079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6055 ( .C ( clk ), .D ( n2198 ), .Q ( new_AGEMA_signal_14083 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6059 ( .C ( clk ), .D ( new_AGEMA_signal_3336 ), .Q ( new_AGEMA_signal_14087 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6063 ( .C ( clk ), .D ( new_AGEMA_signal_3337 ), .Q ( new_AGEMA_signal_14091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6067 ( .C ( clk ), .D ( new_AGEMA_signal_3338 ), .Q ( new_AGEMA_signal_14095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6071 ( .C ( clk ), .D ( n2258 ), .Q ( new_AGEMA_signal_14099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6075 ( .C ( clk ), .D ( new_AGEMA_signal_3459 ), .Q ( new_AGEMA_signal_14103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6079 ( .C ( clk ), .D ( new_AGEMA_signal_3460 ), .Q ( new_AGEMA_signal_14107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6083 ( .C ( clk ), .D ( new_AGEMA_signal_3461 ), .Q ( new_AGEMA_signal_14111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6091 ( .C ( clk ), .D ( new_AGEMA_signal_14118 ), .Q ( new_AGEMA_signal_14119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6099 ( .C ( clk ), .D ( new_AGEMA_signal_14126 ), .Q ( new_AGEMA_signal_14127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6107 ( .C ( clk ), .D ( new_AGEMA_signal_14134 ), .Q ( new_AGEMA_signal_14135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6115 ( .C ( clk ), .D ( new_AGEMA_signal_14142 ), .Q ( new_AGEMA_signal_14143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6121 ( .C ( clk ), .D ( new_AGEMA_signal_14148 ), .Q ( new_AGEMA_signal_14149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6127 ( .C ( clk ), .D ( new_AGEMA_signal_14154 ), .Q ( new_AGEMA_signal_14155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6133 ( .C ( clk ), .D ( new_AGEMA_signal_14160 ), .Q ( new_AGEMA_signal_14161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6139 ( .C ( clk ), .D ( new_AGEMA_signal_14166 ), .Q ( new_AGEMA_signal_14167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6147 ( .C ( clk ), .D ( new_AGEMA_signal_14174 ), .Q ( new_AGEMA_signal_14175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6155 ( .C ( clk ), .D ( new_AGEMA_signal_14182 ), .Q ( new_AGEMA_signal_14183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6163 ( .C ( clk ), .D ( new_AGEMA_signal_14190 ), .Q ( new_AGEMA_signal_14191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6171 ( .C ( clk ), .D ( new_AGEMA_signal_14198 ), .Q ( new_AGEMA_signal_14199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6179 ( .C ( clk ), .D ( new_AGEMA_signal_14206 ), .Q ( new_AGEMA_signal_14207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6187 ( .C ( clk ), .D ( new_AGEMA_signal_14214 ), .Q ( new_AGEMA_signal_14215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6195 ( .C ( clk ), .D ( new_AGEMA_signal_14222 ), .Q ( new_AGEMA_signal_14223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6203 ( .C ( clk ), .D ( new_AGEMA_signal_14230 ), .Q ( new_AGEMA_signal_14231 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6215 ( .C ( clk ), .D ( n2593 ), .Q ( new_AGEMA_signal_14243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6219 ( .C ( clk ), .D ( new_AGEMA_signal_3396 ), .Q ( new_AGEMA_signal_14247 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6223 ( .C ( clk ), .D ( new_AGEMA_signal_3397 ), .Q ( new_AGEMA_signal_14251 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6227 ( .C ( clk ), .D ( new_AGEMA_signal_3398 ), .Q ( new_AGEMA_signal_14255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6231 ( .C ( clk ), .D ( n2636 ), .Q ( new_AGEMA_signal_14259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6235 ( .C ( clk ), .D ( new_AGEMA_signal_3405 ), .Q ( new_AGEMA_signal_14263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6239 ( .C ( clk ), .D ( new_AGEMA_signal_3406 ), .Q ( new_AGEMA_signal_14267 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6243 ( .C ( clk ), .D ( new_AGEMA_signal_3407 ), .Q ( new_AGEMA_signal_14271 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6251 ( .C ( clk ), .D ( new_AGEMA_signal_14278 ), .Q ( new_AGEMA_signal_14279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6259 ( .C ( clk ), .D ( new_AGEMA_signal_14286 ), .Q ( new_AGEMA_signal_14287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6267 ( .C ( clk ), .D ( new_AGEMA_signal_14294 ), .Q ( new_AGEMA_signal_14295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6275 ( .C ( clk ), .D ( new_AGEMA_signal_14302 ), .Q ( new_AGEMA_signal_14303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6279 ( .C ( clk ), .D ( n2806 ), .Q ( new_AGEMA_signal_14307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6283 ( .C ( clk ), .D ( new_AGEMA_signal_3414 ), .Q ( new_AGEMA_signal_14311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6287 ( .C ( clk ), .D ( new_AGEMA_signal_3415 ), .Q ( new_AGEMA_signal_14315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6291 ( .C ( clk ), .D ( new_AGEMA_signal_3416 ), .Q ( new_AGEMA_signal_14319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6297 ( .C ( clk ), .D ( new_AGEMA_signal_14324 ), .Q ( new_AGEMA_signal_14325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6305 ( .C ( clk ), .D ( new_AGEMA_signal_14332 ), .Q ( new_AGEMA_signal_14333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6313 ( .C ( clk ), .D ( new_AGEMA_signal_14340 ), .Q ( new_AGEMA_signal_14341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6321 ( .C ( clk ), .D ( new_AGEMA_signal_14348 ), .Q ( new_AGEMA_signal_14349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6333 ( .C ( clk ), .D ( new_AGEMA_signal_14360 ), .Q ( new_AGEMA_signal_14361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6345 ( .C ( clk ), .D ( new_AGEMA_signal_14372 ), .Q ( new_AGEMA_signal_14373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6357 ( .C ( clk ), .D ( new_AGEMA_signal_14384 ), .Q ( new_AGEMA_signal_14385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6369 ( .C ( clk ), .D ( new_AGEMA_signal_14396 ), .Q ( new_AGEMA_signal_14397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6383 ( .C ( clk ), .D ( new_AGEMA_signal_14410 ), .Q ( new_AGEMA_signal_14411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6397 ( .C ( clk ), .D ( new_AGEMA_signal_14424 ), .Q ( new_AGEMA_signal_14425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6411 ( .C ( clk ), .D ( new_AGEMA_signal_14438 ), .Q ( new_AGEMA_signal_14439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6425 ( .C ( clk ), .D ( new_AGEMA_signal_14452 ), .Q ( new_AGEMA_signal_14453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6433 ( .C ( clk ), .D ( new_AGEMA_signal_14460 ), .Q ( new_AGEMA_signal_14461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6441 ( .C ( clk ), .D ( new_AGEMA_signal_14468 ), .Q ( new_AGEMA_signal_14469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6449 ( .C ( clk ), .D ( new_AGEMA_signal_14476 ), .Q ( new_AGEMA_signal_14477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6457 ( .C ( clk ), .D ( new_AGEMA_signal_14484 ), .Q ( new_AGEMA_signal_14485 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6471 ( .C ( clk ), .D ( new_AGEMA_signal_14498 ), .Q ( new_AGEMA_signal_14499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6485 ( .C ( clk ), .D ( new_AGEMA_signal_14512 ), .Q ( new_AGEMA_signal_14513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6499 ( .C ( clk ), .D ( new_AGEMA_signal_14526 ), .Q ( new_AGEMA_signal_14527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6513 ( .C ( clk ), .D ( new_AGEMA_signal_14540 ), .Q ( new_AGEMA_signal_14541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6521 ( .C ( clk ), .D ( new_AGEMA_signal_14548 ), .Q ( new_AGEMA_signal_14549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6529 ( .C ( clk ), .D ( new_AGEMA_signal_14556 ), .Q ( new_AGEMA_signal_14557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6537 ( .C ( clk ), .D ( new_AGEMA_signal_14564 ), .Q ( new_AGEMA_signal_14565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6545 ( .C ( clk ), .D ( new_AGEMA_signal_14572 ), .Q ( new_AGEMA_signal_14573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6553 ( .C ( clk ), .D ( new_AGEMA_signal_14580 ), .Q ( new_AGEMA_signal_14581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6561 ( .C ( clk ), .D ( new_AGEMA_signal_14588 ), .Q ( new_AGEMA_signal_14589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6569 ( .C ( clk ), .D ( new_AGEMA_signal_14596 ), .Q ( new_AGEMA_signal_14597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6577 ( .C ( clk ), .D ( new_AGEMA_signal_14604 ), .Q ( new_AGEMA_signal_14605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6615 ( .C ( clk ), .D ( new_AGEMA_signal_14642 ), .Q ( new_AGEMA_signal_14643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6631 ( .C ( clk ), .D ( new_AGEMA_signal_14658 ), .Q ( new_AGEMA_signal_14659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6647 ( .C ( clk ), .D ( new_AGEMA_signal_14674 ), .Q ( new_AGEMA_signal_14675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6663 ( .C ( clk ), .D ( new_AGEMA_signal_14690 ), .Q ( new_AGEMA_signal_14691 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6703 ( .C ( clk ), .D ( new_AGEMA_signal_14730 ), .Q ( new_AGEMA_signal_14731 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6719 ( .C ( clk ), .D ( new_AGEMA_signal_14746 ), .Q ( new_AGEMA_signal_14747 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6735 ( .C ( clk ), .D ( new_AGEMA_signal_14762 ), .Q ( new_AGEMA_signal_14763 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6751 ( .C ( clk ), .D ( new_AGEMA_signal_14778 ), .Q ( new_AGEMA_signal_14779 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6761 ( .C ( clk ), .D ( new_AGEMA_signal_14788 ), .Q ( new_AGEMA_signal_14789 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6771 ( .C ( clk ), .D ( new_AGEMA_signal_14798 ), .Q ( new_AGEMA_signal_14799 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6781 ( .C ( clk ), .D ( new_AGEMA_signal_14808 ), .Q ( new_AGEMA_signal_14809 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6791 ( .C ( clk ), .D ( new_AGEMA_signal_14818 ), .Q ( new_AGEMA_signal_14819 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6815 ( .C ( clk ), .D ( n2829 ), .Q ( new_AGEMA_signal_14843 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6823 ( .C ( clk ), .D ( new_AGEMA_signal_3420 ), .Q ( new_AGEMA_signal_14851 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6831 ( .C ( clk ), .D ( new_AGEMA_signal_3421 ), .Q ( new_AGEMA_signal_14859 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6839 ( .C ( clk ), .D ( new_AGEMA_signal_3422 ), .Q ( new_AGEMA_signal_14867 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6901 ( .C ( clk ), .D ( new_AGEMA_signal_14928 ), .Q ( new_AGEMA_signal_14929 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6917 ( .C ( clk ), .D ( new_AGEMA_signal_14944 ), .Q ( new_AGEMA_signal_14945 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6933 ( .C ( clk ), .D ( new_AGEMA_signal_14960 ), .Q ( new_AGEMA_signal_14961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6949 ( .C ( clk ), .D ( new_AGEMA_signal_14976 ), .Q ( new_AGEMA_signal_14977 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6959 ( .C ( clk ), .D ( n2312 ), .Q ( new_AGEMA_signal_14987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6969 ( .C ( clk ), .D ( new_AGEMA_signal_3342 ), .Q ( new_AGEMA_signal_14997 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6979 ( .C ( clk ), .D ( new_AGEMA_signal_3343 ), .Q ( new_AGEMA_signal_15007 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6989 ( .C ( clk ), .D ( new_AGEMA_signal_3344 ), .Q ( new_AGEMA_signal_15017 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7007 ( .C ( clk ), .D ( new_AGEMA_signal_15034 ), .Q ( new_AGEMA_signal_15035 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7025 ( .C ( clk ), .D ( new_AGEMA_signal_15052 ), .Q ( new_AGEMA_signal_15053 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7043 ( .C ( clk ), .D ( new_AGEMA_signal_15070 ), .Q ( new_AGEMA_signal_15071 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7061 ( .C ( clk ), .D ( new_AGEMA_signal_15088 ), .Q ( new_AGEMA_signal_15089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7207 ( .C ( clk ), .D ( new_AGEMA_signal_15234 ), .Q ( new_AGEMA_signal_15235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7227 ( .C ( clk ), .D ( new_AGEMA_signal_15254 ), .Q ( new_AGEMA_signal_15255 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7247 ( .C ( clk ), .D ( new_AGEMA_signal_15274 ), .Q ( new_AGEMA_signal_15275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7267 ( .C ( clk ), .D ( new_AGEMA_signal_15294 ), .Q ( new_AGEMA_signal_15295 ) ) ;

    /* cells in depth 16 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2003 ( .a ({new_AGEMA_signal_12778, new_AGEMA_signal_12772, new_AGEMA_signal_12766, new_AGEMA_signal_12760}), .b ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, n1935}), .clk ( clk ), .r ({Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, n1941}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2059 ( .a ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, new_AGEMA_signal_3297, n1959}), .b ({new_AGEMA_signal_12786, new_AGEMA_signal_12784, new_AGEMA_signal_12782, new_AGEMA_signal_12780}), .clk ( clk ), .r ({Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590]}), .c ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n1960}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2110 ( .a ({new_AGEMA_signal_12802, new_AGEMA_signal_12798, new_AGEMA_signal_12794, new_AGEMA_signal_12790}), .b ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, n1983}), .clk ( clk ), .r ({Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, n1988}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2153 ( .a ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, new_AGEMA_signal_3303, n2014}), .b ({new_AGEMA_signal_12834, new_AGEMA_signal_12826, new_AGEMA_signal_12818, new_AGEMA_signal_12810}), .clk ( clk ), .r ({Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602]}), .c ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, n2015}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2169 ( .a ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, n2029}), .b ({new_AGEMA_signal_12866, new_AGEMA_signal_12858, new_AGEMA_signal_12850, new_AGEMA_signal_12842}), .clk ( clk ), .r ({Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608]}), .c ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2030}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2200 ( .a ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, n2052}), .b ({new_AGEMA_signal_12898, new_AGEMA_signal_12890, new_AGEMA_signal_12882, new_AGEMA_signal_12874}), .clk ( clk ), .r ({Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614]}), .c ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2053}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2222 ( .a ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, n2070}), .b ({new_AGEMA_signal_12930, new_AGEMA_signal_12922, new_AGEMA_signal_12914, new_AGEMA_signal_12906}), .clk ( clk ), .r ({Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620]}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, new_AGEMA_signal_3441, n2071}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2259 ( .a ({new_AGEMA_signal_12954, new_AGEMA_signal_12948, new_AGEMA_signal_12942, new_AGEMA_signal_12936}), .b ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, n2098}), .clk ( clk ), .r ({Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626]}), .c ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, n2103}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2288 ( .a ({new_AGEMA_signal_12994, new_AGEMA_signal_12984, new_AGEMA_signal_12974, new_AGEMA_signal_12964}), .b ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, n2125}), .clk ( clk ), .r ({Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, n2126}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2314 ( .a ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, n2145}), .b ({new_AGEMA_signal_13026, new_AGEMA_signal_13018, new_AGEMA_signal_13010, new_AGEMA_signal_13002}), .clk ( clk ), .r ({Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638]}), .c ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2146}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2334 ( .a ({new_AGEMA_signal_13058, new_AGEMA_signal_13050, new_AGEMA_signal_13042, new_AGEMA_signal_13034}), .b ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, n2169}), .clk ( clk ), .r ({Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644]}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3453, n2173}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2351 ( .a ({new_AGEMA_signal_13090, new_AGEMA_signal_13082, new_AGEMA_signal_13074, new_AGEMA_signal_13066}), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, n2185}), .clk ( clk ), .r ({Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650]}), .c ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, n2187}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2416 ( .a ({new_AGEMA_signal_13098, new_AGEMA_signal_13096, new_AGEMA_signal_13094, new_AGEMA_signal_13092}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, n2251}), .clk ( clk ), .r ({Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656]}), .c ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2256}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2441 ( .a ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, n2274}), .b ({new_AGEMA_signal_13114, new_AGEMA_signal_13110, new_AGEMA_signal_13106, new_AGEMA_signal_13102}), .clk ( clk ), .r ({Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662]}), .c ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, new_AGEMA_signal_3465, n2275}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2474 ( .a ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, n2302}), .b ({new_AGEMA_signal_13138, new_AGEMA_signal_13132, new_AGEMA_signal_13126, new_AGEMA_signal_13120}), .clk ( clk ), .r ({Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668]}), .c ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, n2303}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2504 ( .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, n2339}), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, n2338}), .clk ( clk ), .r ({Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674]}), .c ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, new_AGEMA_signal_3471, n2382}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2516 ( .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, n2351}), .b ({new_AGEMA_signal_13154, new_AGEMA_signal_13150, new_AGEMA_signal_13146, new_AGEMA_signal_13142}), .clk ( clk ), .r ({Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680]}), .c ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, n2380}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2531 ( .a ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, n2365}), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13184, new_AGEMA_signal_13174, new_AGEMA_signal_13164}), .clk ( clk ), .r ({Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686]}), .c ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477, n2366}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2561 ( .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, n2399}), .b ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, n2398}), .clk ( clk ), .r ({Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692]}), .c ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, n2425}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2582 ( .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, n2423}), .b ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, n2422}), .clk ( clk ), .r ({Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698]}), .c ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, n2424}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2597 ( .a ({new_AGEMA_signal_13226, new_AGEMA_signal_13218, new_AGEMA_signal_13210, new_AGEMA_signal_13202}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, n2441}), .clk ( clk ), .r ({Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704]}), .c ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, n2451}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2631 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, n2479}), .b ({new_AGEMA_signal_13242, new_AGEMA_signal_13238, new_AGEMA_signal_13234, new_AGEMA_signal_13230}), .clk ( clk ), .r ({Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710]}), .c ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, n2514}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2658 ( .a ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, n2510}), .b ({new_AGEMA_signal_13250, new_AGEMA_signal_13248, new_AGEMA_signal_13246, new_AGEMA_signal_13244}), .clk ( clk ), .r ({Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716]}), .c ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2511}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2688 ( .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, n2552}), .b ({new_AGEMA_signal_13282, new_AGEMA_signal_13274, new_AGEMA_signal_13266, new_AGEMA_signal_13258}), .clk ( clk ), .r ({Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722]}), .c ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, new_AGEMA_signal_3489, n2671}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2716 ( .a ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, n2589}), .b ({new_AGEMA_signal_13314, new_AGEMA_signal_13306, new_AGEMA_signal_13298, new_AGEMA_signal_13290}), .clk ( clk ), .r ({Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728]}), .c ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, n2590}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2731 ( .a ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, n2608}), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13332, new_AGEMA_signal_13326, new_AGEMA_signal_13320}), .clk ( clk ), .r ({Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734]}), .c ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2623}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2763 ( .a ({new_AGEMA_signal_13354, new_AGEMA_signal_13350, new_AGEMA_signal_13346, new_AGEMA_signal_13342}), .b ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, n2659}), .clk ( clk ), .r ({Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740]}), .c ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2667}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2786 ( .a ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, n2702}), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13378, new_AGEMA_signal_13370, new_AGEMA_signal_13362}), .clk ( clk ), .r ({Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746]}), .c ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501, n2703}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) U2840 ( .s ({new_AGEMA_signal_13114, new_AGEMA_signal_13110, new_AGEMA_signal_13106, new_AGEMA_signal_13102}), .b ({new_AGEMA_signal_13394, new_AGEMA_signal_13392, new_AGEMA_signal_13390, new_AGEMA_signal_13388}), .a ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, n2801}), .clk ( clk ), .r ({Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752]}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, n2803}) ) ;
    buf_clk new_AGEMA_reg_buffer_5372 ( .C ( clk ), .D ( new_AGEMA_signal_13399 ), .Q ( new_AGEMA_signal_13400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5378 ( .C ( clk ), .D ( new_AGEMA_signal_13405 ), .Q ( new_AGEMA_signal_13406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5384 ( .C ( clk ), .D ( new_AGEMA_signal_13411 ), .Q ( new_AGEMA_signal_13412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5390 ( .C ( clk ), .D ( new_AGEMA_signal_13417 ), .Q ( new_AGEMA_signal_13418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5396 ( .C ( clk ), .D ( new_AGEMA_signal_13423 ), .Q ( new_AGEMA_signal_13424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5402 ( .C ( clk ), .D ( new_AGEMA_signal_13429 ), .Q ( new_AGEMA_signal_13430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5408 ( .C ( clk ), .D ( new_AGEMA_signal_13435 ), .Q ( new_AGEMA_signal_13436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5414 ( .C ( clk ), .D ( new_AGEMA_signal_13441 ), .Q ( new_AGEMA_signal_13442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5420 ( .C ( clk ), .D ( new_AGEMA_signal_13447 ), .Q ( new_AGEMA_signal_13448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5426 ( .C ( clk ), .D ( new_AGEMA_signal_13453 ), .Q ( new_AGEMA_signal_13454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5432 ( .C ( clk ), .D ( new_AGEMA_signal_13459 ), .Q ( new_AGEMA_signal_13460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5438 ( .C ( clk ), .D ( new_AGEMA_signal_13465 ), .Q ( new_AGEMA_signal_13466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5442 ( .C ( clk ), .D ( new_AGEMA_signal_13469 ), .Q ( new_AGEMA_signal_13470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5446 ( .C ( clk ), .D ( new_AGEMA_signal_13473 ), .Q ( new_AGEMA_signal_13474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5450 ( .C ( clk ), .D ( new_AGEMA_signal_13477 ), .Q ( new_AGEMA_signal_13478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5454 ( .C ( clk ), .D ( new_AGEMA_signal_13481 ), .Q ( new_AGEMA_signal_13482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5462 ( .C ( clk ), .D ( new_AGEMA_signal_13489 ), .Q ( new_AGEMA_signal_13490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5470 ( .C ( clk ), .D ( new_AGEMA_signal_13497 ), .Q ( new_AGEMA_signal_13498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5478 ( .C ( clk ), .D ( new_AGEMA_signal_13505 ), .Q ( new_AGEMA_signal_13506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5486 ( .C ( clk ), .D ( new_AGEMA_signal_13513 ), .Q ( new_AGEMA_signal_13514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5492 ( .C ( clk ), .D ( new_AGEMA_signal_13519 ), .Q ( new_AGEMA_signal_13520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5498 ( .C ( clk ), .D ( new_AGEMA_signal_13525 ), .Q ( new_AGEMA_signal_13526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5504 ( .C ( clk ), .D ( new_AGEMA_signal_13531 ), .Q ( new_AGEMA_signal_13532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5510 ( .C ( clk ), .D ( new_AGEMA_signal_13537 ), .Q ( new_AGEMA_signal_13538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5514 ( .C ( clk ), .D ( new_AGEMA_signal_13541 ), .Q ( new_AGEMA_signal_13542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5518 ( .C ( clk ), .D ( new_AGEMA_signal_13545 ), .Q ( new_AGEMA_signal_13546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5522 ( .C ( clk ), .D ( new_AGEMA_signal_13549 ), .Q ( new_AGEMA_signal_13550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5526 ( .C ( clk ), .D ( new_AGEMA_signal_13553 ), .Q ( new_AGEMA_signal_13554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5534 ( .C ( clk ), .D ( new_AGEMA_signal_13561 ), .Q ( new_AGEMA_signal_13562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5542 ( .C ( clk ), .D ( new_AGEMA_signal_13569 ), .Q ( new_AGEMA_signal_13570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5550 ( .C ( clk ), .D ( new_AGEMA_signal_13577 ), .Q ( new_AGEMA_signal_13578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5558 ( .C ( clk ), .D ( new_AGEMA_signal_13585 ), .Q ( new_AGEMA_signal_13586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5566 ( .C ( clk ), .D ( new_AGEMA_signal_13593 ), .Q ( new_AGEMA_signal_13594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5574 ( .C ( clk ), .D ( new_AGEMA_signal_13601 ), .Q ( new_AGEMA_signal_13602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5582 ( .C ( clk ), .D ( new_AGEMA_signal_13609 ), .Q ( new_AGEMA_signal_13610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5590 ( .C ( clk ), .D ( new_AGEMA_signal_13617 ), .Q ( new_AGEMA_signal_13618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5600 ( .C ( clk ), .D ( new_AGEMA_signal_13627 ), .Q ( new_AGEMA_signal_13628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5610 ( .C ( clk ), .D ( new_AGEMA_signal_13637 ), .Q ( new_AGEMA_signal_13638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5620 ( .C ( clk ), .D ( new_AGEMA_signal_13647 ), .Q ( new_AGEMA_signal_13648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5630 ( .C ( clk ), .D ( new_AGEMA_signal_13657 ), .Q ( new_AGEMA_signal_13658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5638 ( .C ( clk ), .D ( new_AGEMA_signal_13665 ), .Q ( new_AGEMA_signal_13666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5646 ( .C ( clk ), .D ( new_AGEMA_signal_13673 ), .Q ( new_AGEMA_signal_13674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5654 ( .C ( clk ), .D ( new_AGEMA_signal_13681 ), .Q ( new_AGEMA_signal_13682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5662 ( .C ( clk ), .D ( new_AGEMA_signal_13689 ), .Q ( new_AGEMA_signal_13690 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5668 ( .C ( clk ), .D ( new_AGEMA_signal_13695 ), .Q ( new_AGEMA_signal_13696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5674 ( .C ( clk ), .D ( new_AGEMA_signal_13701 ), .Q ( new_AGEMA_signal_13702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5680 ( .C ( clk ), .D ( new_AGEMA_signal_13707 ), .Q ( new_AGEMA_signal_13708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5686 ( .C ( clk ), .D ( new_AGEMA_signal_13713 ), .Q ( new_AGEMA_signal_13714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5690 ( .C ( clk ), .D ( new_AGEMA_signal_13717 ), .Q ( new_AGEMA_signal_13718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5694 ( .C ( clk ), .D ( new_AGEMA_signal_13721 ), .Q ( new_AGEMA_signal_13722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5698 ( .C ( clk ), .D ( new_AGEMA_signal_13725 ), .Q ( new_AGEMA_signal_13726 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5702 ( .C ( clk ), .D ( new_AGEMA_signal_13729 ), .Q ( new_AGEMA_signal_13730 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5708 ( .C ( clk ), .D ( new_AGEMA_signal_13735 ), .Q ( new_AGEMA_signal_13736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5714 ( .C ( clk ), .D ( new_AGEMA_signal_13741 ), .Q ( new_AGEMA_signal_13742 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5720 ( .C ( clk ), .D ( new_AGEMA_signal_13747 ), .Q ( new_AGEMA_signal_13748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5726 ( .C ( clk ), .D ( new_AGEMA_signal_13753 ), .Q ( new_AGEMA_signal_13754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5734 ( .C ( clk ), .D ( new_AGEMA_signal_13761 ), .Q ( new_AGEMA_signal_13762 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5742 ( .C ( clk ), .D ( new_AGEMA_signal_13769 ), .Q ( new_AGEMA_signal_13770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5750 ( .C ( clk ), .D ( new_AGEMA_signal_13777 ), .Q ( new_AGEMA_signal_13778 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5758 ( .C ( clk ), .D ( new_AGEMA_signal_13785 ), .Q ( new_AGEMA_signal_13786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5764 ( .C ( clk ), .D ( new_AGEMA_signal_13791 ), .Q ( new_AGEMA_signal_13792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5770 ( .C ( clk ), .D ( new_AGEMA_signal_13797 ), .Q ( new_AGEMA_signal_13798 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5776 ( .C ( clk ), .D ( new_AGEMA_signal_13803 ), .Q ( new_AGEMA_signal_13804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5782 ( .C ( clk ), .D ( new_AGEMA_signal_13809 ), .Q ( new_AGEMA_signal_13810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5784 ( .C ( clk ), .D ( new_AGEMA_signal_13811 ), .Q ( new_AGEMA_signal_13812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5786 ( .C ( clk ), .D ( new_AGEMA_signal_13813 ), .Q ( new_AGEMA_signal_13814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5788 ( .C ( clk ), .D ( new_AGEMA_signal_13815 ), .Q ( new_AGEMA_signal_13816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5790 ( .C ( clk ), .D ( new_AGEMA_signal_13817 ), .Q ( new_AGEMA_signal_13818 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5798 ( .C ( clk ), .D ( new_AGEMA_signal_13825 ), .Q ( new_AGEMA_signal_13826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5806 ( .C ( clk ), .D ( new_AGEMA_signal_13833 ), .Q ( new_AGEMA_signal_13834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5814 ( .C ( clk ), .D ( new_AGEMA_signal_13841 ), .Q ( new_AGEMA_signal_13842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5822 ( .C ( clk ), .D ( new_AGEMA_signal_13849 ), .Q ( new_AGEMA_signal_13850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5826 ( .C ( clk ), .D ( new_AGEMA_signal_13853 ), .Q ( new_AGEMA_signal_13854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5830 ( .C ( clk ), .D ( new_AGEMA_signal_13857 ), .Q ( new_AGEMA_signal_13858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5834 ( .C ( clk ), .D ( new_AGEMA_signal_13861 ), .Q ( new_AGEMA_signal_13862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5838 ( .C ( clk ), .D ( new_AGEMA_signal_13865 ), .Q ( new_AGEMA_signal_13866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5844 ( .C ( clk ), .D ( new_AGEMA_signal_13871 ), .Q ( new_AGEMA_signal_13872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5850 ( .C ( clk ), .D ( new_AGEMA_signal_13877 ), .Q ( new_AGEMA_signal_13878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5856 ( .C ( clk ), .D ( new_AGEMA_signal_13883 ), .Q ( new_AGEMA_signal_13884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5862 ( .C ( clk ), .D ( new_AGEMA_signal_13889 ), .Q ( new_AGEMA_signal_13890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5868 ( .C ( clk ), .D ( new_AGEMA_signal_13895 ), .Q ( new_AGEMA_signal_13896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5874 ( .C ( clk ), .D ( new_AGEMA_signal_13901 ), .Q ( new_AGEMA_signal_13902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5880 ( .C ( clk ), .D ( new_AGEMA_signal_13907 ), .Q ( new_AGEMA_signal_13908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5886 ( .C ( clk ), .D ( new_AGEMA_signal_13913 ), .Q ( new_AGEMA_signal_13914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5890 ( .C ( clk ), .D ( new_AGEMA_signal_13917 ), .Q ( new_AGEMA_signal_13918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5894 ( .C ( clk ), .D ( new_AGEMA_signal_13921 ), .Q ( new_AGEMA_signal_13922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5898 ( .C ( clk ), .D ( new_AGEMA_signal_13925 ), .Q ( new_AGEMA_signal_13926 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5902 ( .C ( clk ), .D ( new_AGEMA_signal_13929 ), .Q ( new_AGEMA_signal_13930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5906 ( .C ( clk ), .D ( new_AGEMA_signal_13933 ), .Q ( new_AGEMA_signal_13934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5912 ( .C ( clk ), .D ( new_AGEMA_signal_13939 ), .Q ( new_AGEMA_signal_13940 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5918 ( .C ( clk ), .D ( new_AGEMA_signal_13945 ), .Q ( new_AGEMA_signal_13946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5924 ( .C ( clk ), .D ( new_AGEMA_signal_13951 ), .Q ( new_AGEMA_signal_13952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5928 ( .C ( clk ), .D ( new_AGEMA_signal_13955 ), .Q ( new_AGEMA_signal_13956 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5932 ( .C ( clk ), .D ( new_AGEMA_signal_13959 ), .Q ( new_AGEMA_signal_13960 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5936 ( .C ( clk ), .D ( new_AGEMA_signal_13963 ), .Q ( new_AGEMA_signal_13964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5940 ( .C ( clk ), .D ( new_AGEMA_signal_13967 ), .Q ( new_AGEMA_signal_13968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5946 ( .C ( clk ), .D ( new_AGEMA_signal_13973 ), .Q ( new_AGEMA_signal_13974 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5952 ( .C ( clk ), .D ( new_AGEMA_signal_13979 ), .Q ( new_AGEMA_signal_13980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5958 ( .C ( clk ), .D ( new_AGEMA_signal_13985 ), .Q ( new_AGEMA_signal_13986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5964 ( .C ( clk ), .D ( new_AGEMA_signal_13991 ), .Q ( new_AGEMA_signal_13992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5974 ( .C ( clk ), .D ( new_AGEMA_signal_14001 ), .Q ( new_AGEMA_signal_14002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5984 ( .C ( clk ), .D ( new_AGEMA_signal_14011 ), .Q ( new_AGEMA_signal_14012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5994 ( .C ( clk ), .D ( new_AGEMA_signal_14021 ), .Q ( new_AGEMA_signal_14022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6004 ( .C ( clk ), .D ( new_AGEMA_signal_14031 ), .Q ( new_AGEMA_signal_14032 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6010 ( .C ( clk ), .D ( new_AGEMA_signal_14037 ), .Q ( new_AGEMA_signal_14038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6016 ( .C ( clk ), .D ( new_AGEMA_signal_14043 ), .Q ( new_AGEMA_signal_14044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C ( clk ), .D ( new_AGEMA_signal_14049 ), .Q ( new_AGEMA_signal_14050 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C ( clk ), .D ( new_AGEMA_signal_14055 ), .Q ( new_AGEMA_signal_14056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C ( clk ), .D ( new_AGEMA_signal_14061 ), .Q ( new_AGEMA_signal_14062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C ( clk ), .D ( new_AGEMA_signal_14067 ), .Q ( new_AGEMA_signal_14068 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C ( clk ), .D ( new_AGEMA_signal_14073 ), .Q ( new_AGEMA_signal_14074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6052 ( .C ( clk ), .D ( new_AGEMA_signal_14079 ), .Q ( new_AGEMA_signal_14080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6056 ( .C ( clk ), .D ( new_AGEMA_signal_14083 ), .Q ( new_AGEMA_signal_14084 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6060 ( .C ( clk ), .D ( new_AGEMA_signal_14087 ), .Q ( new_AGEMA_signal_14088 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6064 ( .C ( clk ), .D ( new_AGEMA_signal_14091 ), .Q ( new_AGEMA_signal_14092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6068 ( .C ( clk ), .D ( new_AGEMA_signal_14095 ), .Q ( new_AGEMA_signal_14096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6072 ( .C ( clk ), .D ( new_AGEMA_signal_14099 ), .Q ( new_AGEMA_signal_14100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6076 ( .C ( clk ), .D ( new_AGEMA_signal_14103 ), .Q ( new_AGEMA_signal_14104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6080 ( .C ( clk ), .D ( new_AGEMA_signal_14107 ), .Q ( new_AGEMA_signal_14108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6084 ( .C ( clk ), .D ( new_AGEMA_signal_14111 ), .Q ( new_AGEMA_signal_14112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6092 ( .C ( clk ), .D ( new_AGEMA_signal_14119 ), .Q ( new_AGEMA_signal_14120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6100 ( .C ( clk ), .D ( new_AGEMA_signal_14127 ), .Q ( new_AGEMA_signal_14128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6108 ( .C ( clk ), .D ( new_AGEMA_signal_14135 ), .Q ( new_AGEMA_signal_14136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6116 ( .C ( clk ), .D ( new_AGEMA_signal_14143 ), .Q ( new_AGEMA_signal_14144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6122 ( .C ( clk ), .D ( new_AGEMA_signal_14149 ), .Q ( new_AGEMA_signal_14150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6128 ( .C ( clk ), .D ( new_AGEMA_signal_14155 ), .Q ( new_AGEMA_signal_14156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6134 ( .C ( clk ), .D ( new_AGEMA_signal_14161 ), .Q ( new_AGEMA_signal_14162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6140 ( .C ( clk ), .D ( new_AGEMA_signal_14167 ), .Q ( new_AGEMA_signal_14168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6148 ( .C ( clk ), .D ( new_AGEMA_signal_14175 ), .Q ( new_AGEMA_signal_14176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6156 ( .C ( clk ), .D ( new_AGEMA_signal_14183 ), .Q ( new_AGEMA_signal_14184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6164 ( .C ( clk ), .D ( new_AGEMA_signal_14191 ), .Q ( new_AGEMA_signal_14192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6172 ( .C ( clk ), .D ( new_AGEMA_signal_14199 ), .Q ( new_AGEMA_signal_14200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6180 ( .C ( clk ), .D ( new_AGEMA_signal_14207 ), .Q ( new_AGEMA_signal_14208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6188 ( .C ( clk ), .D ( new_AGEMA_signal_14215 ), .Q ( new_AGEMA_signal_14216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6196 ( .C ( clk ), .D ( new_AGEMA_signal_14223 ), .Q ( new_AGEMA_signal_14224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6204 ( .C ( clk ), .D ( new_AGEMA_signal_14231 ), .Q ( new_AGEMA_signal_14232 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6216 ( .C ( clk ), .D ( new_AGEMA_signal_14243 ), .Q ( new_AGEMA_signal_14244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6220 ( .C ( clk ), .D ( new_AGEMA_signal_14247 ), .Q ( new_AGEMA_signal_14248 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6224 ( .C ( clk ), .D ( new_AGEMA_signal_14251 ), .Q ( new_AGEMA_signal_14252 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6228 ( .C ( clk ), .D ( new_AGEMA_signal_14255 ), .Q ( new_AGEMA_signal_14256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6232 ( .C ( clk ), .D ( new_AGEMA_signal_14259 ), .Q ( new_AGEMA_signal_14260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6236 ( .C ( clk ), .D ( new_AGEMA_signal_14263 ), .Q ( new_AGEMA_signal_14264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6240 ( .C ( clk ), .D ( new_AGEMA_signal_14267 ), .Q ( new_AGEMA_signal_14268 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6244 ( .C ( clk ), .D ( new_AGEMA_signal_14271 ), .Q ( new_AGEMA_signal_14272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6252 ( .C ( clk ), .D ( new_AGEMA_signal_14279 ), .Q ( new_AGEMA_signal_14280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6260 ( .C ( clk ), .D ( new_AGEMA_signal_14287 ), .Q ( new_AGEMA_signal_14288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6268 ( .C ( clk ), .D ( new_AGEMA_signal_14295 ), .Q ( new_AGEMA_signal_14296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6276 ( .C ( clk ), .D ( new_AGEMA_signal_14303 ), .Q ( new_AGEMA_signal_14304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6280 ( .C ( clk ), .D ( new_AGEMA_signal_14307 ), .Q ( new_AGEMA_signal_14308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6284 ( .C ( clk ), .D ( new_AGEMA_signal_14311 ), .Q ( new_AGEMA_signal_14312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6288 ( .C ( clk ), .D ( new_AGEMA_signal_14315 ), .Q ( new_AGEMA_signal_14316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6292 ( .C ( clk ), .D ( new_AGEMA_signal_14319 ), .Q ( new_AGEMA_signal_14320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6298 ( .C ( clk ), .D ( new_AGEMA_signal_14325 ), .Q ( new_AGEMA_signal_14326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6306 ( .C ( clk ), .D ( new_AGEMA_signal_14333 ), .Q ( new_AGEMA_signal_14334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6314 ( .C ( clk ), .D ( new_AGEMA_signal_14341 ), .Q ( new_AGEMA_signal_14342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6322 ( .C ( clk ), .D ( new_AGEMA_signal_14349 ), .Q ( new_AGEMA_signal_14350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6334 ( .C ( clk ), .D ( new_AGEMA_signal_14361 ), .Q ( new_AGEMA_signal_14362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6346 ( .C ( clk ), .D ( new_AGEMA_signal_14373 ), .Q ( new_AGEMA_signal_14374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6358 ( .C ( clk ), .D ( new_AGEMA_signal_14385 ), .Q ( new_AGEMA_signal_14386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6370 ( .C ( clk ), .D ( new_AGEMA_signal_14397 ), .Q ( new_AGEMA_signal_14398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6384 ( .C ( clk ), .D ( new_AGEMA_signal_14411 ), .Q ( new_AGEMA_signal_14412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6398 ( .C ( clk ), .D ( new_AGEMA_signal_14425 ), .Q ( new_AGEMA_signal_14426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6412 ( .C ( clk ), .D ( new_AGEMA_signal_14439 ), .Q ( new_AGEMA_signal_14440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6426 ( .C ( clk ), .D ( new_AGEMA_signal_14453 ), .Q ( new_AGEMA_signal_14454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6434 ( .C ( clk ), .D ( new_AGEMA_signal_14461 ), .Q ( new_AGEMA_signal_14462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6442 ( .C ( clk ), .D ( new_AGEMA_signal_14469 ), .Q ( new_AGEMA_signal_14470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6450 ( .C ( clk ), .D ( new_AGEMA_signal_14477 ), .Q ( new_AGEMA_signal_14478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6458 ( .C ( clk ), .D ( new_AGEMA_signal_14485 ), .Q ( new_AGEMA_signal_14486 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6472 ( .C ( clk ), .D ( new_AGEMA_signal_14499 ), .Q ( new_AGEMA_signal_14500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6486 ( .C ( clk ), .D ( new_AGEMA_signal_14513 ), .Q ( new_AGEMA_signal_14514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6500 ( .C ( clk ), .D ( new_AGEMA_signal_14527 ), .Q ( new_AGEMA_signal_14528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6514 ( .C ( clk ), .D ( new_AGEMA_signal_14541 ), .Q ( new_AGEMA_signal_14542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6522 ( .C ( clk ), .D ( new_AGEMA_signal_14549 ), .Q ( new_AGEMA_signal_14550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6530 ( .C ( clk ), .D ( new_AGEMA_signal_14557 ), .Q ( new_AGEMA_signal_14558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6538 ( .C ( clk ), .D ( new_AGEMA_signal_14565 ), .Q ( new_AGEMA_signal_14566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6546 ( .C ( clk ), .D ( new_AGEMA_signal_14573 ), .Q ( new_AGEMA_signal_14574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6554 ( .C ( clk ), .D ( new_AGEMA_signal_14581 ), .Q ( new_AGEMA_signal_14582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6562 ( .C ( clk ), .D ( new_AGEMA_signal_14589 ), .Q ( new_AGEMA_signal_14590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6570 ( .C ( clk ), .D ( new_AGEMA_signal_14597 ), .Q ( new_AGEMA_signal_14598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6578 ( .C ( clk ), .D ( new_AGEMA_signal_14605 ), .Q ( new_AGEMA_signal_14606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6616 ( .C ( clk ), .D ( new_AGEMA_signal_14643 ), .Q ( new_AGEMA_signal_14644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6632 ( .C ( clk ), .D ( new_AGEMA_signal_14659 ), .Q ( new_AGEMA_signal_14660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6648 ( .C ( clk ), .D ( new_AGEMA_signal_14675 ), .Q ( new_AGEMA_signal_14676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6664 ( .C ( clk ), .D ( new_AGEMA_signal_14691 ), .Q ( new_AGEMA_signal_14692 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6704 ( .C ( clk ), .D ( new_AGEMA_signal_14731 ), .Q ( new_AGEMA_signal_14732 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6720 ( .C ( clk ), .D ( new_AGEMA_signal_14747 ), .Q ( new_AGEMA_signal_14748 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6736 ( .C ( clk ), .D ( new_AGEMA_signal_14763 ), .Q ( new_AGEMA_signal_14764 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6752 ( .C ( clk ), .D ( new_AGEMA_signal_14779 ), .Q ( new_AGEMA_signal_14780 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6762 ( .C ( clk ), .D ( new_AGEMA_signal_14789 ), .Q ( new_AGEMA_signal_14790 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6772 ( .C ( clk ), .D ( new_AGEMA_signal_14799 ), .Q ( new_AGEMA_signal_14800 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6782 ( .C ( clk ), .D ( new_AGEMA_signal_14809 ), .Q ( new_AGEMA_signal_14810 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6792 ( .C ( clk ), .D ( new_AGEMA_signal_14819 ), .Q ( new_AGEMA_signal_14820 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6816 ( .C ( clk ), .D ( new_AGEMA_signal_14843 ), .Q ( new_AGEMA_signal_14844 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6824 ( .C ( clk ), .D ( new_AGEMA_signal_14851 ), .Q ( new_AGEMA_signal_14852 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6832 ( .C ( clk ), .D ( new_AGEMA_signal_14859 ), .Q ( new_AGEMA_signal_14860 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6840 ( .C ( clk ), .D ( new_AGEMA_signal_14867 ), .Q ( new_AGEMA_signal_14868 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6902 ( .C ( clk ), .D ( new_AGEMA_signal_14929 ), .Q ( new_AGEMA_signal_14930 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6918 ( .C ( clk ), .D ( new_AGEMA_signal_14945 ), .Q ( new_AGEMA_signal_14946 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6934 ( .C ( clk ), .D ( new_AGEMA_signal_14961 ), .Q ( new_AGEMA_signal_14962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6950 ( .C ( clk ), .D ( new_AGEMA_signal_14977 ), .Q ( new_AGEMA_signal_14978 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6960 ( .C ( clk ), .D ( new_AGEMA_signal_14987 ), .Q ( new_AGEMA_signal_14988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6970 ( .C ( clk ), .D ( new_AGEMA_signal_14997 ), .Q ( new_AGEMA_signal_14998 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6980 ( .C ( clk ), .D ( new_AGEMA_signal_15007 ), .Q ( new_AGEMA_signal_15008 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6990 ( .C ( clk ), .D ( new_AGEMA_signal_15017 ), .Q ( new_AGEMA_signal_15018 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7008 ( .C ( clk ), .D ( new_AGEMA_signal_15035 ), .Q ( new_AGEMA_signal_15036 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7026 ( .C ( clk ), .D ( new_AGEMA_signal_15053 ), .Q ( new_AGEMA_signal_15054 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7044 ( .C ( clk ), .D ( new_AGEMA_signal_15071 ), .Q ( new_AGEMA_signal_15072 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7062 ( .C ( clk ), .D ( new_AGEMA_signal_15089 ), .Q ( new_AGEMA_signal_15090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7208 ( .C ( clk ), .D ( new_AGEMA_signal_15235 ), .Q ( new_AGEMA_signal_15236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7228 ( .C ( clk ), .D ( new_AGEMA_signal_15255 ), .Q ( new_AGEMA_signal_15256 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7248 ( .C ( clk ), .D ( new_AGEMA_signal_15275 ), .Q ( new_AGEMA_signal_15276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7268 ( .C ( clk ), .D ( new_AGEMA_signal_15295 ), .Q ( new_AGEMA_signal_15296 ) ) ;

    /* cells in depth 17 */
    buf_clk new_AGEMA_reg_buffer_5907 ( .C ( clk ), .D ( new_AGEMA_signal_13934 ), .Q ( new_AGEMA_signal_13935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5913 ( .C ( clk ), .D ( new_AGEMA_signal_13940 ), .Q ( new_AGEMA_signal_13941 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5919 ( .C ( clk ), .D ( new_AGEMA_signal_13946 ), .Q ( new_AGEMA_signal_13947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5925 ( .C ( clk ), .D ( new_AGEMA_signal_13952 ), .Q ( new_AGEMA_signal_13953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5929 ( .C ( clk ), .D ( new_AGEMA_signal_13956 ), .Q ( new_AGEMA_signal_13957 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5933 ( .C ( clk ), .D ( new_AGEMA_signal_13960 ), .Q ( new_AGEMA_signal_13961 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5937 ( .C ( clk ), .D ( new_AGEMA_signal_13964 ), .Q ( new_AGEMA_signal_13965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5941 ( .C ( clk ), .D ( new_AGEMA_signal_13968 ), .Q ( new_AGEMA_signal_13969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5947 ( .C ( clk ), .D ( new_AGEMA_signal_13974 ), .Q ( new_AGEMA_signal_13975 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5953 ( .C ( clk ), .D ( new_AGEMA_signal_13980 ), .Q ( new_AGEMA_signal_13981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5959 ( .C ( clk ), .D ( new_AGEMA_signal_13986 ), .Q ( new_AGEMA_signal_13987 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5965 ( .C ( clk ), .D ( new_AGEMA_signal_13992 ), .Q ( new_AGEMA_signal_13993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5975 ( .C ( clk ), .D ( new_AGEMA_signal_14002 ), .Q ( new_AGEMA_signal_14003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5985 ( .C ( clk ), .D ( new_AGEMA_signal_14012 ), .Q ( new_AGEMA_signal_14013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5995 ( .C ( clk ), .D ( new_AGEMA_signal_14022 ), .Q ( new_AGEMA_signal_14023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6005 ( .C ( clk ), .D ( new_AGEMA_signal_14032 ), .Q ( new_AGEMA_signal_14033 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6011 ( .C ( clk ), .D ( new_AGEMA_signal_14038 ), .Q ( new_AGEMA_signal_14039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6017 ( .C ( clk ), .D ( new_AGEMA_signal_14044 ), .Q ( new_AGEMA_signal_14045 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C ( clk ), .D ( new_AGEMA_signal_14050 ), .Q ( new_AGEMA_signal_14051 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C ( clk ), .D ( new_AGEMA_signal_14056 ), .Q ( new_AGEMA_signal_14057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C ( clk ), .D ( new_AGEMA_signal_14062 ), .Q ( new_AGEMA_signal_14063 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C ( clk ), .D ( new_AGEMA_signal_14068 ), .Q ( new_AGEMA_signal_14069 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C ( clk ), .D ( new_AGEMA_signal_14074 ), .Q ( new_AGEMA_signal_14075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6053 ( .C ( clk ), .D ( new_AGEMA_signal_14080 ), .Q ( new_AGEMA_signal_14081 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6057 ( .C ( clk ), .D ( new_AGEMA_signal_14084 ), .Q ( new_AGEMA_signal_14085 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6061 ( .C ( clk ), .D ( new_AGEMA_signal_14088 ), .Q ( new_AGEMA_signal_14089 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6065 ( .C ( clk ), .D ( new_AGEMA_signal_14092 ), .Q ( new_AGEMA_signal_14093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6069 ( .C ( clk ), .D ( new_AGEMA_signal_14096 ), .Q ( new_AGEMA_signal_14097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6073 ( .C ( clk ), .D ( new_AGEMA_signal_14100 ), .Q ( new_AGEMA_signal_14101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6077 ( .C ( clk ), .D ( new_AGEMA_signal_14104 ), .Q ( new_AGEMA_signal_14105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6081 ( .C ( clk ), .D ( new_AGEMA_signal_14108 ), .Q ( new_AGEMA_signal_14109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6085 ( .C ( clk ), .D ( new_AGEMA_signal_14112 ), .Q ( new_AGEMA_signal_14113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6093 ( .C ( clk ), .D ( new_AGEMA_signal_14120 ), .Q ( new_AGEMA_signal_14121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6101 ( .C ( clk ), .D ( new_AGEMA_signal_14128 ), .Q ( new_AGEMA_signal_14129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6109 ( .C ( clk ), .D ( new_AGEMA_signal_14136 ), .Q ( new_AGEMA_signal_14137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6117 ( .C ( clk ), .D ( new_AGEMA_signal_14144 ), .Q ( new_AGEMA_signal_14145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6123 ( .C ( clk ), .D ( new_AGEMA_signal_14150 ), .Q ( new_AGEMA_signal_14151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6129 ( .C ( clk ), .D ( new_AGEMA_signal_14156 ), .Q ( new_AGEMA_signal_14157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6135 ( .C ( clk ), .D ( new_AGEMA_signal_14162 ), .Q ( new_AGEMA_signal_14163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6141 ( .C ( clk ), .D ( new_AGEMA_signal_14168 ), .Q ( new_AGEMA_signal_14169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6149 ( .C ( clk ), .D ( new_AGEMA_signal_14176 ), .Q ( new_AGEMA_signal_14177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6157 ( .C ( clk ), .D ( new_AGEMA_signal_14184 ), .Q ( new_AGEMA_signal_14185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6165 ( .C ( clk ), .D ( new_AGEMA_signal_14192 ), .Q ( new_AGEMA_signal_14193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6173 ( .C ( clk ), .D ( new_AGEMA_signal_14200 ), .Q ( new_AGEMA_signal_14201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6181 ( .C ( clk ), .D ( new_AGEMA_signal_14208 ), .Q ( new_AGEMA_signal_14209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6189 ( .C ( clk ), .D ( new_AGEMA_signal_14216 ), .Q ( new_AGEMA_signal_14217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6197 ( .C ( clk ), .D ( new_AGEMA_signal_14224 ), .Q ( new_AGEMA_signal_14225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6205 ( .C ( clk ), .D ( new_AGEMA_signal_14232 ), .Q ( new_AGEMA_signal_14233 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6207 ( .C ( clk ), .D ( n2514 ), .Q ( new_AGEMA_signal_14235 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6209 ( .C ( clk ), .D ( new_AGEMA_signal_3378 ), .Q ( new_AGEMA_signal_14237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6211 ( .C ( clk ), .D ( new_AGEMA_signal_3379 ), .Q ( new_AGEMA_signal_14239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6213 ( .C ( clk ), .D ( new_AGEMA_signal_3380 ), .Q ( new_AGEMA_signal_14241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6217 ( .C ( clk ), .D ( new_AGEMA_signal_14244 ), .Q ( new_AGEMA_signal_14245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6221 ( .C ( clk ), .D ( new_AGEMA_signal_14248 ), .Q ( new_AGEMA_signal_14249 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6225 ( .C ( clk ), .D ( new_AGEMA_signal_14252 ), .Q ( new_AGEMA_signal_14253 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6229 ( .C ( clk ), .D ( new_AGEMA_signal_14256 ), .Q ( new_AGEMA_signal_14257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6233 ( .C ( clk ), .D ( new_AGEMA_signal_14260 ), .Q ( new_AGEMA_signal_14261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6237 ( .C ( clk ), .D ( new_AGEMA_signal_14264 ), .Q ( new_AGEMA_signal_14265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6241 ( .C ( clk ), .D ( new_AGEMA_signal_14268 ), .Q ( new_AGEMA_signal_14269 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6245 ( .C ( clk ), .D ( new_AGEMA_signal_14272 ), .Q ( new_AGEMA_signal_14273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6253 ( .C ( clk ), .D ( new_AGEMA_signal_14280 ), .Q ( new_AGEMA_signal_14281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6261 ( .C ( clk ), .D ( new_AGEMA_signal_14288 ), .Q ( new_AGEMA_signal_14289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6269 ( .C ( clk ), .D ( new_AGEMA_signal_14296 ), .Q ( new_AGEMA_signal_14297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6277 ( .C ( clk ), .D ( new_AGEMA_signal_14304 ), .Q ( new_AGEMA_signal_14305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6281 ( .C ( clk ), .D ( new_AGEMA_signal_14308 ), .Q ( new_AGEMA_signal_14309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6285 ( .C ( clk ), .D ( new_AGEMA_signal_14312 ), .Q ( new_AGEMA_signal_14313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6289 ( .C ( clk ), .D ( new_AGEMA_signal_14316 ), .Q ( new_AGEMA_signal_14317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6293 ( .C ( clk ), .D ( new_AGEMA_signal_14320 ), .Q ( new_AGEMA_signal_14321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6299 ( .C ( clk ), .D ( new_AGEMA_signal_14326 ), .Q ( new_AGEMA_signal_14327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6307 ( .C ( clk ), .D ( new_AGEMA_signal_14334 ), .Q ( new_AGEMA_signal_14335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6315 ( .C ( clk ), .D ( new_AGEMA_signal_14342 ), .Q ( new_AGEMA_signal_14343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6323 ( .C ( clk ), .D ( new_AGEMA_signal_14350 ), .Q ( new_AGEMA_signal_14351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6335 ( .C ( clk ), .D ( new_AGEMA_signal_14362 ), .Q ( new_AGEMA_signal_14363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6347 ( .C ( clk ), .D ( new_AGEMA_signal_14374 ), .Q ( new_AGEMA_signal_14375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6359 ( .C ( clk ), .D ( new_AGEMA_signal_14386 ), .Q ( new_AGEMA_signal_14387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6371 ( .C ( clk ), .D ( new_AGEMA_signal_14398 ), .Q ( new_AGEMA_signal_14399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6385 ( .C ( clk ), .D ( new_AGEMA_signal_14412 ), .Q ( new_AGEMA_signal_14413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6399 ( .C ( clk ), .D ( new_AGEMA_signal_14426 ), .Q ( new_AGEMA_signal_14427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6413 ( .C ( clk ), .D ( new_AGEMA_signal_14440 ), .Q ( new_AGEMA_signal_14441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6427 ( .C ( clk ), .D ( new_AGEMA_signal_14454 ), .Q ( new_AGEMA_signal_14455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6435 ( .C ( clk ), .D ( new_AGEMA_signal_14462 ), .Q ( new_AGEMA_signal_14463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6443 ( .C ( clk ), .D ( new_AGEMA_signal_14470 ), .Q ( new_AGEMA_signal_14471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6451 ( .C ( clk ), .D ( new_AGEMA_signal_14478 ), .Q ( new_AGEMA_signal_14479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6459 ( .C ( clk ), .D ( new_AGEMA_signal_14486 ), .Q ( new_AGEMA_signal_14487 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6473 ( .C ( clk ), .D ( new_AGEMA_signal_14500 ), .Q ( new_AGEMA_signal_14501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6487 ( .C ( clk ), .D ( new_AGEMA_signal_14514 ), .Q ( new_AGEMA_signal_14515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6501 ( .C ( clk ), .D ( new_AGEMA_signal_14528 ), .Q ( new_AGEMA_signal_14529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6515 ( .C ( clk ), .D ( new_AGEMA_signal_14542 ), .Q ( new_AGEMA_signal_14543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6523 ( .C ( clk ), .D ( new_AGEMA_signal_14550 ), .Q ( new_AGEMA_signal_14551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6531 ( .C ( clk ), .D ( new_AGEMA_signal_14558 ), .Q ( new_AGEMA_signal_14559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6539 ( .C ( clk ), .D ( new_AGEMA_signal_14566 ), .Q ( new_AGEMA_signal_14567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6547 ( .C ( clk ), .D ( new_AGEMA_signal_14574 ), .Q ( new_AGEMA_signal_14575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6555 ( .C ( clk ), .D ( new_AGEMA_signal_14582 ), .Q ( new_AGEMA_signal_14583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6563 ( .C ( clk ), .D ( new_AGEMA_signal_14590 ), .Q ( new_AGEMA_signal_14591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6571 ( .C ( clk ), .D ( new_AGEMA_signal_14598 ), .Q ( new_AGEMA_signal_14599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6579 ( .C ( clk ), .D ( new_AGEMA_signal_14606 ), .Q ( new_AGEMA_signal_14607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6617 ( .C ( clk ), .D ( new_AGEMA_signal_14644 ), .Q ( new_AGEMA_signal_14645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6633 ( .C ( clk ), .D ( new_AGEMA_signal_14660 ), .Q ( new_AGEMA_signal_14661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6649 ( .C ( clk ), .D ( new_AGEMA_signal_14676 ), .Q ( new_AGEMA_signal_14677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6665 ( .C ( clk ), .D ( new_AGEMA_signal_14692 ), .Q ( new_AGEMA_signal_14693 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6705 ( .C ( clk ), .D ( new_AGEMA_signal_14732 ), .Q ( new_AGEMA_signal_14733 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6721 ( .C ( clk ), .D ( new_AGEMA_signal_14748 ), .Q ( new_AGEMA_signal_14749 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6737 ( .C ( clk ), .D ( new_AGEMA_signal_14764 ), .Q ( new_AGEMA_signal_14765 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6753 ( .C ( clk ), .D ( new_AGEMA_signal_14780 ), .Q ( new_AGEMA_signal_14781 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6763 ( .C ( clk ), .D ( new_AGEMA_signal_14790 ), .Q ( new_AGEMA_signal_14791 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6773 ( .C ( clk ), .D ( new_AGEMA_signal_14800 ), .Q ( new_AGEMA_signal_14801 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6783 ( .C ( clk ), .D ( new_AGEMA_signal_14810 ), .Q ( new_AGEMA_signal_14811 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6793 ( .C ( clk ), .D ( new_AGEMA_signal_14820 ), .Q ( new_AGEMA_signal_14821 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6817 ( .C ( clk ), .D ( new_AGEMA_signal_14844 ), .Q ( new_AGEMA_signal_14845 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6825 ( .C ( clk ), .D ( new_AGEMA_signal_14852 ), .Q ( new_AGEMA_signal_14853 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6833 ( .C ( clk ), .D ( new_AGEMA_signal_14860 ), .Q ( new_AGEMA_signal_14861 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6841 ( .C ( clk ), .D ( new_AGEMA_signal_14868 ), .Q ( new_AGEMA_signal_14869 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6903 ( .C ( clk ), .D ( new_AGEMA_signal_14930 ), .Q ( new_AGEMA_signal_14931 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6919 ( .C ( clk ), .D ( new_AGEMA_signal_14946 ), .Q ( new_AGEMA_signal_14947 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6935 ( .C ( clk ), .D ( new_AGEMA_signal_14962 ), .Q ( new_AGEMA_signal_14963 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6951 ( .C ( clk ), .D ( new_AGEMA_signal_14978 ), .Q ( new_AGEMA_signal_14979 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6961 ( .C ( clk ), .D ( new_AGEMA_signal_14988 ), .Q ( new_AGEMA_signal_14989 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6971 ( .C ( clk ), .D ( new_AGEMA_signal_14998 ), .Q ( new_AGEMA_signal_14999 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6981 ( .C ( clk ), .D ( new_AGEMA_signal_15008 ), .Q ( new_AGEMA_signal_15009 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6991 ( .C ( clk ), .D ( new_AGEMA_signal_15018 ), .Q ( new_AGEMA_signal_15019 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7009 ( .C ( clk ), .D ( new_AGEMA_signal_15036 ), .Q ( new_AGEMA_signal_15037 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7027 ( .C ( clk ), .D ( new_AGEMA_signal_15054 ), .Q ( new_AGEMA_signal_15055 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7045 ( .C ( clk ), .D ( new_AGEMA_signal_15072 ), .Q ( new_AGEMA_signal_15073 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7063 ( .C ( clk ), .D ( new_AGEMA_signal_15090 ), .Q ( new_AGEMA_signal_15091 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7087 ( .C ( clk ), .D ( n2671 ), .Q ( new_AGEMA_signal_15115 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7095 ( .C ( clk ), .D ( new_AGEMA_signal_3489 ), .Q ( new_AGEMA_signal_15123 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7103 ( .C ( clk ), .D ( new_AGEMA_signal_3490 ), .Q ( new_AGEMA_signal_15131 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7111 ( .C ( clk ), .D ( new_AGEMA_signal_3491 ), .Q ( new_AGEMA_signal_15139 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7209 ( .C ( clk ), .D ( new_AGEMA_signal_15236 ), .Q ( new_AGEMA_signal_15237 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7229 ( .C ( clk ), .D ( new_AGEMA_signal_15256 ), .Q ( new_AGEMA_signal_15257 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7249 ( .C ( clk ), .D ( new_AGEMA_signal_15276 ), .Q ( new_AGEMA_signal_15277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7269 ( .C ( clk ), .D ( new_AGEMA_signal_15296 ), .Q ( new_AGEMA_signal_15297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7311 ( .C ( clk ), .D ( n2380 ), .Q ( new_AGEMA_signal_15339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7323 ( .C ( clk ), .D ( new_AGEMA_signal_3474 ), .Q ( new_AGEMA_signal_15351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7335 ( .C ( clk ), .D ( new_AGEMA_signal_3475 ), .Q ( new_AGEMA_signal_15363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7347 ( .C ( clk ), .D ( new_AGEMA_signal_3476 ), .Q ( new_AGEMA_signal_15375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7359 ( .C ( clk ), .D ( n2382 ), .Q ( new_AGEMA_signal_15387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7373 ( .C ( clk ), .D ( new_AGEMA_signal_3471 ), .Q ( new_AGEMA_signal_15401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7387 ( .C ( clk ), .D ( new_AGEMA_signal_3472 ), .Q ( new_AGEMA_signal_15415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7401 ( .C ( clk ), .D ( new_AGEMA_signal_3473 ), .Q ( new_AGEMA_signal_15429 ) ) ;

    /* cells in depth 18 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2016 ( .a ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, n1941}), .b ({new_AGEMA_signal_13418, new_AGEMA_signal_13412, new_AGEMA_signal_13406, new_AGEMA_signal_13400}), .clk ( clk ), .r ({Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758]}), .c ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, new_AGEMA_signal_3507, n2019}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2060 ( .a ({new_AGEMA_signal_13442, new_AGEMA_signal_13436, new_AGEMA_signal_13430, new_AGEMA_signal_13424}), .b ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, n1960}), .clk ( clk ), .r ({Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764]}), .c ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, n2002}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2116 ( .a ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, n1988}), .b ({new_AGEMA_signal_13466, new_AGEMA_signal_13460, new_AGEMA_signal_13454, new_AGEMA_signal_13448}), .clk ( clk ), .r ({Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770]}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, n1989}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2154 ( .a ({new_AGEMA_signal_13482, new_AGEMA_signal_13478, new_AGEMA_signal_13474, new_AGEMA_signal_13470}), .b ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, n2015}), .clk ( clk ), .r ({Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776]}), .c ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, n2016}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2170 ( .a ({new_AGEMA_signal_13514, new_AGEMA_signal_13506, new_AGEMA_signal_13498, new_AGEMA_signal_13490}), .b ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, n2030}), .clk ( clk ), .r ({Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, n2038}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2201 ( .a ({new_AGEMA_signal_13538, new_AGEMA_signal_13532, new_AGEMA_signal_13526, new_AGEMA_signal_13520}), .b ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, n2053}), .clk ( clk ), .r ({Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788]}), .c ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, n2111}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2223 ( .a ({new_AGEMA_signal_13554, new_AGEMA_signal_13550, new_AGEMA_signal_13546, new_AGEMA_signal_13542}), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, new_AGEMA_signal_3441, n2071}), .clk ( clk ), .r ({Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, n2079}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2263 ( .a ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, n2103}), .b ({new_AGEMA_signal_13586, new_AGEMA_signal_13578, new_AGEMA_signal_13570, new_AGEMA_signal_13562}), .clk ( clk ), .r ({Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800]}), .c ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, n2104}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2289 ( .a ({new_AGEMA_signal_13618, new_AGEMA_signal_13610, new_AGEMA_signal_13602, new_AGEMA_signal_13594}), .b ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, new_AGEMA_signal_3447, n2126}), .clk ( clk ), .r ({Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806]}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, n2127}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2315 ( .a ({new_AGEMA_signal_13482, new_AGEMA_signal_13478, new_AGEMA_signal_13474, new_AGEMA_signal_13470}), .b ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, n2146}), .clk ( clk ), .r ({Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812]}), .c ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n2147}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2336 ( .a ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, new_AGEMA_signal_3453, n2173}), .b ({new_AGEMA_signal_13658, new_AGEMA_signal_13648, new_AGEMA_signal_13638, new_AGEMA_signal_13628}), .clk ( clk ), .r ({Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, n2208}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2352 ( .a ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, n2187}), .b ({new_AGEMA_signal_13690, new_AGEMA_signal_13682, new_AGEMA_signal_13674, new_AGEMA_signal_13666}), .clk ( clk ), .r ({Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824]}), .c ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, n2199}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2420 ( .a ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, n2256}), .b ({new_AGEMA_signal_13714, new_AGEMA_signal_13708, new_AGEMA_signal_13702, new_AGEMA_signal_13696}), .clk ( clk ), .r ({Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, n2257}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2442 ( .a ({new_AGEMA_signal_13730, new_AGEMA_signal_13726, new_AGEMA_signal_13722, new_AGEMA_signal_13718}), .b ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, new_AGEMA_signal_3465, n2275}), .clk ( clk ), .r ({Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836]}), .c ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n2281}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2475 ( .a ({new_AGEMA_signal_13754, new_AGEMA_signal_13748, new_AGEMA_signal_13742, new_AGEMA_signal_13736}), .b ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, n2303}), .clk ( clk ), .r ({Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, n2305}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2532 ( .a ({new_AGEMA_signal_13786, new_AGEMA_signal_13778, new_AGEMA_signal_13770, new_AGEMA_signal_13762}), .b ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, new_AGEMA_signal_3477, n2366}), .clk ( clk ), .r ({Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848]}), .c ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, n2368}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2583 ( .a ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, n2425}), .b ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, n2424}), .clk ( clk ), .r ({Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, n2426}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2605 ( .a ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, new_AGEMA_signal_3483, n2451}), .b ({new_AGEMA_signal_13810, new_AGEMA_signal_13804, new_AGEMA_signal_13798, new_AGEMA_signal_13792}), .clk ( clk ), .r ({Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860]}), .c ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2457}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2659 ( .a ({new_AGEMA_signal_13818, new_AGEMA_signal_13816, new_AGEMA_signal_13814, new_AGEMA_signal_13812}), .b ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, n2511}), .clk ( clk ), .r ({Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866]}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, n2513}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2717 ( .a ({new_AGEMA_signal_13850, new_AGEMA_signal_13842, new_AGEMA_signal_13834, new_AGEMA_signal_13826}), .b ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, n2590}), .clk ( clk ), .r ({Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872]}), .c ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, n2592}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2741 ( .a ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, n2623}), .b ({new_AGEMA_signal_13866, new_AGEMA_signal_13862, new_AGEMA_signal_13858, new_AGEMA_signal_13854}), .clk ( clk ), .r ({Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878]}), .c ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, n2637}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2767 ( .a ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, n2667}), .b ({new_AGEMA_signal_13890, new_AGEMA_signal_13884, new_AGEMA_signal_13878, new_AGEMA_signal_13872}), .clk ( clk ), .r ({Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884]}), .c ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, n2668}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2787 ( .a ({new_AGEMA_signal_13914, new_AGEMA_signal_13908, new_AGEMA_signal_13902, new_AGEMA_signal_13896}), .b ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, new_AGEMA_signal_3501, n2703}), .clk ( clk ), .r ({Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890]}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, n2705}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2841 ( .a ({new_AGEMA_signal_13930, new_AGEMA_signal_13926, new_AGEMA_signal_13922, new_AGEMA_signal_13918}), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, n2803}), .clk ( clk ), .r ({Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896]}), .c ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, n2805}) ) ;
    buf_clk new_AGEMA_reg_buffer_5908 ( .C ( clk ), .D ( new_AGEMA_signal_13935 ), .Q ( new_AGEMA_signal_13936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5914 ( .C ( clk ), .D ( new_AGEMA_signal_13941 ), .Q ( new_AGEMA_signal_13942 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5920 ( .C ( clk ), .D ( new_AGEMA_signal_13947 ), .Q ( new_AGEMA_signal_13948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5926 ( .C ( clk ), .D ( new_AGEMA_signal_13953 ), .Q ( new_AGEMA_signal_13954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5930 ( .C ( clk ), .D ( new_AGEMA_signal_13957 ), .Q ( new_AGEMA_signal_13958 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5934 ( .C ( clk ), .D ( new_AGEMA_signal_13961 ), .Q ( new_AGEMA_signal_13962 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5938 ( .C ( clk ), .D ( new_AGEMA_signal_13965 ), .Q ( new_AGEMA_signal_13966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5942 ( .C ( clk ), .D ( new_AGEMA_signal_13969 ), .Q ( new_AGEMA_signal_13970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5948 ( .C ( clk ), .D ( new_AGEMA_signal_13975 ), .Q ( new_AGEMA_signal_13976 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5954 ( .C ( clk ), .D ( new_AGEMA_signal_13981 ), .Q ( new_AGEMA_signal_13982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5960 ( .C ( clk ), .D ( new_AGEMA_signal_13987 ), .Q ( new_AGEMA_signal_13988 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5966 ( .C ( clk ), .D ( new_AGEMA_signal_13993 ), .Q ( new_AGEMA_signal_13994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5976 ( .C ( clk ), .D ( new_AGEMA_signal_14003 ), .Q ( new_AGEMA_signal_14004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5986 ( .C ( clk ), .D ( new_AGEMA_signal_14013 ), .Q ( new_AGEMA_signal_14014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_5996 ( .C ( clk ), .D ( new_AGEMA_signal_14023 ), .Q ( new_AGEMA_signal_14024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6006 ( .C ( clk ), .D ( new_AGEMA_signal_14033 ), .Q ( new_AGEMA_signal_14034 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6012 ( .C ( clk ), .D ( new_AGEMA_signal_14039 ), .Q ( new_AGEMA_signal_14040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6018 ( .C ( clk ), .D ( new_AGEMA_signal_14045 ), .Q ( new_AGEMA_signal_14046 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C ( clk ), .D ( new_AGEMA_signal_14051 ), .Q ( new_AGEMA_signal_14052 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C ( clk ), .D ( new_AGEMA_signal_14057 ), .Q ( new_AGEMA_signal_14058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C ( clk ), .D ( new_AGEMA_signal_14063 ), .Q ( new_AGEMA_signal_14064 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C ( clk ), .D ( new_AGEMA_signal_14069 ), .Q ( new_AGEMA_signal_14070 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C ( clk ), .D ( new_AGEMA_signal_14075 ), .Q ( new_AGEMA_signal_14076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6054 ( .C ( clk ), .D ( new_AGEMA_signal_14081 ), .Q ( new_AGEMA_signal_14082 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6058 ( .C ( clk ), .D ( new_AGEMA_signal_14085 ), .Q ( new_AGEMA_signal_14086 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6062 ( .C ( clk ), .D ( new_AGEMA_signal_14089 ), .Q ( new_AGEMA_signal_14090 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6066 ( .C ( clk ), .D ( new_AGEMA_signal_14093 ), .Q ( new_AGEMA_signal_14094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6070 ( .C ( clk ), .D ( new_AGEMA_signal_14097 ), .Q ( new_AGEMA_signal_14098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6074 ( .C ( clk ), .D ( new_AGEMA_signal_14101 ), .Q ( new_AGEMA_signal_14102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6078 ( .C ( clk ), .D ( new_AGEMA_signal_14105 ), .Q ( new_AGEMA_signal_14106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6082 ( .C ( clk ), .D ( new_AGEMA_signal_14109 ), .Q ( new_AGEMA_signal_14110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6086 ( .C ( clk ), .D ( new_AGEMA_signal_14113 ), .Q ( new_AGEMA_signal_14114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6094 ( .C ( clk ), .D ( new_AGEMA_signal_14121 ), .Q ( new_AGEMA_signal_14122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6102 ( .C ( clk ), .D ( new_AGEMA_signal_14129 ), .Q ( new_AGEMA_signal_14130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6110 ( .C ( clk ), .D ( new_AGEMA_signal_14137 ), .Q ( new_AGEMA_signal_14138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6118 ( .C ( clk ), .D ( new_AGEMA_signal_14145 ), .Q ( new_AGEMA_signal_14146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6124 ( .C ( clk ), .D ( new_AGEMA_signal_14151 ), .Q ( new_AGEMA_signal_14152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6130 ( .C ( clk ), .D ( new_AGEMA_signal_14157 ), .Q ( new_AGEMA_signal_14158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6136 ( .C ( clk ), .D ( new_AGEMA_signal_14163 ), .Q ( new_AGEMA_signal_14164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6142 ( .C ( clk ), .D ( new_AGEMA_signal_14169 ), .Q ( new_AGEMA_signal_14170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6150 ( .C ( clk ), .D ( new_AGEMA_signal_14177 ), .Q ( new_AGEMA_signal_14178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6158 ( .C ( clk ), .D ( new_AGEMA_signal_14185 ), .Q ( new_AGEMA_signal_14186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6166 ( .C ( clk ), .D ( new_AGEMA_signal_14193 ), .Q ( new_AGEMA_signal_14194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6174 ( .C ( clk ), .D ( new_AGEMA_signal_14201 ), .Q ( new_AGEMA_signal_14202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6182 ( .C ( clk ), .D ( new_AGEMA_signal_14209 ), .Q ( new_AGEMA_signal_14210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6190 ( .C ( clk ), .D ( new_AGEMA_signal_14217 ), .Q ( new_AGEMA_signal_14218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6198 ( .C ( clk ), .D ( new_AGEMA_signal_14225 ), .Q ( new_AGEMA_signal_14226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6206 ( .C ( clk ), .D ( new_AGEMA_signal_14233 ), .Q ( new_AGEMA_signal_14234 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6208 ( .C ( clk ), .D ( new_AGEMA_signal_14235 ), .Q ( new_AGEMA_signal_14236 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6210 ( .C ( clk ), .D ( new_AGEMA_signal_14237 ), .Q ( new_AGEMA_signal_14238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6212 ( .C ( clk ), .D ( new_AGEMA_signal_14239 ), .Q ( new_AGEMA_signal_14240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6214 ( .C ( clk ), .D ( new_AGEMA_signal_14241 ), .Q ( new_AGEMA_signal_14242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6218 ( .C ( clk ), .D ( new_AGEMA_signal_14245 ), .Q ( new_AGEMA_signal_14246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6222 ( .C ( clk ), .D ( new_AGEMA_signal_14249 ), .Q ( new_AGEMA_signal_14250 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6226 ( .C ( clk ), .D ( new_AGEMA_signal_14253 ), .Q ( new_AGEMA_signal_14254 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6230 ( .C ( clk ), .D ( new_AGEMA_signal_14257 ), .Q ( new_AGEMA_signal_14258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6234 ( .C ( clk ), .D ( new_AGEMA_signal_14261 ), .Q ( new_AGEMA_signal_14262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6238 ( .C ( clk ), .D ( new_AGEMA_signal_14265 ), .Q ( new_AGEMA_signal_14266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6242 ( .C ( clk ), .D ( new_AGEMA_signal_14269 ), .Q ( new_AGEMA_signal_14270 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6246 ( .C ( clk ), .D ( new_AGEMA_signal_14273 ), .Q ( new_AGEMA_signal_14274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6254 ( .C ( clk ), .D ( new_AGEMA_signal_14281 ), .Q ( new_AGEMA_signal_14282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6262 ( .C ( clk ), .D ( new_AGEMA_signal_14289 ), .Q ( new_AGEMA_signal_14290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6270 ( .C ( clk ), .D ( new_AGEMA_signal_14297 ), .Q ( new_AGEMA_signal_14298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6278 ( .C ( clk ), .D ( new_AGEMA_signal_14305 ), .Q ( new_AGEMA_signal_14306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6282 ( .C ( clk ), .D ( new_AGEMA_signal_14309 ), .Q ( new_AGEMA_signal_14310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6286 ( .C ( clk ), .D ( new_AGEMA_signal_14313 ), .Q ( new_AGEMA_signal_14314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6290 ( .C ( clk ), .D ( new_AGEMA_signal_14317 ), .Q ( new_AGEMA_signal_14318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6294 ( .C ( clk ), .D ( new_AGEMA_signal_14321 ), .Q ( new_AGEMA_signal_14322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6300 ( .C ( clk ), .D ( new_AGEMA_signal_14327 ), .Q ( new_AGEMA_signal_14328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6308 ( .C ( clk ), .D ( new_AGEMA_signal_14335 ), .Q ( new_AGEMA_signal_14336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6316 ( .C ( clk ), .D ( new_AGEMA_signal_14343 ), .Q ( new_AGEMA_signal_14344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6324 ( .C ( clk ), .D ( new_AGEMA_signal_14351 ), .Q ( new_AGEMA_signal_14352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6336 ( .C ( clk ), .D ( new_AGEMA_signal_14363 ), .Q ( new_AGEMA_signal_14364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6348 ( .C ( clk ), .D ( new_AGEMA_signal_14375 ), .Q ( new_AGEMA_signal_14376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6360 ( .C ( clk ), .D ( new_AGEMA_signal_14387 ), .Q ( new_AGEMA_signal_14388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6372 ( .C ( clk ), .D ( new_AGEMA_signal_14399 ), .Q ( new_AGEMA_signal_14400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6386 ( .C ( clk ), .D ( new_AGEMA_signal_14413 ), .Q ( new_AGEMA_signal_14414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6400 ( .C ( clk ), .D ( new_AGEMA_signal_14427 ), .Q ( new_AGEMA_signal_14428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6414 ( .C ( clk ), .D ( new_AGEMA_signal_14441 ), .Q ( new_AGEMA_signal_14442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6428 ( .C ( clk ), .D ( new_AGEMA_signal_14455 ), .Q ( new_AGEMA_signal_14456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6436 ( .C ( clk ), .D ( new_AGEMA_signal_14463 ), .Q ( new_AGEMA_signal_14464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6444 ( .C ( clk ), .D ( new_AGEMA_signal_14471 ), .Q ( new_AGEMA_signal_14472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6452 ( .C ( clk ), .D ( new_AGEMA_signal_14479 ), .Q ( new_AGEMA_signal_14480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6460 ( .C ( clk ), .D ( new_AGEMA_signal_14487 ), .Q ( new_AGEMA_signal_14488 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6474 ( .C ( clk ), .D ( new_AGEMA_signal_14501 ), .Q ( new_AGEMA_signal_14502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6488 ( .C ( clk ), .D ( new_AGEMA_signal_14515 ), .Q ( new_AGEMA_signal_14516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6502 ( .C ( clk ), .D ( new_AGEMA_signal_14529 ), .Q ( new_AGEMA_signal_14530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6516 ( .C ( clk ), .D ( new_AGEMA_signal_14543 ), .Q ( new_AGEMA_signal_14544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6524 ( .C ( clk ), .D ( new_AGEMA_signal_14551 ), .Q ( new_AGEMA_signal_14552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6532 ( .C ( clk ), .D ( new_AGEMA_signal_14559 ), .Q ( new_AGEMA_signal_14560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6540 ( .C ( clk ), .D ( new_AGEMA_signal_14567 ), .Q ( new_AGEMA_signal_14568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6548 ( .C ( clk ), .D ( new_AGEMA_signal_14575 ), .Q ( new_AGEMA_signal_14576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6556 ( .C ( clk ), .D ( new_AGEMA_signal_14583 ), .Q ( new_AGEMA_signal_14584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6564 ( .C ( clk ), .D ( new_AGEMA_signal_14591 ), .Q ( new_AGEMA_signal_14592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6572 ( .C ( clk ), .D ( new_AGEMA_signal_14599 ), .Q ( new_AGEMA_signal_14600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6580 ( .C ( clk ), .D ( new_AGEMA_signal_14607 ), .Q ( new_AGEMA_signal_14608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6618 ( .C ( clk ), .D ( new_AGEMA_signal_14645 ), .Q ( new_AGEMA_signal_14646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6634 ( .C ( clk ), .D ( new_AGEMA_signal_14661 ), .Q ( new_AGEMA_signal_14662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6650 ( .C ( clk ), .D ( new_AGEMA_signal_14677 ), .Q ( new_AGEMA_signal_14678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6666 ( .C ( clk ), .D ( new_AGEMA_signal_14693 ), .Q ( new_AGEMA_signal_14694 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6706 ( .C ( clk ), .D ( new_AGEMA_signal_14733 ), .Q ( new_AGEMA_signal_14734 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6722 ( .C ( clk ), .D ( new_AGEMA_signal_14749 ), .Q ( new_AGEMA_signal_14750 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6738 ( .C ( clk ), .D ( new_AGEMA_signal_14765 ), .Q ( new_AGEMA_signal_14766 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6754 ( .C ( clk ), .D ( new_AGEMA_signal_14781 ), .Q ( new_AGEMA_signal_14782 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6764 ( .C ( clk ), .D ( new_AGEMA_signal_14791 ), .Q ( new_AGEMA_signal_14792 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6774 ( .C ( clk ), .D ( new_AGEMA_signal_14801 ), .Q ( new_AGEMA_signal_14802 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6784 ( .C ( clk ), .D ( new_AGEMA_signal_14811 ), .Q ( new_AGEMA_signal_14812 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6794 ( .C ( clk ), .D ( new_AGEMA_signal_14821 ), .Q ( new_AGEMA_signal_14822 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6818 ( .C ( clk ), .D ( new_AGEMA_signal_14845 ), .Q ( new_AGEMA_signal_14846 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6826 ( .C ( clk ), .D ( new_AGEMA_signal_14853 ), .Q ( new_AGEMA_signal_14854 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6834 ( .C ( clk ), .D ( new_AGEMA_signal_14861 ), .Q ( new_AGEMA_signal_14862 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6842 ( .C ( clk ), .D ( new_AGEMA_signal_14869 ), .Q ( new_AGEMA_signal_14870 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6904 ( .C ( clk ), .D ( new_AGEMA_signal_14931 ), .Q ( new_AGEMA_signal_14932 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6920 ( .C ( clk ), .D ( new_AGEMA_signal_14947 ), .Q ( new_AGEMA_signal_14948 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6936 ( .C ( clk ), .D ( new_AGEMA_signal_14963 ), .Q ( new_AGEMA_signal_14964 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6952 ( .C ( clk ), .D ( new_AGEMA_signal_14979 ), .Q ( new_AGEMA_signal_14980 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6962 ( .C ( clk ), .D ( new_AGEMA_signal_14989 ), .Q ( new_AGEMA_signal_14990 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6972 ( .C ( clk ), .D ( new_AGEMA_signal_14999 ), .Q ( new_AGEMA_signal_15000 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6982 ( .C ( clk ), .D ( new_AGEMA_signal_15009 ), .Q ( new_AGEMA_signal_15010 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6992 ( .C ( clk ), .D ( new_AGEMA_signal_15019 ), .Q ( new_AGEMA_signal_15020 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7010 ( .C ( clk ), .D ( new_AGEMA_signal_15037 ), .Q ( new_AGEMA_signal_15038 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7028 ( .C ( clk ), .D ( new_AGEMA_signal_15055 ), .Q ( new_AGEMA_signal_15056 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7046 ( .C ( clk ), .D ( new_AGEMA_signal_15073 ), .Q ( new_AGEMA_signal_15074 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7064 ( .C ( clk ), .D ( new_AGEMA_signal_15091 ), .Q ( new_AGEMA_signal_15092 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7088 ( .C ( clk ), .D ( new_AGEMA_signal_15115 ), .Q ( new_AGEMA_signal_15116 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7096 ( .C ( clk ), .D ( new_AGEMA_signal_15123 ), .Q ( new_AGEMA_signal_15124 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7104 ( .C ( clk ), .D ( new_AGEMA_signal_15131 ), .Q ( new_AGEMA_signal_15132 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7112 ( .C ( clk ), .D ( new_AGEMA_signal_15139 ), .Q ( new_AGEMA_signal_15140 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7210 ( .C ( clk ), .D ( new_AGEMA_signal_15237 ), .Q ( new_AGEMA_signal_15238 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7230 ( .C ( clk ), .D ( new_AGEMA_signal_15257 ), .Q ( new_AGEMA_signal_15258 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7250 ( .C ( clk ), .D ( new_AGEMA_signal_15277 ), .Q ( new_AGEMA_signal_15278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7270 ( .C ( clk ), .D ( new_AGEMA_signal_15297 ), .Q ( new_AGEMA_signal_15298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7312 ( .C ( clk ), .D ( new_AGEMA_signal_15339 ), .Q ( new_AGEMA_signal_15340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7324 ( .C ( clk ), .D ( new_AGEMA_signal_15351 ), .Q ( new_AGEMA_signal_15352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7336 ( .C ( clk ), .D ( new_AGEMA_signal_15363 ), .Q ( new_AGEMA_signal_15364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7348 ( .C ( clk ), .D ( new_AGEMA_signal_15375 ), .Q ( new_AGEMA_signal_15376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7360 ( .C ( clk ), .D ( new_AGEMA_signal_15387 ), .Q ( new_AGEMA_signal_15388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7374 ( .C ( clk ), .D ( new_AGEMA_signal_15401 ), .Q ( new_AGEMA_signal_15402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7388 ( .C ( clk ), .D ( new_AGEMA_signal_15415 ), .Q ( new_AGEMA_signal_15416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7402 ( .C ( clk ), .D ( new_AGEMA_signal_15429 ), .Q ( new_AGEMA_signal_15430 ) ) ;

    /* cells in depth 19 */
    buf_clk new_AGEMA_reg_buffer_6301 ( .C ( clk ), .D ( new_AGEMA_signal_14328 ), .Q ( new_AGEMA_signal_14329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6309 ( .C ( clk ), .D ( new_AGEMA_signal_14336 ), .Q ( new_AGEMA_signal_14337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6317 ( .C ( clk ), .D ( new_AGEMA_signal_14344 ), .Q ( new_AGEMA_signal_14345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6325 ( .C ( clk ), .D ( new_AGEMA_signal_14352 ), .Q ( new_AGEMA_signal_14353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6337 ( .C ( clk ), .D ( new_AGEMA_signal_14364 ), .Q ( new_AGEMA_signal_14365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6349 ( .C ( clk ), .D ( new_AGEMA_signal_14376 ), .Q ( new_AGEMA_signal_14377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6361 ( .C ( clk ), .D ( new_AGEMA_signal_14388 ), .Q ( new_AGEMA_signal_14389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6373 ( .C ( clk ), .D ( new_AGEMA_signal_14400 ), .Q ( new_AGEMA_signal_14401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6387 ( .C ( clk ), .D ( new_AGEMA_signal_14414 ), .Q ( new_AGEMA_signal_14415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6401 ( .C ( clk ), .D ( new_AGEMA_signal_14428 ), .Q ( new_AGEMA_signal_14429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6415 ( .C ( clk ), .D ( new_AGEMA_signal_14442 ), .Q ( new_AGEMA_signal_14443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6429 ( .C ( clk ), .D ( new_AGEMA_signal_14456 ), .Q ( new_AGEMA_signal_14457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6437 ( .C ( clk ), .D ( new_AGEMA_signal_14464 ), .Q ( new_AGEMA_signal_14465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6445 ( .C ( clk ), .D ( new_AGEMA_signal_14472 ), .Q ( new_AGEMA_signal_14473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6453 ( .C ( clk ), .D ( new_AGEMA_signal_14480 ), .Q ( new_AGEMA_signal_14481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6461 ( .C ( clk ), .D ( new_AGEMA_signal_14488 ), .Q ( new_AGEMA_signal_14489 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6475 ( .C ( clk ), .D ( new_AGEMA_signal_14502 ), .Q ( new_AGEMA_signal_14503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6489 ( .C ( clk ), .D ( new_AGEMA_signal_14516 ), .Q ( new_AGEMA_signal_14517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6503 ( .C ( clk ), .D ( new_AGEMA_signal_14530 ), .Q ( new_AGEMA_signal_14531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6517 ( .C ( clk ), .D ( new_AGEMA_signal_14544 ), .Q ( new_AGEMA_signal_14545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6525 ( .C ( clk ), .D ( new_AGEMA_signal_14552 ), .Q ( new_AGEMA_signal_14553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6533 ( .C ( clk ), .D ( new_AGEMA_signal_14560 ), .Q ( new_AGEMA_signal_14561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6541 ( .C ( clk ), .D ( new_AGEMA_signal_14568 ), .Q ( new_AGEMA_signal_14569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6549 ( .C ( clk ), .D ( new_AGEMA_signal_14576 ), .Q ( new_AGEMA_signal_14577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6557 ( .C ( clk ), .D ( new_AGEMA_signal_14584 ), .Q ( new_AGEMA_signal_14585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6565 ( .C ( clk ), .D ( new_AGEMA_signal_14592 ), .Q ( new_AGEMA_signal_14593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6573 ( .C ( clk ), .D ( new_AGEMA_signal_14600 ), .Q ( new_AGEMA_signal_14601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6581 ( .C ( clk ), .D ( new_AGEMA_signal_14608 ), .Q ( new_AGEMA_signal_14609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6583 ( .C ( clk ), .D ( n2002 ), .Q ( new_AGEMA_signal_14611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6587 ( .C ( clk ), .D ( new_AGEMA_signal_3510 ), .Q ( new_AGEMA_signal_14615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6591 ( .C ( clk ), .D ( new_AGEMA_signal_3511 ), .Q ( new_AGEMA_signal_14619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6595 ( .C ( clk ), .D ( new_AGEMA_signal_3512 ), .Q ( new_AGEMA_signal_14623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6619 ( .C ( clk ), .D ( new_AGEMA_signal_14646 ), .Q ( new_AGEMA_signal_14647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6635 ( .C ( clk ), .D ( new_AGEMA_signal_14662 ), .Q ( new_AGEMA_signal_14663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6651 ( .C ( clk ), .D ( new_AGEMA_signal_14678 ), .Q ( new_AGEMA_signal_14679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6667 ( .C ( clk ), .D ( new_AGEMA_signal_14694 ), .Q ( new_AGEMA_signal_14695 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6671 ( .C ( clk ), .D ( n2208 ), .Q ( new_AGEMA_signal_14699 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6675 ( .C ( clk ), .D ( new_AGEMA_signal_3537 ), .Q ( new_AGEMA_signal_14703 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6679 ( .C ( clk ), .D ( new_AGEMA_signal_3538 ), .Q ( new_AGEMA_signal_14707 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6683 ( .C ( clk ), .D ( new_AGEMA_signal_3539 ), .Q ( new_AGEMA_signal_14711 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6707 ( .C ( clk ), .D ( new_AGEMA_signal_14734 ), .Q ( new_AGEMA_signal_14735 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6723 ( .C ( clk ), .D ( new_AGEMA_signal_14750 ), .Q ( new_AGEMA_signal_14751 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6739 ( .C ( clk ), .D ( new_AGEMA_signal_14766 ), .Q ( new_AGEMA_signal_14767 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6755 ( .C ( clk ), .D ( new_AGEMA_signal_14782 ), .Q ( new_AGEMA_signal_14783 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6765 ( .C ( clk ), .D ( new_AGEMA_signal_14792 ), .Q ( new_AGEMA_signal_14793 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6775 ( .C ( clk ), .D ( new_AGEMA_signal_14802 ), .Q ( new_AGEMA_signal_14803 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6785 ( .C ( clk ), .D ( new_AGEMA_signal_14812 ), .Q ( new_AGEMA_signal_14813 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6795 ( .C ( clk ), .D ( new_AGEMA_signal_14822 ), .Q ( new_AGEMA_signal_14823 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6799 ( .C ( clk ), .D ( n2668 ), .Q ( new_AGEMA_signal_14827 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6803 ( .C ( clk ), .D ( new_AGEMA_signal_3570 ), .Q ( new_AGEMA_signal_14831 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6807 ( .C ( clk ), .D ( new_AGEMA_signal_3571 ), .Q ( new_AGEMA_signal_14835 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6811 ( .C ( clk ), .D ( new_AGEMA_signal_3572 ), .Q ( new_AGEMA_signal_14839 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6819 ( .C ( clk ), .D ( new_AGEMA_signal_14846 ), .Q ( new_AGEMA_signal_14847 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6827 ( .C ( clk ), .D ( new_AGEMA_signal_14854 ), .Q ( new_AGEMA_signal_14855 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6835 ( .C ( clk ), .D ( new_AGEMA_signal_14862 ), .Q ( new_AGEMA_signal_14863 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6843 ( .C ( clk ), .D ( new_AGEMA_signal_14870 ), .Q ( new_AGEMA_signal_14871 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6847 ( .C ( clk ), .D ( n2016 ), .Q ( new_AGEMA_signal_14875 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6853 ( .C ( clk ), .D ( new_AGEMA_signal_3516 ), .Q ( new_AGEMA_signal_14881 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6859 ( .C ( clk ), .D ( new_AGEMA_signal_3517 ), .Q ( new_AGEMA_signal_14887 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6865 ( .C ( clk ), .D ( new_AGEMA_signal_3518 ), .Q ( new_AGEMA_signal_14893 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6871 ( .C ( clk ), .D ( n2111 ), .Q ( new_AGEMA_signal_14899 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6877 ( .C ( clk ), .D ( new_AGEMA_signal_3522 ), .Q ( new_AGEMA_signal_14905 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6883 ( .C ( clk ), .D ( new_AGEMA_signal_3523 ), .Q ( new_AGEMA_signal_14911 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6889 ( .C ( clk ), .D ( new_AGEMA_signal_3524 ), .Q ( new_AGEMA_signal_14917 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6905 ( .C ( clk ), .D ( new_AGEMA_signal_14932 ), .Q ( new_AGEMA_signal_14933 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6921 ( .C ( clk ), .D ( new_AGEMA_signal_14948 ), .Q ( new_AGEMA_signal_14949 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6937 ( .C ( clk ), .D ( new_AGEMA_signal_14964 ), .Q ( new_AGEMA_signal_14965 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6953 ( .C ( clk ), .D ( new_AGEMA_signal_14980 ), .Q ( new_AGEMA_signal_14981 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6963 ( .C ( clk ), .D ( new_AGEMA_signal_14990 ), .Q ( new_AGEMA_signal_14991 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6973 ( .C ( clk ), .D ( new_AGEMA_signal_15000 ), .Q ( new_AGEMA_signal_15001 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6983 ( .C ( clk ), .D ( new_AGEMA_signal_15010 ), .Q ( new_AGEMA_signal_15011 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6993 ( .C ( clk ), .D ( new_AGEMA_signal_15020 ), .Q ( new_AGEMA_signal_15021 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7011 ( .C ( clk ), .D ( new_AGEMA_signal_15038 ), .Q ( new_AGEMA_signal_15039 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7029 ( .C ( clk ), .D ( new_AGEMA_signal_15056 ), .Q ( new_AGEMA_signal_15057 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7047 ( .C ( clk ), .D ( new_AGEMA_signal_15074 ), .Q ( new_AGEMA_signal_15075 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7065 ( .C ( clk ), .D ( new_AGEMA_signal_15092 ), .Q ( new_AGEMA_signal_15093 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7089 ( .C ( clk ), .D ( new_AGEMA_signal_15116 ), .Q ( new_AGEMA_signal_15117 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7097 ( .C ( clk ), .D ( new_AGEMA_signal_15124 ), .Q ( new_AGEMA_signal_15125 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7105 ( .C ( clk ), .D ( new_AGEMA_signal_15132 ), .Q ( new_AGEMA_signal_15133 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7113 ( .C ( clk ), .D ( new_AGEMA_signal_15140 ), .Q ( new_AGEMA_signal_15141 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7135 ( .C ( clk ), .D ( n2019 ), .Q ( new_AGEMA_signal_15163 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7143 ( .C ( clk ), .D ( new_AGEMA_signal_3507 ), .Q ( new_AGEMA_signal_15171 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7151 ( .C ( clk ), .D ( new_AGEMA_signal_3508 ), .Q ( new_AGEMA_signal_15179 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7159 ( .C ( clk ), .D ( new_AGEMA_signal_3509 ), .Q ( new_AGEMA_signal_15187 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7211 ( .C ( clk ), .D ( new_AGEMA_signal_15238 ), .Q ( new_AGEMA_signal_15239 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7231 ( .C ( clk ), .D ( new_AGEMA_signal_15258 ), .Q ( new_AGEMA_signal_15259 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7251 ( .C ( clk ), .D ( new_AGEMA_signal_15278 ), .Q ( new_AGEMA_signal_15279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7271 ( .C ( clk ), .D ( new_AGEMA_signal_15298 ), .Q ( new_AGEMA_signal_15299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7313 ( .C ( clk ), .D ( new_AGEMA_signal_15340 ), .Q ( new_AGEMA_signal_15341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7325 ( .C ( clk ), .D ( new_AGEMA_signal_15352 ), .Q ( new_AGEMA_signal_15353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7337 ( .C ( clk ), .D ( new_AGEMA_signal_15364 ), .Q ( new_AGEMA_signal_15365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7349 ( .C ( clk ), .D ( new_AGEMA_signal_15376 ), .Q ( new_AGEMA_signal_15377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7361 ( .C ( clk ), .D ( new_AGEMA_signal_15388 ), .Q ( new_AGEMA_signal_15389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7375 ( .C ( clk ), .D ( new_AGEMA_signal_15402 ), .Q ( new_AGEMA_signal_15403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7389 ( .C ( clk ), .D ( new_AGEMA_signal_15416 ), .Q ( new_AGEMA_signal_15417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7403 ( .C ( clk ), .D ( new_AGEMA_signal_15430 ), .Q ( new_AGEMA_signal_15431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7415 ( .C ( clk ), .D ( n2426 ), .Q ( new_AGEMA_signal_15443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7429 ( .C ( clk ), .D ( new_AGEMA_signal_3555 ), .Q ( new_AGEMA_signal_15457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7443 ( .C ( clk ), .D ( new_AGEMA_signal_3556 ), .Q ( new_AGEMA_signal_15471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7457 ( .C ( clk ), .D ( new_AGEMA_signal_3557 ), .Q ( new_AGEMA_signal_15485 ) ) ;

    /* cells in depth 20 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2117 ( .a ({new_AGEMA_signal_13954, new_AGEMA_signal_13948, new_AGEMA_signal_13942, new_AGEMA_signal_13936}), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, n1989}), .clk ( clk ), .r ({Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, n2000}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2181 ( .a ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, new_AGEMA_signal_3435, n2038}), .b ({new_AGEMA_signal_13970, new_AGEMA_signal_13966, new_AGEMA_signal_13962, new_AGEMA_signal_13958}), .clk ( clk ), .r ({Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, n2113}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2231 ( .a ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, n2079}), .b ({new_AGEMA_signal_13994, new_AGEMA_signal_13988, new_AGEMA_signal_13982, new_AGEMA_signal_13976}), .clk ( clk ), .r ({Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914]}), .c ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, n2109}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2264 ( .a ({new_AGEMA_signal_14034, new_AGEMA_signal_14024, new_AGEMA_signal_14014, new_AGEMA_signal_14004}), .b ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, n2104}), .clk ( clk ), .r ({Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, n2107}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2290 ( .a ({new_AGEMA_signal_14058, new_AGEMA_signal_14052, new_AGEMA_signal_14046, new_AGEMA_signal_14040}), .b ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, n2127}), .clk ( clk ), .r ({Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926]}), .c ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, n2212}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2316 ( .a ({new_AGEMA_signal_14082, new_AGEMA_signal_14076, new_AGEMA_signal_14070, new_AGEMA_signal_14064}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, n2147}), .clk ( clk ), .r ({Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, n2149}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2366 ( .a ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, n2199}), .b ({new_AGEMA_signal_14098, new_AGEMA_signal_14094, new_AGEMA_signal_14090, new_AGEMA_signal_14086}), .clk ( clk ), .r ({Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938]}), .c ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2206}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2421 ( .a ({new_AGEMA_signal_14114, new_AGEMA_signal_14110, new_AGEMA_signal_14106, new_AGEMA_signal_14102}), .b ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, n2257}), .clk ( clk ), .r ({Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, n2310}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2447 ( .a ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, n2281}), .b ({new_AGEMA_signal_14146, new_AGEMA_signal_14138, new_AGEMA_signal_14130, new_AGEMA_signal_14122}), .clk ( clk ), .r ({Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950]}), .c ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, n2308}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2476 ( .a ({new_AGEMA_signal_14170, new_AGEMA_signal_14164, new_AGEMA_signal_14158, new_AGEMA_signal_14152}), .b ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, n2305}), .clk ( clk ), .r ({Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, n2307}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2533 ( .a ({new_AGEMA_signal_14202, new_AGEMA_signal_14194, new_AGEMA_signal_14186, new_AGEMA_signal_14178}), .b ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, n2368}), .clk ( clk ), .r ({Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962]}), .c ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2370}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2611 ( .a ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, n2457}), .b ({new_AGEMA_signal_14234, new_AGEMA_signal_14226, new_AGEMA_signal_14218, new_AGEMA_signal_14210}), .clk ( clk ), .r ({Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, n2530}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2660 ( .a ({new_AGEMA_signal_14242, new_AGEMA_signal_14240, new_AGEMA_signal_14238, new_AGEMA_signal_14236}), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, n2513}), .clk ( clk ), .r ({Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974]}), .c ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, n2515}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2718 ( .a ({new_AGEMA_signal_14258, new_AGEMA_signal_14254, new_AGEMA_signal_14250, new_AGEMA_signal_14246}), .b ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, n2592}), .clk ( clk ), .r ({Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, n2639}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2749 ( .a ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, new_AGEMA_signal_3495, n2637}), .b ({new_AGEMA_signal_14274, new_AGEMA_signal_14270, new_AGEMA_signal_14266, new_AGEMA_signal_14262}), .clk ( clk ), .r ({Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986]}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, n2638}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2788 ( .a ({new_AGEMA_signal_14306, new_AGEMA_signal_14298, new_AGEMA_signal_14290, new_AGEMA_signal_14282}), .b ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, n2705}), .clk ( clk ), .r ({Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992]}), .c ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, n2832}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2842 ( .a ({new_AGEMA_signal_14322, new_AGEMA_signal_14318, new_AGEMA_signal_14314, new_AGEMA_signal_14310}), .b ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, n2805}), .clk ( clk ), .r ({Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998]}), .c ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, n2807}) ) ;
    buf_clk new_AGEMA_reg_buffer_6302 ( .C ( clk ), .D ( new_AGEMA_signal_14329 ), .Q ( new_AGEMA_signal_14330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6310 ( .C ( clk ), .D ( new_AGEMA_signal_14337 ), .Q ( new_AGEMA_signal_14338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6318 ( .C ( clk ), .D ( new_AGEMA_signal_14345 ), .Q ( new_AGEMA_signal_14346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6326 ( .C ( clk ), .D ( new_AGEMA_signal_14353 ), .Q ( new_AGEMA_signal_14354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6338 ( .C ( clk ), .D ( new_AGEMA_signal_14365 ), .Q ( new_AGEMA_signal_14366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6350 ( .C ( clk ), .D ( new_AGEMA_signal_14377 ), .Q ( new_AGEMA_signal_14378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6362 ( .C ( clk ), .D ( new_AGEMA_signal_14389 ), .Q ( new_AGEMA_signal_14390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6374 ( .C ( clk ), .D ( new_AGEMA_signal_14401 ), .Q ( new_AGEMA_signal_14402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6388 ( .C ( clk ), .D ( new_AGEMA_signal_14415 ), .Q ( new_AGEMA_signal_14416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6402 ( .C ( clk ), .D ( new_AGEMA_signal_14429 ), .Q ( new_AGEMA_signal_14430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6416 ( .C ( clk ), .D ( new_AGEMA_signal_14443 ), .Q ( new_AGEMA_signal_14444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6430 ( .C ( clk ), .D ( new_AGEMA_signal_14457 ), .Q ( new_AGEMA_signal_14458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6438 ( .C ( clk ), .D ( new_AGEMA_signal_14465 ), .Q ( new_AGEMA_signal_14466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6446 ( .C ( clk ), .D ( new_AGEMA_signal_14473 ), .Q ( new_AGEMA_signal_14474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6454 ( .C ( clk ), .D ( new_AGEMA_signal_14481 ), .Q ( new_AGEMA_signal_14482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6462 ( .C ( clk ), .D ( new_AGEMA_signal_14489 ), .Q ( new_AGEMA_signal_14490 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6476 ( .C ( clk ), .D ( new_AGEMA_signal_14503 ), .Q ( new_AGEMA_signal_14504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6490 ( .C ( clk ), .D ( new_AGEMA_signal_14517 ), .Q ( new_AGEMA_signal_14518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6504 ( .C ( clk ), .D ( new_AGEMA_signal_14531 ), .Q ( new_AGEMA_signal_14532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6518 ( .C ( clk ), .D ( new_AGEMA_signal_14545 ), .Q ( new_AGEMA_signal_14546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6526 ( .C ( clk ), .D ( new_AGEMA_signal_14553 ), .Q ( new_AGEMA_signal_14554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6534 ( .C ( clk ), .D ( new_AGEMA_signal_14561 ), .Q ( new_AGEMA_signal_14562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6542 ( .C ( clk ), .D ( new_AGEMA_signal_14569 ), .Q ( new_AGEMA_signal_14570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6550 ( .C ( clk ), .D ( new_AGEMA_signal_14577 ), .Q ( new_AGEMA_signal_14578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6558 ( .C ( clk ), .D ( new_AGEMA_signal_14585 ), .Q ( new_AGEMA_signal_14586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6566 ( .C ( clk ), .D ( new_AGEMA_signal_14593 ), .Q ( new_AGEMA_signal_14594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6574 ( .C ( clk ), .D ( new_AGEMA_signal_14601 ), .Q ( new_AGEMA_signal_14602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6582 ( .C ( clk ), .D ( new_AGEMA_signal_14609 ), .Q ( new_AGEMA_signal_14610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6584 ( .C ( clk ), .D ( new_AGEMA_signal_14611 ), .Q ( new_AGEMA_signal_14612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6588 ( .C ( clk ), .D ( new_AGEMA_signal_14615 ), .Q ( new_AGEMA_signal_14616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6592 ( .C ( clk ), .D ( new_AGEMA_signal_14619 ), .Q ( new_AGEMA_signal_14620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6596 ( .C ( clk ), .D ( new_AGEMA_signal_14623 ), .Q ( new_AGEMA_signal_14624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6620 ( .C ( clk ), .D ( new_AGEMA_signal_14647 ), .Q ( new_AGEMA_signal_14648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6636 ( .C ( clk ), .D ( new_AGEMA_signal_14663 ), .Q ( new_AGEMA_signal_14664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6652 ( .C ( clk ), .D ( new_AGEMA_signal_14679 ), .Q ( new_AGEMA_signal_14680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6668 ( .C ( clk ), .D ( new_AGEMA_signal_14695 ), .Q ( new_AGEMA_signal_14696 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6672 ( .C ( clk ), .D ( new_AGEMA_signal_14699 ), .Q ( new_AGEMA_signal_14700 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6676 ( .C ( clk ), .D ( new_AGEMA_signal_14703 ), .Q ( new_AGEMA_signal_14704 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6680 ( .C ( clk ), .D ( new_AGEMA_signal_14707 ), .Q ( new_AGEMA_signal_14708 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6684 ( .C ( clk ), .D ( new_AGEMA_signal_14711 ), .Q ( new_AGEMA_signal_14712 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6708 ( .C ( clk ), .D ( new_AGEMA_signal_14735 ), .Q ( new_AGEMA_signal_14736 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6724 ( .C ( clk ), .D ( new_AGEMA_signal_14751 ), .Q ( new_AGEMA_signal_14752 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6740 ( .C ( clk ), .D ( new_AGEMA_signal_14767 ), .Q ( new_AGEMA_signal_14768 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6756 ( .C ( clk ), .D ( new_AGEMA_signal_14783 ), .Q ( new_AGEMA_signal_14784 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6766 ( .C ( clk ), .D ( new_AGEMA_signal_14793 ), .Q ( new_AGEMA_signal_14794 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6776 ( .C ( clk ), .D ( new_AGEMA_signal_14803 ), .Q ( new_AGEMA_signal_14804 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6786 ( .C ( clk ), .D ( new_AGEMA_signal_14813 ), .Q ( new_AGEMA_signal_14814 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6796 ( .C ( clk ), .D ( new_AGEMA_signal_14823 ), .Q ( new_AGEMA_signal_14824 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6800 ( .C ( clk ), .D ( new_AGEMA_signal_14827 ), .Q ( new_AGEMA_signal_14828 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6804 ( .C ( clk ), .D ( new_AGEMA_signal_14831 ), .Q ( new_AGEMA_signal_14832 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6808 ( .C ( clk ), .D ( new_AGEMA_signal_14835 ), .Q ( new_AGEMA_signal_14836 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6812 ( .C ( clk ), .D ( new_AGEMA_signal_14839 ), .Q ( new_AGEMA_signal_14840 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6820 ( .C ( clk ), .D ( new_AGEMA_signal_14847 ), .Q ( new_AGEMA_signal_14848 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6828 ( .C ( clk ), .D ( new_AGEMA_signal_14855 ), .Q ( new_AGEMA_signal_14856 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6836 ( .C ( clk ), .D ( new_AGEMA_signal_14863 ), .Q ( new_AGEMA_signal_14864 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6844 ( .C ( clk ), .D ( new_AGEMA_signal_14871 ), .Q ( new_AGEMA_signal_14872 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6848 ( .C ( clk ), .D ( new_AGEMA_signal_14875 ), .Q ( new_AGEMA_signal_14876 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6854 ( .C ( clk ), .D ( new_AGEMA_signal_14881 ), .Q ( new_AGEMA_signal_14882 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6860 ( .C ( clk ), .D ( new_AGEMA_signal_14887 ), .Q ( new_AGEMA_signal_14888 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6866 ( .C ( clk ), .D ( new_AGEMA_signal_14893 ), .Q ( new_AGEMA_signal_14894 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6872 ( .C ( clk ), .D ( new_AGEMA_signal_14899 ), .Q ( new_AGEMA_signal_14900 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6878 ( .C ( clk ), .D ( new_AGEMA_signal_14905 ), .Q ( new_AGEMA_signal_14906 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6884 ( .C ( clk ), .D ( new_AGEMA_signal_14911 ), .Q ( new_AGEMA_signal_14912 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6890 ( .C ( clk ), .D ( new_AGEMA_signal_14917 ), .Q ( new_AGEMA_signal_14918 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6906 ( .C ( clk ), .D ( new_AGEMA_signal_14933 ), .Q ( new_AGEMA_signal_14934 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6922 ( .C ( clk ), .D ( new_AGEMA_signal_14949 ), .Q ( new_AGEMA_signal_14950 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6938 ( .C ( clk ), .D ( new_AGEMA_signal_14965 ), .Q ( new_AGEMA_signal_14966 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6954 ( .C ( clk ), .D ( new_AGEMA_signal_14981 ), .Q ( new_AGEMA_signal_14982 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6964 ( .C ( clk ), .D ( new_AGEMA_signal_14991 ), .Q ( new_AGEMA_signal_14992 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6974 ( .C ( clk ), .D ( new_AGEMA_signal_15001 ), .Q ( new_AGEMA_signal_15002 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6984 ( .C ( clk ), .D ( new_AGEMA_signal_15011 ), .Q ( new_AGEMA_signal_15012 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6994 ( .C ( clk ), .D ( new_AGEMA_signal_15021 ), .Q ( new_AGEMA_signal_15022 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7012 ( .C ( clk ), .D ( new_AGEMA_signal_15039 ), .Q ( new_AGEMA_signal_15040 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7030 ( .C ( clk ), .D ( new_AGEMA_signal_15057 ), .Q ( new_AGEMA_signal_15058 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7048 ( .C ( clk ), .D ( new_AGEMA_signal_15075 ), .Q ( new_AGEMA_signal_15076 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7066 ( .C ( clk ), .D ( new_AGEMA_signal_15093 ), .Q ( new_AGEMA_signal_15094 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7090 ( .C ( clk ), .D ( new_AGEMA_signal_15117 ), .Q ( new_AGEMA_signal_15118 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7098 ( .C ( clk ), .D ( new_AGEMA_signal_15125 ), .Q ( new_AGEMA_signal_15126 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7106 ( .C ( clk ), .D ( new_AGEMA_signal_15133 ), .Q ( new_AGEMA_signal_15134 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7114 ( .C ( clk ), .D ( new_AGEMA_signal_15141 ), .Q ( new_AGEMA_signal_15142 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7136 ( .C ( clk ), .D ( new_AGEMA_signal_15163 ), .Q ( new_AGEMA_signal_15164 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7144 ( .C ( clk ), .D ( new_AGEMA_signal_15171 ), .Q ( new_AGEMA_signal_15172 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7152 ( .C ( clk ), .D ( new_AGEMA_signal_15179 ), .Q ( new_AGEMA_signal_15180 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7160 ( .C ( clk ), .D ( new_AGEMA_signal_15187 ), .Q ( new_AGEMA_signal_15188 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7212 ( .C ( clk ), .D ( new_AGEMA_signal_15239 ), .Q ( new_AGEMA_signal_15240 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7232 ( .C ( clk ), .D ( new_AGEMA_signal_15259 ), .Q ( new_AGEMA_signal_15260 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7252 ( .C ( clk ), .D ( new_AGEMA_signal_15279 ), .Q ( new_AGEMA_signal_15280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7272 ( .C ( clk ), .D ( new_AGEMA_signal_15299 ), .Q ( new_AGEMA_signal_15300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7314 ( .C ( clk ), .D ( new_AGEMA_signal_15341 ), .Q ( new_AGEMA_signal_15342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7326 ( .C ( clk ), .D ( new_AGEMA_signal_15353 ), .Q ( new_AGEMA_signal_15354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7338 ( .C ( clk ), .D ( new_AGEMA_signal_15365 ), .Q ( new_AGEMA_signal_15366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7350 ( .C ( clk ), .D ( new_AGEMA_signal_15377 ), .Q ( new_AGEMA_signal_15378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7362 ( .C ( clk ), .D ( new_AGEMA_signal_15389 ), .Q ( new_AGEMA_signal_15390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7376 ( .C ( clk ), .D ( new_AGEMA_signal_15403 ), .Q ( new_AGEMA_signal_15404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7390 ( .C ( clk ), .D ( new_AGEMA_signal_15417 ), .Q ( new_AGEMA_signal_15418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7404 ( .C ( clk ), .D ( new_AGEMA_signal_15431 ), .Q ( new_AGEMA_signal_15432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7416 ( .C ( clk ), .D ( new_AGEMA_signal_15443 ), .Q ( new_AGEMA_signal_15444 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7430 ( .C ( clk ), .D ( new_AGEMA_signal_15457 ), .Q ( new_AGEMA_signal_15458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7444 ( .C ( clk ), .D ( new_AGEMA_signal_15471 ), .Q ( new_AGEMA_signal_15472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7458 ( .C ( clk ), .D ( new_AGEMA_signal_15485 ), .Q ( new_AGEMA_signal_15486 ) ) ;

    /* cells in depth 21 */
    buf_clk new_AGEMA_reg_buffer_6585 ( .C ( clk ), .D ( new_AGEMA_signal_14612 ), .Q ( new_AGEMA_signal_14613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6589 ( .C ( clk ), .D ( new_AGEMA_signal_14616 ), .Q ( new_AGEMA_signal_14617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6593 ( .C ( clk ), .D ( new_AGEMA_signal_14620 ), .Q ( new_AGEMA_signal_14621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6597 ( .C ( clk ), .D ( new_AGEMA_signal_14624 ), .Q ( new_AGEMA_signal_14625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6599 ( .C ( clk ), .D ( n2109 ), .Q ( new_AGEMA_signal_14627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6601 ( .C ( clk ), .D ( new_AGEMA_signal_3582 ), .Q ( new_AGEMA_signal_14629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6603 ( .C ( clk ), .D ( new_AGEMA_signal_3583 ), .Q ( new_AGEMA_signal_14631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6605 ( .C ( clk ), .D ( new_AGEMA_signal_3584 ), .Q ( new_AGEMA_signal_14633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6621 ( .C ( clk ), .D ( new_AGEMA_signal_14648 ), .Q ( new_AGEMA_signal_14649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6637 ( .C ( clk ), .D ( new_AGEMA_signal_14664 ), .Q ( new_AGEMA_signal_14665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6653 ( .C ( clk ), .D ( new_AGEMA_signal_14680 ), .Q ( new_AGEMA_signal_14681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6669 ( .C ( clk ), .D ( new_AGEMA_signal_14696 ), .Q ( new_AGEMA_signal_14697 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6673 ( .C ( clk ), .D ( new_AGEMA_signal_14700 ), .Q ( new_AGEMA_signal_14701 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6677 ( .C ( clk ), .D ( new_AGEMA_signal_14704 ), .Q ( new_AGEMA_signal_14705 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6681 ( .C ( clk ), .D ( new_AGEMA_signal_14708 ), .Q ( new_AGEMA_signal_14709 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6685 ( .C ( clk ), .D ( new_AGEMA_signal_14712 ), .Q ( new_AGEMA_signal_14713 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6687 ( .C ( clk ), .D ( n2310 ), .Q ( new_AGEMA_signal_14715 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6689 ( .C ( clk ), .D ( new_AGEMA_signal_3597 ), .Q ( new_AGEMA_signal_14717 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6691 ( .C ( clk ), .D ( new_AGEMA_signal_3598 ), .Q ( new_AGEMA_signal_14719 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6693 ( .C ( clk ), .D ( new_AGEMA_signal_3599 ), .Q ( new_AGEMA_signal_14721 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6709 ( .C ( clk ), .D ( new_AGEMA_signal_14736 ), .Q ( new_AGEMA_signal_14737 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6725 ( .C ( clk ), .D ( new_AGEMA_signal_14752 ), .Q ( new_AGEMA_signal_14753 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6741 ( .C ( clk ), .D ( new_AGEMA_signal_14768 ), .Q ( new_AGEMA_signal_14769 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6757 ( .C ( clk ), .D ( new_AGEMA_signal_14784 ), .Q ( new_AGEMA_signal_14785 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6767 ( .C ( clk ), .D ( new_AGEMA_signal_14794 ), .Q ( new_AGEMA_signal_14795 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6777 ( .C ( clk ), .D ( new_AGEMA_signal_14804 ), .Q ( new_AGEMA_signal_14805 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6787 ( .C ( clk ), .D ( new_AGEMA_signal_14814 ), .Q ( new_AGEMA_signal_14815 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6797 ( .C ( clk ), .D ( new_AGEMA_signal_14824 ), .Q ( new_AGEMA_signal_14825 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6801 ( .C ( clk ), .D ( new_AGEMA_signal_14828 ), .Q ( new_AGEMA_signal_14829 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6805 ( .C ( clk ), .D ( new_AGEMA_signal_14832 ), .Q ( new_AGEMA_signal_14833 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6809 ( .C ( clk ), .D ( new_AGEMA_signal_14836 ), .Q ( new_AGEMA_signal_14837 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6813 ( .C ( clk ), .D ( new_AGEMA_signal_14840 ), .Q ( new_AGEMA_signal_14841 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6821 ( .C ( clk ), .D ( new_AGEMA_signal_14848 ), .Q ( new_AGEMA_signal_14849 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6829 ( .C ( clk ), .D ( new_AGEMA_signal_14856 ), .Q ( new_AGEMA_signal_14857 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6837 ( .C ( clk ), .D ( new_AGEMA_signal_14864 ), .Q ( new_AGEMA_signal_14865 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6845 ( .C ( clk ), .D ( new_AGEMA_signal_14872 ), .Q ( new_AGEMA_signal_14873 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6849 ( .C ( clk ), .D ( new_AGEMA_signal_14876 ), .Q ( new_AGEMA_signal_14877 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6855 ( .C ( clk ), .D ( new_AGEMA_signal_14882 ), .Q ( new_AGEMA_signal_14883 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6861 ( .C ( clk ), .D ( new_AGEMA_signal_14888 ), .Q ( new_AGEMA_signal_14889 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6867 ( .C ( clk ), .D ( new_AGEMA_signal_14894 ), .Q ( new_AGEMA_signal_14895 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6873 ( .C ( clk ), .D ( new_AGEMA_signal_14900 ), .Q ( new_AGEMA_signal_14901 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6879 ( .C ( clk ), .D ( new_AGEMA_signal_14906 ), .Q ( new_AGEMA_signal_14907 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6885 ( .C ( clk ), .D ( new_AGEMA_signal_14912 ), .Q ( new_AGEMA_signal_14913 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6891 ( .C ( clk ), .D ( new_AGEMA_signal_14918 ), .Q ( new_AGEMA_signal_14919 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6907 ( .C ( clk ), .D ( new_AGEMA_signal_14934 ), .Q ( new_AGEMA_signal_14935 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6923 ( .C ( clk ), .D ( new_AGEMA_signal_14950 ), .Q ( new_AGEMA_signal_14951 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6939 ( .C ( clk ), .D ( new_AGEMA_signal_14966 ), .Q ( new_AGEMA_signal_14967 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6955 ( .C ( clk ), .D ( new_AGEMA_signal_14982 ), .Q ( new_AGEMA_signal_14983 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6965 ( .C ( clk ), .D ( new_AGEMA_signal_14992 ), .Q ( new_AGEMA_signal_14993 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6975 ( .C ( clk ), .D ( new_AGEMA_signal_15002 ), .Q ( new_AGEMA_signal_15003 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6985 ( .C ( clk ), .D ( new_AGEMA_signal_15012 ), .Q ( new_AGEMA_signal_15013 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6995 ( .C ( clk ), .D ( new_AGEMA_signal_15022 ), .Q ( new_AGEMA_signal_15023 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7013 ( .C ( clk ), .D ( new_AGEMA_signal_15040 ), .Q ( new_AGEMA_signal_15041 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7031 ( .C ( clk ), .D ( new_AGEMA_signal_15058 ), .Q ( new_AGEMA_signal_15059 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7049 ( .C ( clk ), .D ( new_AGEMA_signal_15076 ), .Q ( new_AGEMA_signal_15077 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7067 ( .C ( clk ), .D ( new_AGEMA_signal_15094 ), .Q ( new_AGEMA_signal_15095 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7071 ( .C ( clk ), .D ( n2530 ), .Q ( new_AGEMA_signal_15099 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7075 ( .C ( clk ), .D ( new_AGEMA_signal_3609 ), .Q ( new_AGEMA_signal_15103 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7079 ( .C ( clk ), .D ( new_AGEMA_signal_3610 ), .Q ( new_AGEMA_signal_15107 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7083 ( .C ( clk ), .D ( new_AGEMA_signal_3611 ), .Q ( new_AGEMA_signal_15111 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7091 ( .C ( clk ), .D ( new_AGEMA_signal_15118 ), .Q ( new_AGEMA_signal_15119 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7099 ( .C ( clk ), .D ( new_AGEMA_signal_15126 ), .Q ( new_AGEMA_signal_15127 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7107 ( .C ( clk ), .D ( new_AGEMA_signal_15134 ), .Q ( new_AGEMA_signal_15135 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7115 ( .C ( clk ), .D ( new_AGEMA_signal_15142 ), .Q ( new_AGEMA_signal_15143 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7119 ( .C ( clk ), .D ( n2832 ), .Q ( new_AGEMA_signal_15147 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7123 ( .C ( clk ), .D ( new_AGEMA_signal_3618 ), .Q ( new_AGEMA_signal_15151 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7127 ( .C ( clk ), .D ( new_AGEMA_signal_3619 ), .Q ( new_AGEMA_signal_15155 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7131 ( .C ( clk ), .D ( new_AGEMA_signal_3620 ), .Q ( new_AGEMA_signal_15159 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7137 ( .C ( clk ), .D ( new_AGEMA_signal_15164 ), .Q ( new_AGEMA_signal_15165 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7145 ( .C ( clk ), .D ( new_AGEMA_signal_15172 ), .Q ( new_AGEMA_signal_15173 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7153 ( .C ( clk ), .D ( new_AGEMA_signal_15180 ), .Q ( new_AGEMA_signal_15181 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7161 ( .C ( clk ), .D ( new_AGEMA_signal_15188 ), .Q ( new_AGEMA_signal_15189 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7167 ( .C ( clk ), .D ( n2113 ), .Q ( new_AGEMA_signal_15195 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7173 ( .C ( clk ), .D ( new_AGEMA_signal_3519 ), .Q ( new_AGEMA_signal_15201 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7179 ( .C ( clk ), .D ( new_AGEMA_signal_3520 ), .Q ( new_AGEMA_signal_15207 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7185 ( .C ( clk ), .D ( new_AGEMA_signal_3521 ), .Q ( new_AGEMA_signal_15213 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7213 ( .C ( clk ), .D ( new_AGEMA_signal_15240 ), .Q ( new_AGEMA_signal_15241 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7233 ( .C ( clk ), .D ( new_AGEMA_signal_15260 ), .Q ( new_AGEMA_signal_15261 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7253 ( .C ( clk ), .D ( new_AGEMA_signal_15280 ), .Q ( new_AGEMA_signal_15281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7273 ( .C ( clk ), .D ( new_AGEMA_signal_15300 ), .Q ( new_AGEMA_signal_15301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7279 ( .C ( clk ), .D ( n2212 ), .Q ( new_AGEMA_signal_15307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7287 ( .C ( clk ), .D ( new_AGEMA_signal_3588 ), .Q ( new_AGEMA_signal_15315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7295 ( .C ( clk ), .D ( new_AGEMA_signal_3589 ), .Q ( new_AGEMA_signal_15323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7303 ( .C ( clk ), .D ( new_AGEMA_signal_3590 ), .Q ( new_AGEMA_signal_15331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7315 ( .C ( clk ), .D ( new_AGEMA_signal_15342 ), .Q ( new_AGEMA_signal_15343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7327 ( .C ( clk ), .D ( new_AGEMA_signal_15354 ), .Q ( new_AGEMA_signal_15355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7339 ( .C ( clk ), .D ( new_AGEMA_signal_15366 ), .Q ( new_AGEMA_signal_15367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7351 ( .C ( clk ), .D ( new_AGEMA_signal_15378 ), .Q ( new_AGEMA_signal_15379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7363 ( .C ( clk ), .D ( new_AGEMA_signal_15390 ), .Q ( new_AGEMA_signal_15391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7377 ( .C ( clk ), .D ( new_AGEMA_signal_15404 ), .Q ( new_AGEMA_signal_15405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7391 ( .C ( clk ), .D ( new_AGEMA_signal_15418 ), .Q ( new_AGEMA_signal_15419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7405 ( .C ( clk ), .D ( new_AGEMA_signal_15432 ), .Q ( new_AGEMA_signal_15433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7417 ( .C ( clk ), .D ( new_AGEMA_signal_15444 ), .Q ( new_AGEMA_signal_15445 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7431 ( .C ( clk ), .D ( new_AGEMA_signal_15458 ), .Q ( new_AGEMA_signal_15459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7445 ( .C ( clk ), .D ( new_AGEMA_signal_15472 ), .Q ( new_AGEMA_signal_15473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7459 ( .C ( clk ), .D ( new_AGEMA_signal_15486 ), .Q ( new_AGEMA_signal_15487 ) ) ;

    /* cells in depth 22 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2129 ( .a ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, n2000}), .b ({new_AGEMA_signal_14354, new_AGEMA_signal_14346, new_AGEMA_signal_14338, new_AGEMA_signal_14330}), .clk ( clk ), .r ({Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004]}), .c ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, n2001}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2267 ( .a ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, n2107}), .b ({new_AGEMA_signal_14402, new_AGEMA_signal_14390, new_AGEMA_signal_14378, new_AGEMA_signal_14366}), .clk ( clk ), .r ({Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, n2108}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2317 ( .a ({new_AGEMA_signal_14458, new_AGEMA_signal_14444, new_AGEMA_signal_14430, new_AGEMA_signal_14416}), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, n2149}), .clk ( clk ), .r ({Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016]}), .c ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2153}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2374 ( .a ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, n2206}), .b ({new_AGEMA_signal_14490, new_AGEMA_signal_14482, new_AGEMA_signal_14474, new_AGEMA_signal_14466}), .clk ( clk ), .r ({Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022]}), .c ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633, n2207}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2477 ( .a ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, n2308}), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, n2307}), .clk ( clk ), .r ({Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028]}), .c ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, n2309}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2535 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, n2370}), .b ({new_AGEMA_signal_14546, new_AGEMA_signal_14532, new_AGEMA_signal_14518, new_AGEMA_signal_14504}), .clk ( clk ), .r ({Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, n2373}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2661 ( .a ({new_AGEMA_signal_14578, new_AGEMA_signal_14570, new_AGEMA_signal_14562, new_AGEMA_signal_14554}), .b ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, n2515}), .clk ( clk ), .r ({Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040]}), .c ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2528}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2750 ( .a ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, new_AGEMA_signal_3615, n2639}), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, n2638}), .clk ( clk ), .r ({Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046]}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645, n2669}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2843 ( .a ({new_AGEMA_signal_14610, new_AGEMA_signal_14602, new_AGEMA_signal_14594, new_AGEMA_signal_14586}), .b ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, n2807}), .clk ( clk ), .r ({Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052]}), .c ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621, n2830}) ) ;
    buf_clk new_AGEMA_reg_buffer_6586 ( .C ( clk ), .D ( new_AGEMA_signal_14613 ), .Q ( new_AGEMA_signal_14614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6590 ( .C ( clk ), .D ( new_AGEMA_signal_14617 ), .Q ( new_AGEMA_signal_14618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6594 ( .C ( clk ), .D ( new_AGEMA_signal_14621 ), .Q ( new_AGEMA_signal_14622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6598 ( .C ( clk ), .D ( new_AGEMA_signal_14625 ), .Q ( new_AGEMA_signal_14626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6600 ( .C ( clk ), .D ( new_AGEMA_signal_14627 ), .Q ( new_AGEMA_signal_14628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6602 ( .C ( clk ), .D ( new_AGEMA_signal_14629 ), .Q ( new_AGEMA_signal_14630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6604 ( .C ( clk ), .D ( new_AGEMA_signal_14631 ), .Q ( new_AGEMA_signal_14632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6606 ( .C ( clk ), .D ( new_AGEMA_signal_14633 ), .Q ( new_AGEMA_signal_14634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6622 ( .C ( clk ), .D ( new_AGEMA_signal_14649 ), .Q ( new_AGEMA_signal_14650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6638 ( .C ( clk ), .D ( new_AGEMA_signal_14665 ), .Q ( new_AGEMA_signal_14666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6654 ( .C ( clk ), .D ( new_AGEMA_signal_14681 ), .Q ( new_AGEMA_signal_14682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6670 ( .C ( clk ), .D ( new_AGEMA_signal_14697 ), .Q ( new_AGEMA_signal_14698 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6674 ( .C ( clk ), .D ( new_AGEMA_signal_14701 ), .Q ( new_AGEMA_signal_14702 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6678 ( .C ( clk ), .D ( new_AGEMA_signal_14705 ), .Q ( new_AGEMA_signal_14706 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6682 ( .C ( clk ), .D ( new_AGEMA_signal_14709 ), .Q ( new_AGEMA_signal_14710 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6686 ( .C ( clk ), .D ( new_AGEMA_signal_14713 ), .Q ( new_AGEMA_signal_14714 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6688 ( .C ( clk ), .D ( new_AGEMA_signal_14715 ), .Q ( new_AGEMA_signal_14716 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6690 ( .C ( clk ), .D ( new_AGEMA_signal_14717 ), .Q ( new_AGEMA_signal_14718 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6692 ( .C ( clk ), .D ( new_AGEMA_signal_14719 ), .Q ( new_AGEMA_signal_14720 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6694 ( .C ( clk ), .D ( new_AGEMA_signal_14721 ), .Q ( new_AGEMA_signal_14722 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6710 ( .C ( clk ), .D ( new_AGEMA_signal_14737 ), .Q ( new_AGEMA_signal_14738 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6726 ( .C ( clk ), .D ( new_AGEMA_signal_14753 ), .Q ( new_AGEMA_signal_14754 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6742 ( .C ( clk ), .D ( new_AGEMA_signal_14769 ), .Q ( new_AGEMA_signal_14770 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6758 ( .C ( clk ), .D ( new_AGEMA_signal_14785 ), .Q ( new_AGEMA_signal_14786 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6768 ( .C ( clk ), .D ( new_AGEMA_signal_14795 ), .Q ( new_AGEMA_signal_14796 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6778 ( .C ( clk ), .D ( new_AGEMA_signal_14805 ), .Q ( new_AGEMA_signal_14806 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6788 ( .C ( clk ), .D ( new_AGEMA_signal_14815 ), .Q ( new_AGEMA_signal_14816 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6798 ( .C ( clk ), .D ( new_AGEMA_signal_14825 ), .Q ( new_AGEMA_signal_14826 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6802 ( .C ( clk ), .D ( new_AGEMA_signal_14829 ), .Q ( new_AGEMA_signal_14830 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6806 ( .C ( clk ), .D ( new_AGEMA_signal_14833 ), .Q ( new_AGEMA_signal_14834 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6810 ( .C ( clk ), .D ( new_AGEMA_signal_14837 ), .Q ( new_AGEMA_signal_14838 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6814 ( .C ( clk ), .D ( new_AGEMA_signal_14841 ), .Q ( new_AGEMA_signal_14842 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6822 ( .C ( clk ), .D ( new_AGEMA_signal_14849 ), .Q ( new_AGEMA_signal_14850 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6830 ( .C ( clk ), .D ( new_AGEMA_signal_14857 ), .Q ( new_AGEMA_signal_14858 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6838 ( .C ( clk ), .D ( new_AGEMA_signal_14865 ), .Q ( new_AGEMA_signal_14866 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6846 ( .C ( clk ), .D ( new_AGEMA_signal_14873 ), .Q ( new_AGEMA_signal_14874 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6850 ( .C ( clk ), .D ( new_AGEMA_signal_14877 ), .Q ( new_AGEMA_signal_14878 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6856 ( .C ( clk ), .D ( new_AGEMA_signal_14883 ), .Q ( new_AGEMA_signal_14884 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6862 ( .C ( clk ), .D ( new_AGEMA_signal_14889 ), .Q ( new_AGEMA_signal_14890 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6868 ( .C ( clk ), .D ( new_AGEMA_signal_14895 ), .Q ( new_AGEMA_signal_14896 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6874 ( .C ( clk ), .D ( new_AGEMA_signal_14901 ), .Q ( new_AGEMA_signal_14902 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6880 ( .C ( clk ), .D ( new_AGEMA_signal_14907 ), .Q ( new_AGEMA_signal_14908 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6886 ( .C ( clk ), .D ( new_AGEMA_signal_14913 ), .Q ( new_AGEMA_signal_14914 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6892 ( .C ( clk ), .D ( new_AGEMA_signal_14919 ), .Q ( new_AGEMA_signal_14920 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6908 ( .C ( clk ), .D ( new_AGEMA_signal_14935 ), .Q ( new_AGEMA_signal_14936 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6924 ( .C ( clk ), .D ( new_AGEMA_signal_14951 ), .Q ( new_AGEMA_signal_14952 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6940 ( .C ( clk ), .D ( new_AGEMA_signal_14967 ), .Q ( new_AGEMA_signal_14968 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6956 ( .C ( clk ), .D ( new_AGEMA_signal_14983 ), .Q ( new_AGEMA_signal_14984 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6966 ( .C ( clk ), .D ( new_AGEMA_signal_14993 ), .Q ( new_AGEMA_signal_14994 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6976 ( .C ( clk ), .D ( new_AGEMA_signal_15003 ), .Q ( new_AGEMA_signal_15004 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6986 ( .C ( clk ), .D ( new_AGEMA_signal_15013 ), .Q ( new_AGEMA_signal_15014 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6996 ( .C ( clk ), .D ( new_AGEMA_signal_15023 ), .Q ( new_AGEMA_signal_15024 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7014 ( .C ( clk ), .D ( new_AGEMA_signal_15041 ), .Q ( new_AGEMA_signal_15042 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7032 ( .C ( clk ), .D ( new_AGEMA_signal_15059 ), .Q ( new_AGEMA_signal_15060 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7050 ( .C ( clk ), .D ( new_AGEMA_signal_15077 ), .Q ( new_AGEMA_signal_15078 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7068 ( .C ( clk ), .D ( new_AGEMA_signal_15095 ), .Q ( new_AGEMA_signal_15096 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7072 ( .C ( clk ), .D ( new_AGEMA_signal_15099 ), .Q ( new_AGEMA_signal_15100 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7076 ( .C ( clk ), .D ( new_AGEMA_signal_15103 ), .Q ( new_AGEMA_signal_15104 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7080 ( .C ( clk ), .D ( new_AGEMA_signal_15107 ), .Q ( new_AGEMA_signal_15108 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7084 ( .C ( clk ), .D ( new_AGEMA_signal_15111 ), .Q ( new_AGEMA_signal_15112 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7092 ( .C ( clk ), .D ( new_AGEMA_signal_15119 ), .Q ( new_AGEMA_signal_15120 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7100 ( .C ( clk ), .D ( new_AGEMA_signal_15127 ), .Q ( new_AGEMA_signal_15128 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7108 ( .C ( clk ), .D ( new_AGEMA_signal_15135 ), .Q ( new_AGEMA_signal_15136 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7116 ( .C ( clk ), .D ( new_AGEMA_signal_15143 ), .Q ( new_AGEMA_signal_15144 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7120 ( .C ( clk ), .D ( new_AGEMA_signal_15147 ), .Q ( new_AGEMA_signal_15148 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7124 ( .C ( clk ), .D ( new_AGEMA_signal_15151 ), .Q ( new_AGEMA_signal_15152 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7128 ( .C ( clk ), .D ( new_AGEMA_signal_15155 ), .Q ( new_AGEMA_signal_15156 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7132 ( .C ( clk ), .D ( new_AGEMA_signal_15159 ), .Q ( new_AGEMA_signal_15160 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7138 ( .C ( clk ), .D ( new_AGEMA_signal_15165 ), .Q ( new_AGEMA_signal_15166 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7146 ( .C ( clk ), .D ( new_AGEMA_signal_15173 ), .Q ( new_AGEMA_signal_15174 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7154 ( .C ( clk ), .D ( new_AGEMA_signal_15181 ), .Q ( new_AGEMA_signal_15182 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7162 ( .C ( clk ), .D ( new_AGEMA_signal_15189 ), .Q ( new_AGEMA_signal_15190 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7168 ( .C ( clk ), .D ( new_AGEMA_signal_15195 ), .Q ( new_AGEMA_signal_15196 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7174 ( .C ( clk ), .D ( new_AGEMA_signal_15201 ), .Q ( new_AGEMA_signal_15202 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7180 ( .C ( clk ), .D ( new_AGEMA_signal_15207 ), .Q ( new_AGEMA_signal_15208 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7186 ( .C ( clk ), .D ( new_AGEMA_signal_15213 ), .Q ( new_AGEMA_signal_15214 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7214 ( .C ( clk ), .D ( new_AGEMA_signal_15241 ), .Q ( new_AGEMA_signal_15242 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7234 ( .C ( clk ), .D ( new_AGEMA_signal_15261 ), .Q ( new_AGEMA_signal_15262 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7254 ( .C ( clk ), .D ( new_AGEMA_signal_15281 ), .Q ( new_AGEMA_signal_15282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7274 ( .C ( clk ), .D ( new_AGEMA_signal_15301 ), .Q ( new_AGEMA_signal_15302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7280 ( .C ( clk ), .D ( new_AGEMA_signal_15307 ), .Q ( new_AGEMA_signal_15308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7288 ( .C ( clk ), .D ( new_AGEMA_signal_15315 ), .Q ( new_AGEMA_signal_15316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7296 ( .C ( clk ), .D ( new_AGEMA_signal_15323 ), .Q ( new_AGEMA_signal_15324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7304 ( .C ( clk ), .D ( new_AGEMA_signal_15331 ), .Q ( new_AGEMA_signal_15332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7316 ( .C ( clk ), .D ( new_AGEMA_signal_15343 ), .Q ( new_AGEMA_signal_15344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7328 ( .C ( clk ), .D ( new_AGEMA_signal_15355 ), .Q ( new_AGEMA_signal_15356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7340 ( .C ( clk ), .D ( new_AGEMA_signal_15367 ), .Q ( new_AGEMA_signal_15368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7352 ( .C ( clk ), .D ( new_AGEMA_signal_15379 ), .Q ( new_AGEMA_signal_15380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7364 ( .C ( clk ), .D ( new_AGEMA_signal_15391 ), .Q ( new_AGEMA_signal_15392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7378 ( .C ( clk ), .D ( new_AGEMA_signal_15405 ), .Q ( new_AGEMA_signal_15406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7392 ( .C ( clk ), .D ( new_AGEMA_signal_15419 ), .Q ( new_AGEMA_signal_15420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7406 ( .C ( clk ), .D ( new_AGEMA_signal_15433 ), .Q ( new_AGEMA_signal_15434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7418 ( .C ( clk ), .D ( new_AGEMA_signal_15445 ), .Q ( new_AGEMA_signal_15446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7432 ( .C ( clk ), .D ( new_AGEMA_signal_15459 ), .Q ( new_AGEMA_signal_15460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7446 ( .C ( clk ), .D ( new_AGEMA_signal_15473 ), .Q ( new_AGEMA_signal_15474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7460 ( .C ( clk ), .D ( new_AGEMA_signal_15487 ), .Q ( new_AGEMA_signal_15488 ) ) ;

    /* cells in depth 23 */
    buf_clk new_AGEMA_reg_buffer_6851 ( .C ( clk ), .D ( new_AGEMA_signal_14878 ), .Q ( new_AGEMA_signal_14879 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6857 ( .C ( clk ), .D ( new_AGEMA_signal_14884 ), .Q ( new_AGEMA_signal_14885 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6863 ( .C ( clk ), .D ( new_AGEMA_signal_14890 ), .Q ( new_AGEMA_signal_14891 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6869 ( .C ( clk ), .D ( new_AGEMA_signal_14896 ), .Q ( new_AGEMA_signal_14897 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6875 ( .C ( clk ), .D ( new_AGEMA_signal_14902 ), .Q ( new_AGEMA_signal_14903 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6881 ( .C ( clk ), .D ( new_AGEMA_signal_14908 ), .Q ( new_AGEMA_signal_14909 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6887 ( .C ( clk ), .D ( new_AGEMA_signal_14914 ), .Q ( new_AGEMA_signal_14915 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6893 ( .C ( clk ), .D ( new_AGEMA_signal_14920 ), .Q ( new_AGEMA_signal_14921 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6909 ( .C ( clk ), .D ( new_AGEMA_signal_14936 ), .Q ( new_AGEMA_signal_14937 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6925 ( .C ( clk ), .D ( new_AGEMA_signal_14952 ), .Q ( new_AGEMA_signal_14953 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6941 ( .C ( clk ), .D ( new_AGEMA_signal_14968 ), .Q ( new_AGEMA_signal_14969 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6957 ( .C ( clk ), .D ( new_AGEMA_signal_14984 ), .Q ( new_AGEMA_signal_14985 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6967 ( .C ( clk ), .D ( new_AGEMA_signal_14994 ), .Q ( new_AGEMA_signal_14995 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6977 ( .C ( clk ), .D ( new_AGEMA_signal_15004 ), .Q ( new_AGEMA_signal_15005 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6987 ( .C ( clk ), .D ( new_AGEMA_signal_15014 ), .Q ( new_AGEMA_signal_15015 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6997 ( .C ( clk ), .D ( new_AGEMA_signal_15024 ), .Q ( new_AGEMA_signal_15025 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7015 ( .C ( clk ), .D ( new_AGEMA_signal_15042 ), .Q ( new_AGEMA_signal_15043 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7033 ( .C ( clk ), .D ( new_AGEMA_signal_15060 ), .Q ( new_AGEMA_signal_15061 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7051 ( .C ( clk ), .D ( new_AGEMA_signal_15078 ), .Q ( new_AGEMA_signal_15079 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7069 ( .C ( clk ), .D ( new_AGEMA_signal_15096 ), .Q ( new_AGEMA_signal_15097 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7073 ( .C ( clk ), .D ( new_AGEMA_signal_15100 ), .Q ( new_AGEMA_signal_15101 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7077 ( .C ( clk ), .D ( new_AGEMA_signal_15104 ), .Q ( new_AGEMA_signal_15105 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7081 ( .C ( clk ), .D ( new_AGEMA_signal_15108 ), .Q ( new_AGEMA_signal_15109 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7085 ( .C ( clk ), .D ( new_AGEMA_signal_15112 ), .Q ( new_AGEMA_signal_15113 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7093 ( .C ( clk ), .D ( new_AGEMA_signal_15120 ), .Q ( new_AGEMA_signal_15121 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7101 ( .C ( clk ), .D ( new_AGEMA_signal_15128 ), .Q ( new_AGEMA_signal_15129 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7109 ( .C ( clk ), .D ( new_AGEMA_signal_15136 ), .Q ( new_AGEMA_signal_15137 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7117 ( .C ( clk ), .D ( new_AGEMA_signal_15144 ), .Q ( new_AGEMA_signal_15145 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7121 ( .C ( clk ), .D ( new_AGEMA_signal_15148 ), .Q ( new_AGEMA_signal_15149 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7125 ( .C ( clk ), .D ( new_AGEMA_signal_15152 ), .Q ( new_AGEMA_signal_15153 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7129 ( .C ( clk ), .D ( new_AGEMA_signal_15156 ), .Q ( new_AGEMA_signal_15157 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7133 ( .C ( clk ), .D ( new_AGEMA_signal_15160 ), .Q ( new_AGEMA_signal_15161 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7139 ( .C ( clk ), .D ( new_AGEMA_signal_15166 ), .Q ( new_AGEMA_signal_15167 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7147 ( .C ( clk ), .D ( new_AGEMA_signal_15174 ), .Q ( new_AGEMA_signal_15175 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7155 ( .C ( clk ), .D ( new_AGEMA_signal_15182 ), .Q ( new_AGEMA_signal_15183 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7163 ( .C ( clk ), .D ( new_AGEMA_signal_15190 ), .Q ( new_AGEMA_signal_15191 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7169 ( .C ( clk ), .D ( new_AGEMA_signal_15196 ), .Q ( new_AGEMA_signal_15197 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7175 ( .C ( clk ), .D ( new_AGEMA_signal_15202 ), .Q ( new_AGEMA_signal_15203 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7181 ( .C ( clk ), .D ( new_AGEMA_signal_15208 ), .Q ( new_AGEMA_signal_15209 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7187 ( .C ( clk ), .D ( new_AGEMA_signal_15214 ), .Q ( new_AGEMA_signal_15215 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7215 ( .C ( clk ), .D ( new_AGEMA_signal_15242 ), .Q ( new_AGEMA_signal_15243 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7235 ( .C ( clk ), .D ( new_AGEMA_signal_15262 ), .Q ( new_AGEMA_signal_15263 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7255 ( .C ( clk ), .D ( new_AGEMA_signal_15282 ), .Q ( new_AGEMA_signal_15283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7275 ( .C ( clk ), .D ( new_AGEMA_signal_15302 ), .Q ( new_AGEMA_signal_15303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7281 ( .C ( clk ), .D ( new_AGEMA_signal_15308 ), .Q ( new_AGEMA_signal_15309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7289 ( .C ( clk ), .D ( new_AGEMA_signal_15316 ), .Q ( new_AGEMA_signal_15317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7297 ( .C ( clk ), .D ( new_AGEMA_signal_15324 ), .Q ( new_AGEMA_signal_15325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7305 ( .C ( clk ), .D ( new_AGEMA_signal_15332 ), .Q ( new_AGEMA_signal_15333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7317 ( .C ( clk ), .D ( new_AGEMA_signal_15344 ), .Q ( new_AGEMA_signal_15345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7329 ( .C ( clk ), .D ( new_AGEMA_signal_15356 ), .Q ( new_AGEMA_signal_15357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7341 ( .C ( clk ), .D ( new_AGEMA_signal_15368 ), .Q ( new_AGEMA_signal_15369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7353 ( .C ( clk ), .D ( new_AGEMA_signal_15380 ), .Q ( new_AGEMA_signal_15381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7365 ( .C ( clk ), .D ( new_AGEMA_signal_15392 ), .Q ( new_AGEMA_signal_15393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7379 ( .C ( clk ), .D ( new_AGEMA_signal_15406 ), .Q ( new_AGEMA_signal_15407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7393 ( .C ( clk ), .D ( new_AGEMA_signal_15420 ), .Q ( new_AGEMA_signal_15421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7407 ( .C ( clk ), .D ( new_AGEMA_signal_15434 ), .Q ( new_AGEMA_signal_15435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7419 ( .C ( clk ), .D ( new_AGEMA_signal_15446 ), .Q ( new_AGEMA_signal_15447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7433 ( .C ( clk ), .D ( new_AGEMA_signal_15460 ), .Q ( new_AGEMA_signal_15461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7447 ( .C ( clk ), .D ( new_AGEMA_signal_15474 ), .Q ( new_AGEMA_signal_15475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7461 ( .C ( clk ), .D ( new_AGEMA_signal_15488 ), .Q ( new_AGEMA_signal_15489 ) ) ;

    /* cells in depth 24 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2130 ( .a ({new_AGEMA_signal_14626, new_AGEMA_signal_14622, new_AGEMA_signal_14618, new_AGEMA_signal_14614}), .b ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, n2001}), .clk ( clk ), .r ({Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058]}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, n2017}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2268 ( .a ({new_AGEMA_signal_14634, new_AGEMA_signal_14632, new_AGEMA_signal_14630, new_AGEMA_signal_14628}), .b ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, new_AGEMA_signal_3627, n2108}), .clk ( clk ), .r ({Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064]}), .c ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2110}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2319 ( .a ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, n2153}), .b ({new_AGEMA_signal_14698, new_AGEMA_signal_14682, new_AGEMA_signal_14666, new_AGEMA_signal_14650}), .clk ( clk ), .r ({Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070]}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657, n2154}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2375 ( .a ({new_AGEMA_signal_14714, new_AGEMA_signal_14710, new_AGEMA_signal_14706, new_AGEMA_signal_14702}), .b ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, new_AGEMA_signal_3633, n2207}), .clk ( clk ), .r ({Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076]}), .c ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, n2209}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2478 ( .a ({new_AGEMA_signal_14722, new_AGEMA_signal_14720, new_AGEMA_signal_14718, new_AGEMA_signal_14716}), .b ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, n2309}), .clk ( clk ), .r ({Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082]}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, n2311}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2537 ( .a ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, new_AGEMA_signal_3639, n2373}), .b ({new_AGEMA_signal_14786, new_AGEMA_signal_14770, new_AGEMA_signal_14754, new_AGEMA_signal_14738}), .clk ( clk ), .r ({Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088]}), .c ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2374}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2672 ( .a ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, n2528}), .b ({new_AGEMA_signal_14826, new_AGEMA_signal_14816, new_AGEMA_signal_14806, new_AGEMA_signal_14796}), .clk ( clk ), .r ({Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094]}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669, n2529}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2768 ( .a ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, new_AGEMA_signal_3645, n2669}), .b ({new_AGEMA_signal_14842, new_AGEMA_signal_14838, new_AGEMA_signal_14834, new_AGEMA_signal_14830}), .clk ( clk ), .r ({Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100]}), .c ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, n2670}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2854 ( .a ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, new_AGEMA_signal_3621, n2830}), .b ({new_AGEMA_signal_14874, new_AGEMA_signal_14866, new_AGEMA_signal_14858, new_AGEMA_signal_14850}), .clk ( clk ), .r ({Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106]}), .c ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, n2831}) ) ;
    buf_clk new_AGEMA_reg_buffer_6852 ( .C ( clk ), .D ( new_AGEMA_signal_14879 ), .Q ( new_AGEMA_signal_14880 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6858 ( .C ( clk ), .D ( new_AGEMA_signal_14885 ), .Q ( new_AGEMA_signal_14886 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6864 ( .C ( clk ), .D ( new_AGEMA_signal_14891 ), .Q ( new_AGEMA_signal_14892 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6870 ( .C ( clk ), .D ( new_AGEMA_signal_14897 ), .Q ( new_AGEMA_signal_14898 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6876 ( .C ( clk ), .D ( new_AGEMA_signal_14903 ), .Q ( new_AGEMA_signal_14904 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6882 ( .C ( clk ), .D ( new_AGEMA_signal_14909 ), .Q ( new_AGEMA_signal_14910 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6888 ( .C ( clk ), .D ( new_AGEMA_signal_14915 ), .Q ( new_AGEMA_signal_14916 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6894 ( .C ( clk ), .D ( new_AGEMA_signal_14921 ), .Q ( new_AGEMA_signal_14922 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6910 ( .C ( clk ), .D ( new_AGEMA_signal_14937 ), .Q ( new_AGEMA_signal_14938 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6926 ( .C ( clk ), .D ( new_AGEMA_signal_14953 ), .Q ( new_AGEMA_signal_14954 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6942 ( .C ( clk ), .D ( new_AGEMA_signal_14969 ), .Q ( new_AGEMA_signal_14970 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6958 ( .C ( clk ), .D ( new_AGEMA_signal_14985 ), .Q ( new_AGEMA_signal_14986 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6968 ( .C ( clk ), .D ( new_AGEMA_signal_14995 ), .Q ( new_AGEMA_signal_14996 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6978 ( .C ( clk ), .D ( new_AGEMA_signal_15005 ), .Q ( new_AGEMA_signal_15006 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6988 ( .C ( clk ), .D ( new_AGEMA_signal_15015 ), .Q ( new_AGEMA_signal_15016 ) ) ;
    buf_clk new_AGEMA_reg_buffer_6998 ( .C ( clk ), .D ( new_AGEMA_signal_15025 ), .Q ( new_AGEMA_signal_15026 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7016 ( .C ( clk ), .D ( new_AGEMA_signal_15043 ), .Q ( new_AGEMA_signal_15044 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7034 ( .C ( clk ), .D ( new_AGEMA_signal_15061 ), .Q ( new_AGEMA_signal_15062 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7052 ( .C ( clk ), .D ( new_AGEMA_signal_15079 ), .Q ( new_AGEMA_signal_15080 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7070 ( .C ( clk ), .D ( new_AGEMA_signal_15097 ), .Q ( new_AGEMA_signal_15098 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7074 ( .C ( clk ), .D ( new_AGEMA_signal_15101 ), .Q ( new_AGEMA_signal_15102 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7078 ( .C ( clk ), .D ( new_AGEMA_signal_15105 ), .Q ( new_AGEMA_signal_15106 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7082 ( .C ( clk ), .D ( new_AGEMA_signal_15109 ), .Q ( new_AGEMA_signal_15110 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7086 ( .C ( clk ), .D ( new_AGEMA_signal_15113 ), .Q ( new_AGEMA_signal_15114 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7094 ( .C ( clk ), .D ( new_AGEMA_signal_15121 ), .Q ( new_AGEMA_signal_15122 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7102 ( .C ( clk ), .D ( new_AGEMA_signal_15129 ), .Q ( new_AGEMA_signal_15130 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7110 ( .C ( clk ), .D ( new_AGEMA_signal_15137 ), .Q ( new_AGEMA_signal_15138 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7118 ( .C ( clk ), .D ( new_AGEMA_signal_15145 ), .Q ( new_AGEMA_signal_15146 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7122 ( .C ( clk ), .D ( new_AGEMA_signal_15149 ), .Q ( new_AGEMA_signal_15150 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7126 ( .C ( clk ), .D ( new_AGEMA_signal_15153 ), .Q ( new_AGEMA_signal_15154 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7130 ( .C ( clk ), .D ( new_AGEMA_signal_15157 ), .Q ( new_AGEMA_signal_15158 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7134 ( .C ( clk ), .D ( new_AGEMA_signal_15161 ), .Q ( new_AGEMA_signal_15162 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7140 ( .C ( clk ), .D ( new_AGEMA_signal_15167 ), .Q ( new_AGEMA_signal_15168 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7148 ( .C ( clk ), .D ( new_AGEMA_signal_15175 ), .Q ( new_AGEMA_signal_15176 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7156 ( .C ( clk ), .D ( new_AGEMA_signal_15183 ), .Q ( new_AGEMA_signal_15184 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7164 ( .C ( clk ), .D ( new_AGEMA_signal_15191 ), .Q ( new_AGEMA_signal_15192 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7170 ( .C ( clk ), .D ( new_AGEMA_signal_15197 ), .Q ( new_AGEMA_signal_15198 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7176 ( .C ( clk ), .D ( new_AGEMA_signal_15203 ), .Q ( new_AGEMA_signal_15204 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7182 ( .C ( clk ), .D ( new_AGEMA_signal_15209 ), .Q ( new_AGEMA_signal_15210 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7188 ( .C ( clk ), .D ( new_AGEMA_signal_15215 ), .Q ( new_AGEMA_signal_15216 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7216 ( .C ( clk ), .D ( new_AGEMA_signal_15243 ), .Q ( new_AGEMA_signal_15244 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7236 ( .C ( clk ), .D ( new_AGEMA_signal_15263 ), .Q ( new_AGEMA_signal_15264 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7256 ( .C ( clk ), .D ( new_AGEMA_signal_15283 ), .Q ( new_AGEMA_signal_15284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7276 ( .C ( clk ), .D ( new_AGEMA_signal_15303 ), .Q ( new_AGEMA_signal_15304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7282 ( .C ( clk ), .D ( new_AGEMA_signal_15309 ), .Q ( new_AGEMA_signal_15310 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7290 ( .C ( clk ), .D ( new_AGEMA_signal_15317 ), .Q ( new_AGEMA_signal_15318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7298 ( .C ( clk ), .D ( new_AGEMA_signal_15325 ), .Q ( new_AGEMA_signal_15326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7306 ( .C ( clk ), .D ( new_AGEMA_signal_15333 ), .Q ( new_AGEMA_signal_15334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7318 ( .C ( clk ), .D ( new_AGEMA_signal_15345 ), .Q ( new_AGEMA_signal_15346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7330 ( .C ( clk ), .D ( new_AGEMA_signal_15357 ), .Q ( new_AGEMA_signal_15358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7342 ( .C ( clk ), .D ( new_AGEMA_signal_15369 ), .Q ( new_AGEMA_signal_15370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7354 ( .C ( clk ), .D ( new_AGEMA_signal_15381 ), .Q ( new_AGEMA_signal_15382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7366 ( .C ( clk ), .D ( new_AGEMA_signal_15393 ), .Q ( new_AGEMA_signal_15394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7380 ( .C ( clk ), .D ( new_AGEMA_signal_15407 ), .Q ( new_AGEMA_signal_15408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7394 ( .C ( clk ), .D ( new_AGEMA_signal_15421 ), .Q ( new_AGEMA_signal_15422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7408 ( .C ( clk ), .D ( new_AGEMA_signal_15435 ), .Q ( new_AGEMA_signal_15436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7420 ( .C ( clk ), .D ( new_AGEMA_signal_15447 ), .Q ( new_AGEMA_signal_15448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7434 ( .C ( clk ), .D ( new_AGEMA_signal_15461 ), .Q ( new_AGEMA_signal_15462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7448 ( .C ( clk ), .D ( new_AGEMA_signal_15475 ), .Q ( new_AGEMA_signal_15476 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7462 ( .C ( clk ), .D ( new_AGEMA_signal_15489 ), .Q ( new_AGEMA_signal_15490 ) ) ;

    /* cells in depth 25 */
    buf_clk new_AGEMA_reg_buffer_7141 ( .C ( clk ), .D ( new_AGEMA_signal_15168 ), .Q ( new_AGEMA_signal_15169 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7149 ( .C ( clk ), .D ( new_AGEMA_signal_15176 ), .Q ( new_AGEMA_signal_15177 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7157 ( .C ( clk ), .D ( new_AGEMA_signal_15184 ), .Q ( new_AGEMA_signal_15185 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7165 ( .C ( clk ), .D ( new_AGEMA_signal_15192 ), .Q ( new_AGEMA_signal_15193 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7171 ( .C ( clk ), .D ( new_AGEMA_signal_15198 ), .Q ( new_AGEMA_signal_15199 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7177 ( .C ( clk ), .D ( new_AGEMA_signal_15204 ), .Q ( new_AGEMA_signal_15205 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7183 ( .C ( clk ), .D ( new_AGEMA_signal_15210 ), .Q ( new_AGEMA_signal_15211 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7189 ( .C ( clk ), .D ( new_AGEMA_signal_15216 ), .Q ( new_AGEMA_signal_15217 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7191 ( .C ( clk ), .D ( n2209 ), .Q ( new_AGEMA_signal_15219 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7193 ( .C ( clk ), .D ( new_AGEMA_signal_3660 ), .Q ( new_AGEMA_signal_15221 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7195 ( .C ( clk ), .D ( new_AGEMA_signal_3661 ), .Q ( new_AGEMA_signal_15223 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7197 ( .C ( clk ), .D ( new_AGEMA_signal_3662 ), .Q ( new_AGEMA_signal_15225 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7217 ( .C ( clk ), .D ( new_AGEMA_signal_15244 ), .Q ( new_AGEMA_signal_15245 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7237 ( .C ( clk ), .D ( new_AGEMA_signal_15264 ), .Q ( new_AGEMA_signal_15265 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7257 ( .C ( clk ), .D ( new_AGEMA_signal_15284 ), .Q ( new_AGEMA_signal_15285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7277 ( .C ( clk ), .D ( new_AGEMA_signal_15304 ), .Q ( new_AGEMA_signal_15305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7283 ( .C ( clk ), .D ( new_AGEMA_signal_15310 ), .Q ( new_AGEMA_signal_15311 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7291 ( .C ( clk ), .D ( new_AGEMA_signal_15318 ), .Q ( new_AGEMA_signal_15319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7299 ( .C ( clk ), .D ( new_AGEMA_signal_15326 ), .Q ( new_AGEMA_signal_15327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7307 ( .C ( clk ), .D ( new_AGEMA_signal_15334 ), .Q ( new_AGEMA_signal_15335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7319 ( .C ( clk ), .D ( new_AGEMA_signal_15346 ), .Q ( new_AGEMA_signal_15347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7331 ( .C ( clk ), .D ( new_AGEMA_signal_15358 ), .Q ( new_AGEMA_signal_15359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7343 ( .C ( clk ), .D ( new_AGEMA_signal_15370 ), .Q ( new_AGEMA_signal_15371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7355 ( .C ( clk ), .D ( new_AGEMA_signal_15382 ), .Q ( new_AGEMA_signal_15383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7367 ( .C ( clk ), .D ( new_AGEMA_signal_15394 ), .Q ( new_AGEMA_signal_15395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7381 ( .C ( clk ), .D ( new_AGEMA_signal_15408 ), .Q ( new_AGEMA_signal_15409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7395 ( .C ( clk ), .D ( new_AGEMA_signal_15422 ), .Q ( new_AGEMA_signal_15423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7409 ( .C ( clk ), .D ( new_AGEMA_signal_15436 ), .Q ( new_AGEMA_signal_15437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7421 ( .C ( clk ), .D ( new_AGEMA_signal_15448 ), .Q ( new_AGEMA_signal_15449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7435 ( .C ( clk ), .D ( new_AGEMA_signal_15462 ), .Q ( new_AGEMA_signal_15463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7449 ( .C ( clk ), .D ( new_AGEMA_signal_15476 ), .Q ( new_AGEMA_signal_15477 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7463 ( .C ( clk ), .D ( new_AGEMA_signal_15490 ), .Q ( new_AGEMA_signal_15491 ) ) ;

    /* cells in depth 26 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2155 ( .a ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, new_AGEMA_signal_3651, n2017}), .b ({new_AGEMA_signal_14898, new_AGEMA_signal_14892, new_AGEMA_signal_14886, new_AGEMA_signal_14880}), .clk ( clk ), .r ({Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112]}), .c ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2018}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2269 ( .a ({new_AGEMA_signal_14922, new_AGEMA_signal_14916, new_AGEMA_signal_14910, new_AGEMA_signal_14904}), .b ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, n2110}), .clk ( clk ), .r ({Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118]}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681, n2112}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2320 ( .a ({new_AGEMA_signal_14986, new_AGEMA_signal_14970, new_AGEMA_signal_14954, new_AGEMA_signal_14938}), .b ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, new_AGEMA_signal_3657, n2154}), .clk ( clk ), .r ({Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124]}), .c ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, n2210}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2479 ( .a ({new_AGEMA_signal_15026, new_AGEMA_signal_15016, new_AGEMA_signal_15006, new_AGEMA_signal_14996}), .b ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, new_AGEMA_signal_3663, n2311}), .clk ( clk ), .r ({Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130]}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, new_AGEMA_signal_3687, N470}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2538 ( .a ({new_AGEMA_signal_15098, new_AGEMA_signal_15080, new_AGEMA_signal_15062, new_AGEMA_signal_15044}), .b ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, n2374}), .clk ( clk ), .r ({Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136]}), .c ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2378}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2673 ( .a ({new_AGEMA_signal_15114, new_AGEMA_signal_15110, new_AGEMA_signal_15106, new_AGEMA_signal_15102}), .b ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, new_AGEMA_signal_3669, n2529}), .clk ( clk ), .r ({Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142]}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, N639}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2769 ( .a ({new_AGEMA_signal_15146, new_AGEMA_signal_15138, new_AGEMA_signal_15130, new_AGEMA_signal_15122}), .b ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, n2670}), .clk ( clk ), .r ({Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148]}), .c ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, N723}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2855 ( .a ({new_AGEMA_signal_15162, new_AGEMA_signal_15158, new_AGEMA_signal_15154, new_AGEMA_signal_15150}), .b ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, n2831}), .clk ( clk ), .r ({Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154]}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, new_AGEMA_signal_3675, N789}) ) ;
    buf_clk new_AGEMA_reg_buffer_7142 ( .C ( clk ), .D ( new_AGEMA_signal_15169 ), .Q ( new_AGEMA_signal_15170 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7150 ( .C ( clk ), .D ( new_AGEMA_signal_15177 ), .Q ( new_AGEMA_signal_15178 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7158 ( .C ( clk ), .D ( new_AGEMA_signal_15185 ), .Q ( new_AGEMA_signal_15186 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7166 ( .C ( clk ), .D ( new_AGEMA_signal_15193 ), .Q ( new_AGEMA_signal_15194 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7172 ( .C ( clk ), .D ( new_AGEMA_signal_15199 ), .Q ( new_AGEMA_signal_15200 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7178 ( .C ( clk ), .D ( new_AGEMA_signal_15205 ), .Q ( new_AGEMA_signal_15206 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7184 ( .C ( clk ), .D ( new_AGEMA_signal_15211 ), .Q ( new_AGEMA_signal_15212 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7190 ( .C ( clk ), .D ( new_AGEMA_signal_15217 ), .Q ( new_AGEMA_signal_15218 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7192 ( .C ( clk ), .D ( new_AGEMA_signal_15219 ), .Q ( new_AGEMA_signal_15220 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7194 ( .C ( clk ), .D ( new_AGEMA_signal_15221 ), .Q ( new_AGEMA_signal_15222 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7196 ( .C ( clk ), .D ( new_AGEMA_signal_15223 ), .Q ( new_AGEMA_signal_15224 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7198 ( .C ( clk ), .D ( new_AGEMA_signal_15225 ), .Q ( new_AGEMA_signal_15226 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7218 ( .C ( clk ), .D ( new_AGEMA_signal_15245 ), .Q ( new_AGEMA_signal_15246 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7238 ( .C ( clk ), .D ( new_AGEMA_signal_15265 ), .Q ( new_AGEMA_signal_15266 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7258 ( .C ( clk ), .D ( new_AGEMA_signal_15285 ), .Q ( new_AGEMA_signal_15286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7278 ( .C ( clk ), .D ( new_AGEMA_signal_15305 ), .Q ( new_AGEMA_signal_15306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7284 ( .C ( clk ), .D ( new_AGEMA_signal_15311 ), .Q ( new_AGEMA_signal_15312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7292 ( .C ( clk ), .D ( new_AGEMA_signal_15319 ), .Q ( new_AGEMA_signal_15320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7300 ( .C ( clk ), .D ( new_AGEMA_signal_15327 ), .Q ( new_AGEMA_signal_15328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7308 ( .C ( clk ), .D ( new_AGEMA_signal_15335 ), .Q ( new_AGEMA_signal_15336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7320 ( .C ( clk ), .D ( new_AGEMA_signal_15347 ), .Q ( new_AGEMA_signal_15348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7332 ( .C ( clk ), .D ( new_AGEMA_signal_15359 ), .Q ( new_AGEMA_signal_15360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7344 ( .C ( clk ), .D ( new_AGEMA_signal_15371 ), .Q ( new_AGEMA_signal_15372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7356 ( .C ( clk ), .D ( new_AGEMA_signal_15383 ), .Q ( new_AGEMA_signal_15384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7368 ( .C ( clk ), .D ( new_AGEMA_signal_15395 ), .Q ( new_AGEMA_signal_15396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7382 ( .C ( clk ), .D ( new_AGEMA_signal_15409 ), .Q ( new_AGEMA_signal_15410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7396 ( .C ( clk ), .D ( new_AGEMA_signal_15423 ), .Q ( new_AGEMA_signal_15424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7410 ( .C ( clk ), .D ( new_AGEMA_signal_15437 ), .Q ( new_AGEMA_signal_15438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7422 ( .C ( clk ), .D ( new_AGEMA_signal_15449 ), .Q ( new_AGEMA_signal_15450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7436 ( .C ( clk ), .D ( new_AGEMA_signal_15463 ), .Q ( new_AGEMA_signal_15464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7450 ( .C ( clk ), .D ( new_AGEMA_signal_15477 ), .Q ( new_AGEMA_signal_15478 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7464 ( .C ( clk ), .D ( new_AGEMA_signal_15491 ), .Q ( new_AGEMA_signal_15492 ) ) ;

    /* cells in depth 27 */
    buf_clk new_AGEMA_reg_buffer_7285 ( .C ( clk ), .D ( new_AGEMA_signal_15312 ), .Q ( new_AGEMA_signal_15313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7293 ( .C ( clk ), .D ( new_AGEMA_signal_15320 ), .Q ( new_AGEMA_signal_15321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7301 ( .C ( clk ), .D ( new_AGEMA_signal_15328 ), .Q ( new_AGEMA_signal_15329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7309 ( .C ( clk ), .D ( new_AGEMA_signal_15336 ), .Q ( new_AGEMA_signal_15337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7321 ( .C ( clk ), .D ( new_AGEMA_signal_15348 ), .Q ( new_AGEMA_signal_15349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7333 ( .C ( clk ), .D ( new_AGEMA_signal_15360 ), .Q ( new_AGEMA_signal_15361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7345 ( .C ( clk ), .D ( new_AGEMA_signal_15372 ), .Q ( new_AGEMA_signal_15373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7357 ( .C ( clk ), .D ( new_AGEMA_signal_15384 ), .Q ( new_AGEMA_signal_15385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7369 ( .C ( clk ), .D ( new_AGEMA_signal_15396 ), .Q ( new_AGEMA_signal_15397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7383 ( .C ( clk ), .D ( new_AGEMA_signal_15410 ), .Q ( new_AGEMA_signal_15411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7397 ( .C ( clk ), .D ( new_AGEMA_signal_15424 ), .Q ( new_AGEMA_signal_15425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7411 ( .C ( clk ), .D ( new_AGEMA_signal_15438 ), .Q ( new_AGEMA_signal_15439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7423 ( .C ( clk ), .D ( new_AGEMA_signal_15450 ), .Q ( new_AGEMA_signal_15451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7437 ( .C ( clk ), .D ( new_AGEMA_signal_15464 ), .Q ( new_AGEMA_signal_15465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7451 ( .C ( clk ), .D ( new_AGEMA_signal_15478 ), .Q ( new_AGEMA_signal_15479 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7465 ( .C ( clk ), .D ( new_AGEMA_signal_15492 ), .Q ( new_AGEMA_signal_15493 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7535 ( .C ( clk ), .D ( N470 ), .Q ( new_AGEMA_signal_15563 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7543 ( .C ( clk ), .D ( new_AGEMA_signal_3687 ), .Q ( new_AGEMA_signal_15571 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7551 ( .C ( clk ), .D ( new_AGEMA_signal_3688 ), .Q ( new_AGEMA_signal_15579 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7559 ( .C ( clk ), .D ( new_AGEMA_signal_3689 ), .Q ( new_AGEMA_signal_15587 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7567 ( .C ( clk ), .D ( N639 ), .Q ( new_AGEMA_signal_15595 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7575 ( .C ( clk ), .D ( new_AGEMA_signal_3693 ), .Q ( new_AGEMA_signal_15603 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7583 ( .C ( clk ), .D ( new_AGEMA_signal_3694 ), .Q ( new_AGEMA_signal_15611 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7591 ( .C ( clk ), .D ( new_AGEMA_signal_3695 ), .Q ( new_AGEMA_signal_15619 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7599 ( .C ( clk ), .D ( N723 ), .Q ( new_AGEMA_signal_15627 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7607 ( .C ( clk ), .D ( new_AGEMA_signal_3696 ), .Q ( new_AGEMA_signal_15635 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7615 ( .C ( clk ), .D ( new_AGEMA_signal_3697 ), .Q ( new_AGEMA_signal_15643 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7623 ( .C ( clk ), .D ( new_AGEMA_signal_3698 ), .Q ( new_AGEMA_signal_15651 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7631 ( .C ( clk ), .D ( N789 ), .Q ( new_AGEMA_signal_15659 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7639 ( .C ( clk ), .D ( new_AGEMA_signal_3675 ), .Q ( new_AGEMA_signal_15667 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7647 ( .C ( clk ), .D ( new_AGEMA_signal_3676 ), .Q ( new_AGEMA_signal_15675 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7655 ( .C ( clk ), .D ( new_AGEMA_signal_3677 ), .Q ( new_AGEMA_signal_15683 ) ) ;

    /* cells in depth 28 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2156 ( .a ({new_AGEMA_signal_15194, new_AGEMA_signal_15186, new_AGEMA_signal_15178, new_AGEMA_signal_15170}), .b ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, n2018}), .clk ( clk ), .r ({Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160]}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, N169}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2270 ( .a ({new_AGEMA_signal_15218, new_AGEMA_signal_15212, new_AGEMA_signal_15206, new_AGEMA_signal_15200}), .b ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, new_AGEMA_signal_3681, n2112}), .clk ( clk ), .r ({Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166]}), .c ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, N277}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2376 ( .a ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, n2210}), .b ({new_AGEMA_signal_15226, new_AGEMA_signal_15224, new_AGEMA_signal_15222, new_AGEMA_signal_15220}), .clk ( clk ), .r ({Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172]}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, n2211}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2540 ( .a ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, n2378}), .b ({new_AGEMA_signal_15306, new_AGEMA_signal_15286, new_AGEMA_signal_15266, new_AGEMA_signal_15246}), .clk ( clk ), .r ({Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178]}), .c ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, n2379}) ) ;
    buf_clk new_AGEMA_reg_buffer_7286 ( .C ( clk ), .D ( new_AGEMA_signal_15313 ), .Q ( new_AGEMA_signal_15314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7294 ( .C ( clk ), .D ( new_AGEMA_signal_15321 ), .Q ( new_AGEMA_signal_15322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7302 ( .C ( clk ), .D ( new_AGEMA_signal_15329 ), .Q ( new_AGEMA_signal_15330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7310 ( .C ( clk ), .D ( new_AGEMA_signal_15337 ), .Q ( new_AGEMA_signal_15338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7322 ( .C ( clk ), .D ( new_AGEMA_signal_15349 ), .Q ( new_AGEMA_signal_15350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7334 ( .C ( clk ), .D ( new_AGEMA_signal_15361 ), .Q ( new_AGEMA_signal_15362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7346 ( .C ( clk ), .D ( new_AGEMA_signal_15373 ), .Q ( new_AGEMA_signal_15374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7358 ( .C ( clk ), .D ( new_AGEMA_signal_15385 ), .Q ( new_AGEMA_signal_15386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7370 ( .C ( clk ), .D ( new_AGEMA_signal_15397 ), .Q ( new_AGEMA_signal_15398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7384 ( .C ( clk ), .D ( new_AGEMA_signal_15411 ), .Q ( new_AGEMA_signal_15412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7398 ( .C ( clk ), .D ( new_AGEMA_signal_15425 ), .Q ( new_AGEMA_signal_15426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7412 ( .C ( clk ), .D ( new_AGEMA_signal_15439 ), .Q ( new_AGEMA_signal_15440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7424 ( .C ( clk ), .D ( new_AGEMA_signal_15451 ), .Q ( new_AGEMA_signal_15452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7438 ( .C ( clk ), .D ( new_AGEMA_signal_15465 ), .Q ( new_AGEMA_signal_15466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7452 ( .C ( clk ), .D ( new_AGEMA_signal_15479 ), .Q ( new_AGEMA_signal_15480 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7466 ( .C ( clk ), .D ( new_AGEMA_signal_15493 ), .Q ( new_AGEMA_signal_15494 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7536 ( .C ( clk ), .D ( new_AGEMA_signal_15563 ), .Q ( new_AGEMA_signal_15564 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7544 ( .C ( clk ), .D ( new_AGEMA_signal_15571 ), .Q ( new_AGEMA_signal_15572 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7552 ( .C ( clk ), .D ( new_AGEMA_signal_15579 ), .Q ( new_AGEMA_signal_15580 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7560 ( .C ( clk ), .D ( new_AGEMA_signal_15587 ), .Q ( new_AGEMA_signal_15588 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7568 ( .C ( clk ), .D ( new_AGEMA_signal_15595 ), .Q ( new_AGEMA_signal_15596 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7576 ( .C ( clk ), .D ( new_AGEMA_signal_15603 ), .Q ( new_AGEMA_signal_15604 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7584 ( .C ( clk ), .D ( new_AGEMA_signal_15611 ), .Q ( new_AGEMA_signal_15612 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7592 ( .C ( clk ), .D ( new_AGEMA_signal_15619 ), .Q ( new_AGEMA_signal_15620 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7600 ( .C ( clk ), .D ( new_AGEMA_signal_15627 ), .Q ( new_AGEMA_signal_15628 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7608 ( .C ( clk ), .D ( new_AGEMA_signal_15635 ), .Q ( new_AGEMA_signal_15636 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7616 ( .C ( clk ), .D ( new_AGEMA_signal_15643 ), .Q ( new_AGEMA_signal_15644 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7624 ( .C ( clk ), .D ( new_AGEMA_signal_15651 ), .Q ( new_AGEMA_signal_15652 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7632 ( .C ( clk ), .D ( new_AGEMA_signal_15659 ), .Q ( new_AGEMA_signal_15660 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7640 ( .C ( clk ), .D ( new_AGEMA_signal_15667 ), .Q ( new_AGEMA_signal_15668 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7648 ( .C ( clk ), .D ( new_AGEMA_signal_15675 ), .Q ( new_AGEMA_signal_15676 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7656 ( .C ( clk ), .D ( new_AGEMA_signal_15683 ), .Q ( new_AGEMA_signal_15684 ) ) ;

    /* cells in depth 29 */
    buf_clk new_AGEMA_reg_buffer_7371 ( .C ( clk ), .D ( new_AGEMA_signal_15398 ), .Q ( new_AGEMA_signal_15399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7385 ( .C ( clk ), .D ( new_AGEMA_signal_15412 ), .Q ( new_AGEMA_signal_15413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7399 ( .C ( clk ), .D ( new_AGEMA_signal_15426 ), .Q ( new_AGEMA_signal_15427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7413 ( .C ( clk ), .D ( new_AGEMA_signal_15440 ), .Q ( new_AGEMA_signal_15441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7425 ( .C ( clk ), .D ( new_AGEMA_signal_15452 ), .Q ( new_AGEMA_signal_15453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7439 ( .C ( clk ), .D ( new_AGEMA_signal_15466 ), .Q ( new_AGEMA_signal_15467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7453 ( .C ( clk ), .D ( new_AGEMA_signal_15480 ), .Q ( new_AGEMA_signal_15481 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7467 ( .C ( clk ), .D ( new_AGEMA_signal_15494 ), .Q ( new_AGEMA_signal_15495 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7471 ( .C ( clk ), .D ( N169 ), .Q ( new_AGEMA_signal_15499 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7477 ( .C ( clk ), .D ( new_AGEMA_signal_3699 ), .Q ( new_AGEMA_signal_15505 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7483 ( .C ( clk ), .D ( new_AGEMA_signal_3700 ), .Q ( new_AGEMA_signal_15511 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7489 ( .C ( clk ), .D ( new_AGEMA_signal_3701 ), .Q ( new_AGEMA_signal_15517 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7495 ( .C ( clk ), .D ( N277 ), .Q ( new_AGEMA_signal_15523 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7501 ( .C ( clk ), .D ( new_AGEMA_signal_3702 ), .Q ( new_AGEMA_signal_15529 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7507 ( .C ( clk ), .D ( new_AGEMA_signal_3703 ), .Q ( new_AGEMA_signal_15535 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7513 ( .C ( clk ), .D ( new_AGEMA_signal_3704 ), .Q ( new_AGEMA_signal_15541 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7537 ( .C ( clk ), .D ( new_AGEMA_signal_15564 ), .Q ( new_AGEMA_signal_15565 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7545 ( .C ( clk ), .D ( new_AGEMA_signal_15572 ), .Q ( new_AGEMA_signal_15573 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7553 ( .C ( clk ), .D ( new_AGEMA_signal_15580 ), .Q ( new_AGEMA_signal_15581 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7561 ( .C ( clk ), .D ( new_AGEMA_signal_15588 ), .Q ( new_AGEMA_signal_15589 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7569 ( .C ( clk ), .D ( new_AGEMA_signal_15596 ), .Q ( new_AGEMA_signal_15597 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7577 ( .C ( clk ), .D ( new_AGEMA_signal_15604 ), .Q ( new_AGEMA_signal_15605 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7585 ( .C ( clk ), .D ( new_AGEMA_signal_15612 ), .Q ( new_AGEMA_signal_15613 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7593 ( .C ( clk ), .D ( new_AGEMA_signal_15620 ), .Q ( new_AGEMA_signal_15621 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7601 ( .C ( clk ), .D ( new_AGEMA_signal_15628 ), .Q ( new_AGEMA_signal_15629 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7609 ( .C ( clk ), .D ( new_AGEMA_signal_15636 ), .Q ( new_AGEMA_signal_15637 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7617 ( .C ( clk ), .D ( new_AGEMA_signal_15644 ), .Q ( new_AGEMA_signal_15645 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7625 ( .C ( clk ), .D ( new_AGEMA_signal_15652 ), .Q ( new_AGEMA_signal_15653 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7633 ( .C ( clk ), .D ( new_AGEMA_signal_15660 ), .Q ( new_AGEMA_signal_15661 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7641 ( .C ( clk ), .D ( new_AGEMA_signal_15668 ), .Q ( new_AGEMA_signal_15669 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7649 ( .C ( clk ), .D ( new_AGEMA_signal_15676 ), .Q ( new_AGEMA_signal_15677 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7657 ( .C ( clk ), .D ( new_AGEMA_signal_15684 ), .Q ( new_AGEMA_signal_15685 ) ) ;

    /* cells in depth 30 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2377 ( .a ({new_AGEMA_signal_15338, new_AGEMA_signal_15330, new_AGEMA_signal_15322, new_AGEMA_signal_15314}), .b ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, n2211}), .clk ( clk ), .r ({Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184]}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, N379}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2541 ( .a ({new_AGEMA_signal_15386, new_AGEMA_signal_15374, new_AGEMA_signal_15362, new_AGEMA_signal_15350}), .b ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, n2379}), .clk ( clk ), .r ({Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190]}), .c ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2381}) ) ;
    buf_clk new_AGEMA_reg_buffer_7372 ( .C ( clk ), .D ( new_AGEMA_signal_15399 ), .Q ( new_AGEMA_signal_15400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7386 ( .C ( clk ), .D ( new_AGEMA_signal_15413 ), .Q ( new_AGEMA_signal_15414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7400 ( .C ( clk ), .D ( new_AGEMA_signal_15427 ), .Q ( new_AGEMA_signal_15428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7414 ( .C ( clk ), .D ( new_AGEMA_signal_15441 ), .Q ( new_AGEMA_signal_15442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7426 ( .C ( clk ), .D ( new_AGEMA_signal_15453 ), .Q ( new_AGEMA_signal_15454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7440 ( .C ( clk ), .D ( new_AGEMA_signal_15467 ), .Q ( new_AGEMA_signal_15468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7454 ( .C ( clk ), .D ( new_AGEMA_signal_15481 ), .Q ( new_AGEMA_signal_15482 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7468 ( .C ( clk ), .D ( new_AGEMA_signal_15495 ), .Q ( new_AGEMA_signal_15496 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7472 ( .C ( clk ), .D ( new_AGEMA_signal_15499 ), .Q ( new_AGEMA_signal_15500 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7478 ( .C ( clk ), .D ( new_AGEMA_signal_15505 ), .Q ( new_AGEMA_signal_15506 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7484 ( .C ( clk ), .D ( new_AGEMA_signal_15511 ), .Q ( new_AGEMA_signal_15512 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7490 ( .C ( clk ), .D ( new_AGEMA_signal_15517 ), .Q ( new_AGEMA_signal_15518 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7496 ( .C ( clk ), .D ( new_AGEMA_signal_15523 ), .Q ( new_AGEMA_signal_15524 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7502 ( .C ( clk ), .D ( new_AGEMA_signal_15529 ), .Q ( new_AGEMA_signal_15530 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7508 ( .C ( clk ), .D ( new_AGEMA_signal_15535 ), .Q ( new_AGEMA_signal_15536 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7514 ( .C ( clk ), .D ( new_AGEMA_signal_15541 ), .Q ( new_AGEMA_signal_15542 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7538 ( .C ( clk ), .D ( new_AGEMA_signal_15565 ), .Q ( new_AGEMA_signal_15566 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7546 ( .C ( clk ), .D ( new_AGEMA_signal_15573 ), .Q ( new_AGEMA_signal_15574 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7554 ( .C ( clk ), .D ( new_AGEMA_signal_15581 ), .Q ( new_AGEMA_signal_15582 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7562 ( .C ( clk ), .D ( new_AGEMA_signal_15589 ), .Q ( new_AGEMA_signal_15590 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7570 ( .C ( clk ), .D ( new_AGEMA_signal_15597 ), .Q ( new_AGEMA_signal_15598 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7578 ( .C ( clk ), .D ( new_AGEMA_signal_15605 ), .Q ( new_AGEMA_signal_15606 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7586 ( .C ( clk ), .D ( new_AGEMA_signal_15613 ), .Q ( new_AGEMA_signal_15614 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7594 ( .C ( clk ), .D ( new_AGEMA_signal_15621 ), .Q ( new_AGEMA_signal_15622 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7602 ( .C ( clk ), .D ( new_AGEMA_signal_15629 ), .Q ( new_AGEMA_signal_15630 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7610 ( .C ( clk ), .D ( new_AGEMA_signal_15637 ), .Q ( new_AGEMA_signal_15638 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7618 ( .C ( clk ), .D ( new_AGEMA_signal_15645 ), .Q ( new_AGEMA_signal_15646 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7626 ( .C ( clk ), .D ( new_AGEMA_signal_15653 ), .Q ( new_AGEMA_signal_15654 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7634 ( .C ( clk ), .D ( new_AGEMA_signal_15661 ), .Q ( new_AGEMA_signal_15662 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7642 ( .C ( clk ), .D ( new_AGEMA_signal_15669 ), .Q ( new_AGEMA_signal_15670 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7650 ( .C ( clk ), .D ( new_AGEMA_signal_15677 ), .Q ( new_AGEMA_signal_15678 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7658 ( .C ( clk ), .D ( new_AGEMA_signal_15685 ), .Q ( new_AGEMA_signal_15686 ) ) ;

    /* cells in depth 31 */
    buf_clk new_AGEMA_reg_buffer_7427 ( .C ( clk ), .D ( new_AGEMA_signal_15454 ), .Q ( new_AGEMA_signal_15455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7441 ( .C ( clk ), .D ( new_AGEMA_signal_15468 ), .Q ( new_AGEMA_signal_15469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7455 ( .C ( clk ), .D ( new_AGEMA_signal_15482 ), .Q ( new_AGEMA_signal_15483 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7469 ( .C ( clk ), .D ( new_AGEMA_signal_15496 ), .Q ( new_AGEMA_signal_15497 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7473 ( .C ( clk ), .D ( new_AGEMA_signal_15500 ), .Q ( new_AGEMA_signal_15501 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7479 ( .C ( clk ), .D ( new_AGEMA_signal_15506 ), .Q ( new_AGEMA_signal_15507 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7485 ( .C ( clk ), .D ( new_AGEMA_signal_15512 ), .Q ( new_AGEMA_signal_15513 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7491 ( .C ( clk ), .D ( new_AGEMA_signal_15518 ), .Q ( new_AGEMA_signal_15519 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7497 ( .C ( clk ), .D ( new_AGEMA_signal_15524 ), .Q ( new_AGEMA_signal_15525 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7503 ( .C ( clk ), .D ( new_AGEMA_signal_15530 ), .Q ( new_AGEMA_signal_15531 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7509 ( .C ( clk ), .D ( new_AGEMA_signal_15536 ), .Q ( new_AGEMA_signal_15537 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7515 ( .C ( clk ), .D ( new_AGEMA_signal_15542 ), .Q ( new_AGEMA_signal_15543 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7519 ( .C ( clk ), .D ( N379 ), .Q ( new_AGEMA_signal_15547 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7523 ( .C ( clk ), .D ( new_AGEMA_signal_3711 ), .Q ( new_AGEMA_signal_15551 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7527 ( .C ( clk ), .D ( new_AGEMA_signal_3712 ), .Q ( new_AGEMA_signal_15555 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7531 ( .C ( clk ), .D ( new_AGEMA_signal_3713 ), .Q ( new_AGEMA_signal_15559 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7539 ( .C ( clk ), .D ( new_AGEMA_signal_15566 ), .Q ( new_AGEMA_signal_15567 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7547 ( .C ( clk ), .D ( new_AGEMA_signal_15574 ), .Q ( new_AGEMA_signal_15575 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7555 ( .C ( clk ), .D ( new_AGEMA_signal_15582 ), .Q ( new_AGEMA_signal_15583 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7563 ( .C ( clk ), .D ( new_AGEMA_signal_15590 ), .Q ( new_AGEMA_signal_15591 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7571 ( .C ( clk ), .D ( new_AGEMA_signal_15598 ), .Q ( new_AGEMA_signal_15599 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7579 ( .C ( clk ), .D ( new_AGEMA_signal_15606 ), .Q ( new_AGEMA_signal_15607 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7587 ( .C ( clk ), .D ( new_AGEMA_signal_15614 ), .Q ( new_AGEMA_signal_15615 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7595 ( .C ( clk ), .D ( new_AGEMA_signal_15622 ), .Q ( new_AGEMA_signal_15623 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7603 ( .C ( clk ), .D ( new_AGEMA_signal_15630 ), .Q ( new_AGEMA_signal_15631 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7611 ( .C ( clk ), .D ( new_AGEMA_signal_15638 ), .Q ( new_AGEMA_signal_15639 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7619 ( .C ( clk ), .D ( new_AGEMA_signal_15646 ), .Q ( new_AGEMA_signal_15647 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7627 ( .C ( clk ), .D ( new_AGEMA_signal_15654 ), .Q ( new_AGEMA_signal_15655 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7635 ( .C ( clk ), .D ( new_AGEMA_signal_15662 ), .Q ( new_AGEMA_signal_15663 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7643 ( .C ( clk ), .D ( new_AGEMA_signal_15670 ), .Q ( new_AGEMA_signal_15671 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7651 ( .C ( clk ), .D ( new_AGEMA_signal_15678 ), .Q ( new_AGEMA_signal_15679 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7659 ( .C ( clk ), .D ( new_AGEMA_signal_15686 ), .Q ( new_AGEMA_signal_15687 ) ) ;

    /* cells in depth 32 */
    nor_HPC2 #(.security_order(3), .pipeline(1)) U2542 ( .a ({new_AGEMA_signal_15442, new_AGEMA_signal_15428, new_AGEMA_signal_15414, new_AGEMA_signal_15400}), .b ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, n2381}), .clk ( clk ), .r ({Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196]}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, n2427}) ) ;
    buf_clk new_AGEMA_reg_buffer_7428 ( .C ( clk ), .D ( new_AGEMA_signal_15455 ), .Q ( new_AGEMA_signal_15456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7442 ( .C ( clk ), .D ( new_AGEMA_signal_15469 ), .Q ( new_AGEMA_signal_15470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7456 ( .C ( clk ), .D ( new_AGEMA_signal_15483 ), .Q ( new_AGEMA_signal_15484 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7470 ( .C ( clk ), .D ( new_AGEMA_signal_15497 ), .Q ( new_AGEMA_signal_15498 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7474 ( .C ( clk ), .D ( new_AGEMA_signal_15501 ), .Q ( new_AGEMA_signal_15502 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7480 ( .C ( clk ), .D ( new_AGEMA_signal_15507 ), .Q ( new_AGEMA_signal_15508 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7486 ( .C ( clk ), .D ( new_AGEMA_signal_15513 ), .Q ( new_AGEMA_signal_15514 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7492 ( .C ( clk ), .D ( new_AGEMA_signal_15519 ), .Q ( new_AGEMA_signal_15520 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7498 ( .C ( clk ), .D ( new_AGEMA_signal_15525 ), .Q ( new_AGEMA_signal_15526 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7504 ( .C ( clk ), .D ( new_AGEMA_signal_15531 ), .Q ( new_AGEMA_signal_15532 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7510 ( .C ( clk ), .D ( new_AGEMA_signal_15537 ), .Q ( new_AGEMA_signal_15538 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7516 ( .C ( clk ), .D ( new_AGEMA_signal_15543 ), .Q ( new_AGEMA_signal_15544 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7520 ( .C ( clk ), .D ( new_AGEMA_signal_15547 ), .Q ( new_AGEMA_signal_15548 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7524 ( .C ( clk ), .D ( new_AGEMA_signal_15551 ), .Q ( new_AGEMA_signal_15552 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7528 ( .C ( clk ), .D ( new_AGEMA_signal_15555 ), .Q ( new_AGEMA_signal_15556 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7532 ( .C ( clk ), .D ( new_AGEMA_signal_15559 ), .Q ( new_AGEMA_signal_15560 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7540 ( .C ( clk ), .D ( new_AGEMA_signal_15567 ), .Q ( new_AGEMA_signal_15568 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7548 ( .C ( clk ), .D ( new_AGEMA_signal_15575 ), .Q ( new_AGEMA_signal_15576 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7556 ( .C ( clk ), .D ( new_AGEMA_signal_15583 ), .Q ( new_AGEMA_signal_15584 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7564 ( .C ( clk ), .D ( new_AGEMA_signal_15591 ), .Q ( new_AGEMA_signal_15592 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7572 ( .C ( clk ), .D ( new_AGEMA_signal_15599 ), .Q ( new_AGEMA_signal_15600 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7580 ( .C ( clk ), .D ( new_AGEMA_signal_15607 ), .Q ( new_AGEMA_signal_15608 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7588 ( .C ( clk ), .D ( new_AGEMA_signal_15615 ), .Q ( new_AGEMA_signal_15616 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7596 ( .C ( clk ), .D ( new_AGEMA_signal_15623 ), .Q ( new_AGEMA_signal_15624 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7604 ( .C ( clk ), .D ( new_AGEMA_signal_15631 ), .Q ( new_AGEMA_signal_15632 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7612 ( .C ( clk ), .D ( new_AGEMA_signal_15639 ), .Q ( new_AGEMA_signal_15640 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7620 ( .C ( clk ), .D ( new_AGEMA_signal_15647 ), .Q ( new_AGEMA_signal_15648 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7628 ( .C ( clk ), .D ( new_AGEMA_signal_15655 ), .Q ( new_AGEMA_signal_15656 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7636 ( .C ( clk ), .D ( new_AGEMA_signal_15663 ), .Q ( new_AGEMA_signal_15664 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7644 ( .C ( clk ), .D ( new_AGEMA_signal_15671 ), .Q ( new_AGEMA_signal_15672 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7652 ( .C ( clk ), .D ( new_AGEMA_signal_15679 ), .Q ( new_AGEMA_signal_15680 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7660 ( .C ( clk ), .D ( new_AGEMA_signal_15687 ), .Q ( new_AGEMA_signal_15688 ) ) ;

    /* cells in depth 33 */
    buf_clk new_AGEMA_reg_buffer_7475 ( .C ( clk ), .D ( new_AGEMA_signal_15502 ), .Q ( new_AGEMA_signal_15503 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7481 ( .C ( clk ), .D ( new_AGEMA_signal_15508 ), .Q ( new_AGEMA_signal_15509 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7487 ( .C ( clk ), .D ( new_AGEMA_signal_15514 ), .Q ( new_AGEMA_signal_15515 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7493 ( .C ( clk ), .D ( new_AGEMA_signal_15520 ), .Q ( new_AGEMA_signal_15521 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7499 ( .C ( clk ), .D ( new_AGEMA_signal_15526 ), .Q ( new_AGEMA_signal_15527 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7505 ( .C ( clk ), .D ( new_AGEMA_signal_15532 ), .Q ( new_AGEMA_signal_15533 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7511 ( .C ( clk ), .D ( new_AGEMA_signal_15538 ), .Q ( new_AGEMA_signal_15539 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7517 ( .C ( clk ), .D ( new_AGEMA_signal_15544 ), .Q ( new_AGEMA_signal_15545 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7521 ( .C ( clk ), .D ( new_AGEMA_signal_15548 ), .Q ( new_AGEMA_signal_15549 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7525 ( .C ( clk ), .D ( new_AGEMA_signal_15552 ), .Q ( new_AGEMA_signal_15553 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7529 ( .C ( clk ), .D ( new_AGEMA_signal_15556 ), .Q ( new_AGEMA_signal_15557 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7533 ( .C ( clk ), .D ( new_AGEMA_signal_15560 ), .Q ( new_AGEMA_signal_15561 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7541 ( .C ( clk ), .D ( new_AGEMA_signal_15568 ), .Q ( new_AGEMA_signal_15569 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7549 ( .C ( clk ), .D ( new_AGEMA_signal_15576 ), .Q ( new_AGEMA_signal_15577 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7557 ( .C ( clk ), .D ( new_AGEMA_signal_15584 ), .Q ( new_AGEMA_signal_15585 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7565 ( .C ( clk ), .D ( new_AGEMA_signal_15592 ), .Q ( new_AGEMA_signal_15593 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7573 ( .C ( clk ), .D ( new_AGEMA_signal_15600 ), .Q ( new_AGEMA_signal_15601 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7581 ( .C ( clk ), .D ( new_AGEMA_signal_15608 ), .Q ( new_AGEMA_signal_15609 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7589 ( .C ( clk ), .D ( new_AGEMA_signal_15616 ), .Q ( new_AGEMA_signal_15617 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7597 ( .C ( clk ), .D ( new_AGEMA_signal_15624 ), .Q ( new_AGEMA_signal_15625 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7605 ( .C ( clk ), .D ( new_AGEMA_signal_15632 ), .Q ( new_AGEMA_signal_15633 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7613 ( .C ( clk ), .D ( new_AGEMA_signal_15640 ), .Q ( new_AGEMA_signal_15641 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7621 ( .C ( clk ), .D ( new_AGEMA_signal_15648 ), .Q ( new_AGEMA_signal_15649 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7629 ( .C ( clk ), .D ( new_AGEMA_signal_15656 ), .Q ( new_AGEMA_signal_15657 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7637 ( .C ( clk ), .D ( new_AGEMA_signal_15664 ), .Q ( new_AGEMA_signal_15665 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7645 ( .C ( clk ), .D ( new_AGEMA_signal_15672 ), .Q ( new_AGEMA_signal_15673 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7653 ( .C ( clk ), .D ( new_AGEMA_signal_15680 ), .Q ( new_AGEMA_signal_15681 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7661 ( .C ( clk ), .D ( new_AGEMA_signal_15688 ), .Q ( new_AGEMA_signal_15689 ) ) ;

    /* cells in depth 34 */
    nand_HPC2 #(.security_order(3), .pipeline(1)) U2584 ( .a ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, n2427}), .b ({new_AGEMA_signal_15498, new_AGEMA_signal_15484, new_AGEMA_signal_15470, new_AGEMA_signal_15456}), .clk ( clk ), .r ({Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202]}), .c ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, N563}) ) ;
    buf_clk new_AGEMA_reg_buffer_7476 ( .C ( clk ), .D ( new_AGEMA_signal_15503 ), .Q ( new_AGEMA_signal_15504 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7482 ( .C ( clk ), .D ( new_AGEMA_signal_15509 ), .Q ( new_AGEMA_signal_15510 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7488 ( .C ( clk ), .D ( new_AGEMA_signal_15515 ), .Q ( new_AGEMA_signal_15516 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7494 ( .C ( clk ), .D ( new_AGEMA_signal_15521 ), .Q ( new_AGEMA_signal_15522 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7500 ( .C ( clk ), .D ( new_AGEMA_signal_15527 ), .Q ( new_AGEMA_signal_15528 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7506 ( .C ( clk ), .D ( new_AGEMA_signal_15533 ), .Q ( new_AGEMA_signal_15534 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7512 ( .C ( clk ), .D ( new_AGEMA_signal_15539 ), .Q ( new_AGEMA_signal_15540 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7518 ( .C ( clk ), .D ( new_AGEMA_signal_15545 ), .Q ( new_AGEMA_signal_15546 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7522 ( .C ( clk ), .D ( new_AGEMA_signal_15549 ), .Q ( new_AGEMA_signal_15550 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7526 ( .C ( clk ), .D ( new_AGEMA_signal_15553 ), .Q ( new_AGEMA_signal_15554 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7530 ( .C ( clk ), .D ( new_AGEMA_signal_15557 ), .Q ( new_AGEMA_signal_15558 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7534 ( .C ( clk ), .D ( new_AGEMA_signal_15561 ), .Q ( new_AGEMA_signal_15562 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7542 ( .C ( clk ), .D ( new_AGEMA_signal_15569 ), .Q ( new_AGEMA_signal_15570 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7550 ( .C ( clk ), .D ( new_AGEMA_signal_15577 ), .Q ( new_AGEMA_signal_15578 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7558 ( .C ( clk ), .D ( new_AGEMA_signal_15585 ), .Q ( new_AGEMA_signal_15586 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7566 ( .C ( clk ), .D ( new_AGEMA_signal_15593 ), .Q ( new_AGEMA_signal_15594 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7574 ( .C ( clk ), .D ( new_AGEMA_signal_15601 ), .Q ( new_AGEMA_signal_15602 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7582 ( .C ( clk ), .D ( new_AGEMA_signal_15609 ), .Q ( new_AGEMA_signal_15610 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7590 ( .C ( clk ), .D ( new_AGEMA_signal_15617 ), .Q ( new_AGEMA_signal_15618 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7598 ( .C ( clk ), .D ( new_AGEMA_signal_15625 ), .Q ( new_AGEMA_signal_15626 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7606 ( .C ( clk ), .D ( new_AGEMA_signal_15633 ), .Q ( new_AGEMA_signal_15634 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7614 ( .C ( clk ), .D ( new_AGEMA_signal_15641 ), .Q ( new_AGEMA_signal_15642 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7622 ( .C ( clk ), .D ( new_AGEMA_signal_15649 ), .Q ( new_AGEMA_signal_15650 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7630 ( .C ( clk ), .D ( new_AGEMA_signal_15657 ), .Q ( new_AGEMA_signal_15658 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7638 ( .C ( clk ), .D ( new_AGEMA_signal_15665 ), .Q ( new_AGEMA_signal_15666 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7646 ( .C ( clk ), .D ( new_AGEMA_signal_15673 ), .Q ( new_AGEMA_signal_15674 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7654 ( .C ( clk ), .D ( new_AGEMA_signal_15681 ), .Q ( new_AGEMA_signal_15682 ) ) ;
    buf_clk new_AGEMA_reg_buffer_7662 ( .C ( clk ), .D ( new_AGEMA_signal_15689 ), .Q ( new_AGEMA_signal_15690 ) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_7_ ( .clk ( clk ), .D ({new_AGEMA_signal_15522, new_AGEMA_signal_15516, new_AGEMA_signal_15510, new_AGEMA_signal_15504}), .Q ({SO_s3[7], SO_s2[7], SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_6_ ( .clk ( clk ), .D ({new_AGEMA_signal_15546, new_AGEMA_signal_15540, new_AGEMA_signal_15534, new_AGEMA_signal_15528}), .Q ({SO_s3[6], SO_s2[6], SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_5_ ( .clk ( clk ), .D ({new_AGEMA_signal_15562, new_AGEMA_signal_15558, new_AGEMA_signal_15554, new_AGEMA_signal_15550}), .Q ({SO_s3[5], SO_s2[5], SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_4_ ( .clk ( clk ), .D ({new_AGEMA_signal_15594, new_AGEMA_signal_15586, new_AGEMA_signal_15578, new_AGEMA_signal_15570}), .Q ({SO_s3[4], SO_s2[4], SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, N563}), .Q ({SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_15626, new_AGEMA_signal_15618, new_AGEMA_signal_15610, new_AGEMA_signal_15602}), .Q ({SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_15658, new_AGEMA_signal_15650, new_AGEMA_signal_15642, new_AGEMA_signal_15634}), .Q ({SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_15690, new_AGEMA_signal_15682, new_AGEMA_signal_15674, new_AGEMA_signal_15666}), .Q ({SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
