/* modified netlist. Source: module AES in file AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_GHPC_ClockGating_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [135:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output Synch ;
    wire AKSRnotDone ;
    wire LastRoundorDone ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire n55 ;
    wire n56 ;
    wire n57 ;
    wire n58 ;
    wire n59 ;
    wire n60 ;
    wire n61 ;
    wire n62 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire MuxSboxIn_n7 ;
    wire MuxSboxIn_n6 ;
    wire MuxSboxIn_n5 ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire MixColumnsIns_n64 ;
    wire MixColumnsIns_n63 ;
    wire MixColumnsIns_n62 ;
    wire MixColumnsIns_n61 ;
    wire MixColumnsIns_n60 ;
    wire MixColumnsIns_n59 ;
    wire MixColumnsIns_n58 ;
    wire MixColumnsIns_n57 ;
    wire MixColumnsIns_n56 ;
    wire MixColumnsIns_n55 ;
    wire MixColumnsIns_n54 ;
    wire MixColumnsIns_n53 ;
    wire MixColumnsIns_n52 ;
    wire MixColumnsIns_n51 ;
    wire MixColumnsIns_n50 ;
    wire MixColumnsIns_n49 ;
    wire MixColumnsIns_n48 ;
    wire MixColumnsIns_n47 ;
    wire MixColumnsIns_n46 ;
    wire MixColumnsIns_n45 ;
    wire MixColumnsIns_n44 ;
    wire MixColumnsIns_n43 ;
    wire MixColumnsIns_n42 ;
    wire MixColumnsIns_n41 ;
    wire MixColumnsIns_n40 ;
    wire MixColumnsIns_n39 ;
    wire MixColumnsIns_n38 ;
    wire MixColumnsIns_n37 ;
    wire MixColumnsIns_n36 ;
    wire MixColumnsIns_n35 ;
    wire MixColumnsIns_n34 ;
    wire MixColumnsIns_n33 ;
    wire MixColumnsIns_n32 ;
    wire MixColumnsIns_n31 ;
    wire MixColumnsIns_n30 ;
    wire MixColumnsIns_n29 ;
    wire MixColumnsIns_n28 ;
    wire MixColumnsIns_n27 ;
    wire MixColumnsIns_n26 ;
    wire MixColumnsIns_n25 ;
    wire MixColumnsIns_n24 ;
    wire MixColumnsIns_n23 ;
    wire MixColumnsIns_n22 ;
    wire MixColumnsIns_n21 ;
    wire MixColumnsIns_n20 ;
    wire MixColumnsIns_n19 ;
    wire MixColumnsIns_n18 ;
    wire MixColumnsIns_n17 ;
    wire MixColumnsIns_n16 ;
    wire MixColumnsIns_n15 ;
    wire MixColumnsIns_n14 ;
    wire MixColumnsIns_n13 ;
    wire MixColumnsIns_n12 ;
    wire MixColumnsIns_n11 ;
    wire MixColumnsIns_n10 ;
    wire MixColumnsIns_n9 ;
    wire MixColumnsIns_n8 ;
    wire MixColumnsIns_n7 ;
    wire MixColumnsIns_n6 ;
    wire MixColumnsIns_n5 ;
    wire MixColumnsIns_n4 ;
    wire MixColumnsIns_n3 ;
    wire MixColumnsIns_n2 ;
    wire MixColumnsIns_n1 ;
    wire MuxMCOut_n6 ;
    wire MuxMCOut_n5 ;
    wire MuxMCOut_n4 ;
    wire MuxRound_n19 ;
    wire MuxRound_n18 ;
    wire MuxRound_n17 ;
    wire MuxRound_n16 ;
    wire MuxRound_n15 ;
    wire MuxRound_n14 ;
    wire MuxRound_n13 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire MuxKeyExpansion_n21 ;
    wire MuxKeyExpansion_n20 ;
    wire MuxKeyExpansion_n19 ;
    wire MuxKeyExpansion_n18 ;
    wire MuxKeyExpansion_n17 ;
    wire MuxKeyExpansion_n16 ;
    wire MuxKeyExpansion_n15 ;
    wire MuxKeyExpansion_n14 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n42 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n44 ;
    wire RoundCounterIns_n45 ;
    wire InRoundCounterIns_n12 ;
    wire InRoundCounterIns_n11 ;
    wire InRoundCounterIns_n10 ;
    wire InRoundCounterIns_n9 ;
    wire InRoundCounterIns_n8 ;
    wire InRoundCounterIns_n7 ;
    wire InRoundCounterIns_n5 ;
    wire InRoundCounterIns_n4 ;
    wire InRoundCounterIns_n3 ;
    wire InRoundCounterIns_n2 ;
    wire InRoundCounterIns_n1 ;
    wire InRoundCounterIns_n6 ;
    wire InRoundCounterIns_n39 ;
    wire InRoundCounterIns_n40 ;
    wire InRoundCounterIns_n41 ;
    wire [127:0] RoundOutput ;
    wire [127:0] ShiftRowsOutput ;
    wire [31:0] KSSubBytesInput ;
    wire [31:0] SubBytesInput ;
    wire [3:0] SubBytesOutput ;
    wire [31:0] MixColumnsOutput ;
    wire [31:0] ColumnOutput ;
    wire [127:0] RoundKeyOutput ;
    wire [127:32] RoundKey ;
    wire [7:0] Rcon ;
    wire [127:0] KeyExpansionOutput ;
    wire [3:0] RoundCounter ;
    wire [2:0] InRoundCounter ;
    wire [28:0] MixColumnsIns_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4309 ;
    wire clk_gated ;

    /* cells in depth 0 */
    AND2_X1 U323 ( .A1 (n45), .A2 (n44), .ZN (AKSRnotDone) ) ;
    NOR2_X1 U324 ( .A1 (n60), .A2 (n49), .ZN (LastRoundorDone) ) ;
    AND2_X1 U325 ( .A1 (RoundCounter[0]), .A2 (LastRoundorDone), .ZN (done) ) ;
    INV_X1 U326 ( .A (RoundCounter[3]), .ZN (n60) ) ;
    NOR2_X1 U327 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (n45) ) ;
    INV_X1 U328 ( .A (RoundCounter[2]), .ZN (n46) ) ;
    NAND2_X1 U329 ( .A1 (RoundCounter[1]), .A2 (n46), .ZN (n49) ) ;
    NOR2_X1 U330 ( .A1 (done), .A2 (InRoundCounter[2]), .ZN (n44) ) ;
    INV_X1 U331 ( .A (RoundCounter[1]), .ZN (n55) ) ;
    NAND2_X1 U332 ( .A1 (n55), .A2 (n46), .ZN (n47) ) ;
    NOR2_X1 U333 ( .A1 (RoundCounter[0]), .A2 (n47), .ZN (Rcon[0]) ) ;
    NOR2_X1 U334 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n58) ) ;
    NOR2_X1 U335 ( .A1 (n58), .A2 (n47), .ZN (Rcon[1]) ) ;
    NOR2_X1 U336 ( .A1 (RoundCounter[3]), .A2 (n49), .ZN (n48) ) ;
    NOR2_X1 U337 ( .A1 (n60), .A2 (n47), .ZN (n54) ) ;
    MUX2_X1 U338 ( .S (RoundCounter[0]), .A (n48), .B (n54), .Z (Rcon[2]) ) ;
    INV_X1 U339 ( .A (RoundCounter[0]), .ZN (n50) ) ;
    NOR2_X1 U340 ( .A1 (n50), .A2 (n49), .ZN (n51) ) ;
    MUX2_X1 U341 ( .S (RoundCounter[3]), .A (n51), .B (Rcon[0]), .Z (Rcon[3]) ) ;
    NAND2_X1 U342 ( .A1 (RoundCounter[2]), .A2 (n58), .ZN (n52) ) ;
    NOR2_X1 U343 ( .A1 (RoundCounter[1]), .A2 (n52), .ZN (n53) ) ;
    OR2_X1 U344 ( .A1 (n54), .A2 (n53), .ZN (Rcon[4]) ) ;
    XNOR2_X1 U345 ( .A (RoundCounter[2]), .B (RoundCounter[3]), .ZN (n57) ) ;
    NAND2_X1 U346 ( .A1 (RoundCounter[0]), .A2 (n55), .ZN (n56) ) ;
    NOR2_X1 U347 ( .A1 (n57), .A2 (n56), .ZN (Rcon[5]) ) ;
    INV_X1 U348 ( .A (n58), .ZN (n59) ) ;
    NAND2_X1 U349 ( .A1 (RoundCounter[1]), .A2 (RoundCounter[2]), .ZN (n61) ) ;
    NOR2_X1 U350 ( .A1 (n59), .A2 (n61), .ZN (Rcon[6]) ) ;
    NAND2_X1 U351 ( .A1 (RoundCounter[0]), .A2 (n60), .ZN (n62) ) ;
    NOR2_X1 U352 ( .A1 (n62), .A2 (n61), .ZN (Rcon[7]) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U353 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_2339, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2340, ShiftRowsOutput[96]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U354 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_2342, RoundKey[100]}), .c ({new_AGEMA_signal_2343, ShiftRowsOutput[68]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U355 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_2345, RoundKey[101]}), .c ({new_AGEMA_signal_2346, ShiftRowsOutput[69]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U356 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_2348, RoundKey[102]}), .c ({new_AGEMA_signal_2349, ShiftRowsOutput[70]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U357 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_2351, RoundKey[103]}), .c ({new_AGEMA_signal_2352, ShiftRowsOutput[71]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U358 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_2354, RoundKey[104]}), .c ({new_AGEMA_signal_2355, ShiftRowsOutput[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U359 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_2357, RoundKey[105]}), .c ({new_AGEMA_signal_2358, ShiftRowsOutput[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U360 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_2360, RoundKey[106]}), .c ({new_AGEMA_signal_2361, ShiftRowsOutput[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U361 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_2363, RoundKey[107]}), .c ({new_AGEMA_signal_2364, ShiftRowsOutput[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U362 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_2366, RoundKey[108]}), .c ({new_AGEMA_signal_2367, ShiftRowsOutput[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U363 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_2369, RoundKey[109]}), .c ({new_AGEMA_signal_2370, ShiftRowsOutput[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U364 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({new_AGEMA_signal_2372, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2373, ShiftRowsOutput[74]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U365 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_2375, RoundKey[110]}), .c ({new_AGEMA_signal_2376, ShiftRowsOutput[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U366 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_2378, RoundKey[111]}), .c ({new_AGEMA_signal_2379, ShiftRowsOutput[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U367 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_2381, RoundKey[112]}), .c ({new_AGEMA_signal_2382, ShiftRowsOutput[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U368 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({new_AGEMA_signal_2384, RoundKey[113]}), .c ({new_AGEMA_signal_2385, ShiftRowsOutput[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U369 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({new_AGEMA_signal_2387, RoundKey[114]}), .c ({new_AGEMA_signal_2388, ShiftRowsOutput[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U370 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({new_AGEMA_signal_2390, RoundKey[115]}), .c ({new_AGEMA_signal_2391, ShiftRowsOutput[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U371 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({new_AGEMA_signal_2393, RoundKey[116]}), .c ({new_AGEMA_signal_2394, ShiftRowsOutput[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U372 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({new_AGEMA_signal_2396, RoundKey[117]}), .c ({new_AGEMA_signal_2397, ShiftRowsOutput[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U373 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({new_AGEMA_signal_2399, RoundKey[118]}), .c ({new_AGEMA_signal_2400, ShiftRowsOutput[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U374 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({new_AGEMA_signal_2402, RoundKey[119]}), .c ({new_AGEMA_signal_2403, ShiftRowsOutput[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U375 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({new_AGEMA_signal_2405, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2406, ShiftRowsOutput[75]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U376 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2408, RoundKey[120]}), .c ({new_AGEMA_signal_2409, ShiftRowsOutput[120]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U377 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2411, RoundKey[121]}), .c ({new_AGEMA_signal_2412, ShiftRowsOutput[121]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U378 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2414, RoundKey[122]}), .c ({new_AGEMA_signal_2415, ShiftRowsOutput[122]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U379 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2417, RoundKey[123]}), .c ({new_AGEMA_signal_2418, ShiftRowsOutput[123]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U380 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2420, RoundKey[124]}), .c ({new_AGEMA_signal_2421, ShiftRowsOutput[124]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U381 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2423, RoundKey[125]}), .c ({new_AGEMA_signal_2424, ShiftRowsOutput[125]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U382 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2426, RoundKey[126]}), .c ({new_AGEMA_signal_2427, ShiftRowsOutput[126]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U383 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2429, RoundKey[127]}), .c ({new_AGEMA_signal_2430, ShiftRowsOutput[127]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U384 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({new_AGEMA_signal_2432, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2433, ShiftRowsOutput[76]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U385 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({new_AGEMA_signal_2435, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2436, ShiftRowsOutput[77]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U386 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({new_AGEMA_signal_2438, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2439, ShiftRowsOutput[78]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U387 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({new_AGEMA_signal_2441, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2442, ShiftRowsOutput[79]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U388 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_2444, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2445, ShiftRowsOutput[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U389 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({new_AGEMA_signal_2447, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2448, ShiftRowsOutput[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U390 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({new_AGEMA_signal_2450, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2451, ShiftRowsOutput[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U391 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({new_AGEMA_signal_2453, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2454, ShiftRowsOutput[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U392 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_2456, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2457, ShiftRowsOutput[97]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U393 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({new_AGEMA_signal_2459, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2460, ShiftRowsOutput[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U394 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({new_AGEMA_signal_2462, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2463, ShiftRowsOutput[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U395 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({new_AGEMA_signal_2465, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2466, ShiftRowsOutput[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U396 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({new_AGEMA_signal_2468, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2469, ShiftRowsOutput[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U397 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2471, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2472, ShiftRowsOutput[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U398 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2474, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2475, ShiftRowsOutput[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U399 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_2477, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2478, ShiftRowsOutput[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U400 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2480, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2481, ShiftRowsOutput[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U401 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2483, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2484, ShiftRowsOutput[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U402 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2486, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2487, ShiftRowsOutput[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U403 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_2489, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2490, ShiftRowsOutput[98]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U404 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2492, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2493, ShiftRowsOutput[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U405 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2495, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2496, ShiftRowsOutput[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U406 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_2498, RoundKey[32]}), .c ({new_AGEMA_signal_2499, ShiftRowsOutput[0]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U407 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({new_AGEMA_signal_2501, RoundKey[33]}), .c ({new_AGEMA_signal_2502, ShiftRowsOutput[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U408 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({new_AGEMA_signal_2504, RoundKey[34]}), .c ({new_AGEMA_signal_2505, ShiftRowsOutput[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U409 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({new_AGEMA_signal_2507, RoundKey[35]}), .c ({new_AGEMA_signal_2508, ShiftRowsOutput[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U410 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({new_AGEMA_signal_2510, RoundKey[36]}), .c ({new_AGEMA_signal_2511, ShiftRowsOutput[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U411 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({new_AGEMA_signal_2513, RoundKey[37]}), .c ({new_AGEMA_signal_2514, ShiftRowsOutput[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U412 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({new_AGEMA_signal_2516, RoundKey[38]}), .c ({new_AGEMA_signal_2517, ShiftRowsOutput[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U413 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({new_AGEMA_signal_2519, RoundKey[39]}), .c ({new_AGEMA_signal_2520, ShiftRowsOutput[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U414 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_2522, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2523, ShiftRowsOutput[99]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U415 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_2525, RoundKey[40]}), .c ({new_AGEMA_signal_2526, ShiftRowsOutput[104]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U416 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({new_AGEMA_signal_2528, RoundKey[41]}), .c ({new_AGEMA_signal_2529, ShiftRowsOutput[105]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U417 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({new_AGEMA_signal_2531, RoundKey[42]}), .c ({new_AGEMA_signal_2532, ShiftRowsOutput[106]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U418 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({new_AGEMA_signal_2534, RoundKey[43]}), .c ({new_AGEMA_signal_2535, ShiftRowsOutput[107]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U419 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({new_AGEMA_signal_2537, RoundKey[44]}), .c ({new_AGEMA_signal_2538, ShiftRowsOutput[108]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U420 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({new_AGEMA_signal_2540, RoundKey[45]}), .c ({new_AGEMA_signal_2541, ShiftRowsOutput[109]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U421 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({new_AGEMA_signal_2543, RoundKey[46]}), .c ({new_AGEMA_signal_2544, ShiftRowsOutput[110]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U422 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({new_AGEMA_signal_2546, RoundKey[47]}), .c ({new_AGEMA_signal_2547, ShiftRowsOutput[111]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U423 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_2549, RoundKey[48]}), .c ({new_AGEMA_signal_2550, ShiftRowsOutput[80]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U424 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_2552, RoundKey[49]}), .c ({new_AGEMA_signal_2553, ShiftRowsOutput[81]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U425 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_2555, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2556, ShiftRowsOutput[100]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U426 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_2558, RoundKey[50]}), .c ({new_AGEMA_signal_2559, ShiftRowsOutput[82]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U427 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_2561, RoundKey[51]}), .c ({new_AGEMA_signal_2562, ShiftRowsOutput[83]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U428 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_2564, RoundKey[52]}), .c ({new_AGEMA_signal_2565, ShiftRowsOutput[84]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U429 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_2567, RoundKey[53]}), .c ({new_AGEMA_signal_2568, ShiftRowsOutput[85]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U430 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_2570, RoundKey[54]}), .c ({new_AGEMA_signal_2571, ShiftRowsOutput[86]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U431 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_2573, RoundKey[55]}), .c ({new_AGEMA_signal_2574, ShiftRowsOutput[87]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U432 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_2576, RoundKey[56]}), .c ({new_AGEMA_signal_2577, ShiftRowsOutput[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U433 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2579, RoundKey[57]}), .c ({new_AGEMA_signal_2580, ShiftRowsOutput[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U434 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_2582, RoundKey[58]}), .c ({new_AGEMA_signal_2583, ShiftRowsOutput[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U435 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2585, RoundKey[59]}), .c ({new_AGEMA_signal_2586, ShiftRowsOutput[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U436 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_2588, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_2589, ShiftRowsOutput[101]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U437 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2591, RoundKey[60]}), .c ({new_AGEMA_signal_2592, ShiftRowsOutput[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U438 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2594, RoundKey[61]}), .c ({new_AGEMA_signal_2595, ShiftRowsOutput[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U439 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2597, RoundKey[62]}), .c ({new_AGEMA_signal_2598, ShiftRowsOutput[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U440 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2600, RoundKey[63]}), .c ({new_AGEMA_signal_2601, ShiftRowsOutput[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U441 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_2603, RoundKey[64]}), .c ({new_AGEMA_signal_2604, ShiftRowsOutput[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U442 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({new_AGEMA_signal_2606, RoundKey[65]}), .c ({new_AGEMA_signal_2607, ShiftRowsOutput[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U443 ( .a ({ciphertext_s1[98], ciphertext_s0[98]}), .b ({new_AGEMA_signal_2609, RoundKey[66]}), .c ({new_AGEMA_signal_2610, ShiftRowsOutput[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U444 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({new_AGEMA_signal_2612, RoundKey[67]}), .c ({new_AGEMA_signal_2613, ShiftRowsOutput[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U445 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({new_AGEMA_signal_2615, RoundKey[68]}), .c ({new_AGEMA_signal_2616, ShiftRowsOutput[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U446 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({new_AGEMA_signal_2618, RoundKey[69]}), .c ({new_AGEMA_signal_2619, ShiftRowsOutput[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U447 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_2621, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_2622, ShiftRowsOutput[102]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U448 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({new_AGEMA_signal_2624, RoundKey[70]}), .c ({new_AGEMA_signal_2625, ShiftRowsOutput[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U449 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({new_AGEMA_signal_2627, RoundKey[71]}), .c ({new_AGEMA_signal_2628, ShiftRowsOutput[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U450 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_2630, RoundKey[72]}), .c ({new_AGEMA_signal_2631, ShiftRowsOutput[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U451 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_2633, RoundKey[73]}), .c ({new_AGEMA_signal_2634, ShiftRowsOutput[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U452 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_2636, RoundKey[74]}), .c ({new_AGEMA_signal_2637, ShiftRowsOutput[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U453 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_2639, RoundKey[75]}), .c ({new_AGEMA_signal_2640, ShiftRowsOutput[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U454 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_2642, RoundKey[76]}), .c ({new_AGEMA_signal_2643, ShiftRowsOutput[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U455 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_2645, RoundKey[77]}), .c ({new_AGEMA_signal_2646, ShiftRowsOutput[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U456 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_2648, RoundKey[78]}), .c ({new_AGEMA_signal_2649, ShiftRowsOutput[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U457 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_2651, RoundKey[79]}), .c ({new_AGEMA_signal_2652, ShiftRowsOutput[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U458 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_2654, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_2655, ShiftRowsOutput[103]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U459 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_2657, RoundKey[80]}), .c ({new_AGEMA_signal_2658, ShiftRowsOutput[112]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U460 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_2660, RoundKey[81]}), .c ({new_AGEMA_signal_2661, ShiftRowsOutput[113]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U461 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_2663, RoundKey[82]}), .c ({new_AGEMA_signal_2664, ShiftRowsOutput[114]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U462 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_2666, RoundKey[83]}), .c ({new_AGEMA_signal_2667, ShiftRowsOutput[115]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U463 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_2669, RoundKey[84]}), .c ({new_AGEMA_signal_2670, ShiftRowsOutput[116]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U464 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_2672, RoundKey[85]}), .c ({new_AGEMA_signal_2673, ShiftRowsOutput[117]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U465 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_2675, RoundKey[86]}), .c ({new_AGEMA_signal_2676, ShiftRowsOutput[118]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U466 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_2678, RoundKey[87]}), .c ({new_AGEMA_signal_2679, ShiftRowsOutput[119]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U467 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_2681, RoundKey[88]}), .c ({new_AGEMA_signal_2682, ShiftRowsOutput[88]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U468 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2684, RoundKey[89]}), .c ({new_AGEMA_signal_2685, ShiftRowsOutput[89]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U469 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_2687, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_2688, ShiftRowsOutput[72]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U470 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_2690, RoundKey[90]}), .c ({new_AGEMA_signal_2691, ShiftRowsOutput[90]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U471 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2693, RoundKey[91]}), .c ({new_AGEMA_signal_2694, ShiftRowsOutput[91]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U472 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2696, RoundKey[92]}), .c ({new_AGEMA_signal_2697, ShiftRowsOutput[92]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U473 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2699, RoundKey[93]}), .c ({new_AGEMA_signal_2700, ShiftRowsOutput[93]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U474 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2702, RoundKey[94]}), .c ({new_AGEMA_signal_2703, ShiftRowsOutput[94]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U475 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2705, RoundKey[95]}), .c ({new_AGEMA_signal_2706, ShiftRowsOutput[95]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U476 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_2708, RoundKey[96]}), .c ({new_AGEMA_signal_2709, ShiftRowsOutput[64]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U477 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_2711, RoundKey[97]}), .c ({new_AGEMA_signal_2712, ShiftRowsOutput[65]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U478 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_2714, RoundKey[98]}), .c ({new_AGEMA_signal_2715, ShiftRowsOutput[66]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U479 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_2717, RoundKey[99]}), .c ({new_AGEMA_signal_2718, ShiftRowsOutput[67]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) U480 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({new_AGEMA_signal_2720, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_2721, ShiftRowsOutput[73]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2754, RoundOutput[32]}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_2851, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2755, RoundOutput[33]}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_2853, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2756, RoundOutput[34]}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_2855, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2757, RoundOutput[35]}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_2857, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2758, RoundOutput[36]}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_2859, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2759, RoundOutput[37]}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_2861, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2760, RoundOutput[38]}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_2863, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2761, RoundOutput[39]}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_2865, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2762, RoundOutput[40]}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_2867, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2763, RoundOutput[41]}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_2869, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2764, RoundOutput[42]}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_2871, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2765, RoundOutput[43]}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_2873, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2766, RoundOutput[44]}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_2875, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2767, RoundOutput[45]}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_2877, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2768, RoundOutput[46]}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_2879, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2769, RoundOutput[47]}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_2881, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2770, RoundOutput[48]}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_2883, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2771, RoundOutput[49]}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_2885, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2772, RoundOutput[50]}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_2887, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2773, RoundOutput[51]}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_2889, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2774, RoundOutput[52]}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_2891, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2775, RoundOutput[53]}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_2893, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2776, RoundOutput[54]}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_2895, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2777, RoundOutput[55]}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_2897, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2778, RoundOutput[56]}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_2899, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2779, RoundOutput[57]}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_2901, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2780, RoundOutput[58]}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_2903, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2781, RoundOutput[59]}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_2905, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2782, RoundOutput[60]}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_2907, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2783, RoundOutput[61]}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_2909, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2784, RoundOutput[62]}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_2911, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2785, RoundOutput[63]}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_2913, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2786, RoundOutput[64]}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_2915, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2787, RoundOutput[65]}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_2917, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2788, RoundOutput[66]}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_2919, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2789, RoundOutput[67]}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_2921, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2790, RoundOutput[68]}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_2923, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2791, RoundOutput[69]}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_2925, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2792, RoundOutput[70]}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_2927, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2793, RoundOutput[71]}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_2929, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2794, RoundOutput[72]}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_2931, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2795, RoundOutput[73]}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_2933, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2796, RoundOutput[74]}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_2935, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2797, RoundOutput[75]}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_2937, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2798, RoundOutput[76]}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_2939, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2799, RoundOutput[77]}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_2941, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2800, RoundOutput[78]}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_2943, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2801, RoundOutput[79]}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_2945, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2802, RoundOutput[80]}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_2947, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2803, RoundOutput[81]}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_2949, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2804, RoundOutput[82]}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_2951, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2805, RoundOutput[83]}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_2953, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2806, RoundOutput[84]}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_2955, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2807, RoundOutput[85]}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_2957, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2808, RoundOutput[86]}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_2959, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2809, RoundOutput[87]}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_2961, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2810, RoundOutput[88]}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_2963, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2811, RoundOutput[89]}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_2965, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2812, RoundOutput[90]}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_2967, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2813, RoundOutput[91]}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_2969, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2814, RoundOutput[92]}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_2971, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2815, RoundOutput[93]}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_2973, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2816, RoundOutput[94]}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_2975, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2817, RoundOutput[95]}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_2977, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2818, RoundOutput[96]}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_2979, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2819, RoundOutput[97]}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_2981, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2820, RoundOutput[98]}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_2983, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2821, RoundOutput[99]}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_2985, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2822, RoundOutput[100]}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_2987, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2823, RoundOutput[101]}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_2989, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2824, RoundOutput[102]}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_2991, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2825, RoundOutput[103]}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_2993, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2826, RoundOutput[104]}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_2995, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2827, RoundOutput[105]}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_2997, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2828, RoundOutput[106]}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_2999, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2829, RoundOutput[107]}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_3001, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2830, RoundOutput[108]}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_3003, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2831, RoundOutput[109]}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_3005, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2832, RoundOutput[110]}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_3007, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2833, RoundOutput[111]}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_3009, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2834, RoundOutput[112]}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_3011, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2835, RoundOutput[113]}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_3013, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2836, RoundOutput[114]}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_3015, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2837, RoundOutput[115]}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_3017, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2838, RoundOutput[116]}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_3019, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2839, RoundOutput[117]}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_3021, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2840, RoundOutput[118]}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_3023, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2841, RoundOutput[119]}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_3025, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2842, RoundOutput[120]}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_3027, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2843, RoundOutput[121]}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_3029, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2844, RoundOutput[122]}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_3031, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2845, RoundOutput[123]}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_3033, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2846, RoundOutput[124]}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_3035, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2847, RoundOutput[125]}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_3037, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2848, RoundOutput[126]}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_3039, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2849, RoundOutput[127]}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_3041, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    INV_X1 MuxSboxIn_U3 ( .A (AKSRnotDone), .ZN (MuxSboxIn_n7) ) ;
    INV_X1 MuxSboxIn_U2 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n5) ) ;
    INV_X1 MuxSboxIn_U1 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n6) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_0_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .a ({new_AGEMA_signal_2444, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2723, SubBytesInput[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_1_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .a ({new_AGEMA_signal_2447, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2724, SubBytesInput[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_2_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .a ({new_AGEMA_signal_2450, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2725, SubBytesInput[2]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_3_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .a ({new_AGEMA_signal_2453, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2726, SubBytesInput[3]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_4_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .a ({new_AGEMA_signal_2459, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2727, SubBytesInput[4]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_5_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .a ({new_AGEMA_signal_2462, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2728, SubBytesInput[5]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_6_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .a ({new_AGEMA_signal_2465, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2729, SubBytesInput[6]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_7_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .a ({new_AGEMA_signal_2468, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2730, SubBytesInput[7]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_8_U1 ( .s (AKSRnotDone), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .a ({new_AGEMA_signal_2687, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_2722, SubBytesInput[8]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_9_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .a ({new_AGEMA_signal_2720, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_2731, SubBytesInput[9]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_10_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .a ({new_AGEMA_signal_2372, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2732, SubBytesInput[10]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_11_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .a ({new_AGEMA_signal_2405, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2733, SubBytesInput[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_12_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .a ({new_AGEMA_signal_2432, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2734, SubBytesInput[12]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_13_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .a ({new_AGEMA_signal_2435, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2735, SubBytesInput[13]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_14_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .a ({new_AGEMA_signal_2438, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2736, SubBytesInput[14]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_15_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .a ({new_AGEMA_signal_2441, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2737, SubBytesInput[15]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_16_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .a ({new_AGEMA_signal_2339, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2738, SubBytesInput[16]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_17_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .a ({new_AGEMA_signal_2456, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2739, SubBytesInput[17]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_18_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .a ({new_AGEMA_signal_2489, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2740, SubBytesInput[18]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_19_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .a ({new_AGEMA_signal_2522, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2741, SubBytesInput[19]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_20_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .a ({new_AGEMA_signal_2555, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2742, SubBytesInput[20]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_21_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .a ({new_AGEMA_signal_2588, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_2743, SubBytesInput[21]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_22_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .a ({new_AGEMA_signal_2621, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_2744, SubBytesInput[22]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_23_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .a ({new_AGEMA_signal_2654, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_2745, SubBytesInput[23]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_24_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .a ({new_AGEMA_signal_2471, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2746, SubBytesInput[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_25_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .a ({new_AGEMA_signal_2474, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2747, SubBytesInput[25]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_26_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .a ({new_AGEMA_signal_2477, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2748, SubBytesInput[26]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_27_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .a ({new_AGEMA_signal_2480, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2749, SubBytesInput[27]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_28_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .a ({new_AGEMA_signal_2483, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2750, SubBytesInput[28]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_29_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .a ({new_AGEMA_signal_2486, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2751, SubBytesInput[29]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_30_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .a ({new_AGEMA_signal_2492, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2752, SubBytesInput[30]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxSboxIn_mux_inst_31_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .a ({new_AGEMA_signal_2495, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2753, SubBytesInput[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_2730, SubBytesInput[7]}), .b ({new_AGEMA_signal_2727, SubBytesInput[4]}), .c ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_2730, SubBytesInput[7]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_2730, SubBytesInput[7]}), .b ({new_AGEMA_signal_2724, SubBytesInput[1]}), .c ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_2727, SubBytesInput[4]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_2726, SubBytesInput[3]}), .b ({new_AGEMA_signal_2724, SubBytesInput[1]}), .c ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_2729, SubBytesInput[6]}), .b ({new_AGEMA_signal_2728, SubBytesInput[5]}), .c ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_2723, SubBytesInput[0]}), .b ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_3114, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_2723, SubBytesInput[0]}), .b ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_2729, SubBytesInput[6]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3048, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_2728, SubBytesInput[5]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3049, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_3084, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3048, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3116, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3048, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3085, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3049, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_2727, SubBytesInput[4]}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .c ({new_AGEMA_signal_3050, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3050, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_2724, SubBytesInput[1]}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .c ({new_AGEMA_signal_3051, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3051, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_3119, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_3166, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_3167, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3120, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3049, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3089, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_2737, SubBytesInput[15]}), .b ({new_AGEMA_signal_2734, SubBytesInput[12]}), .c ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_2737, SubBytesInput[15]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_2737, SubBytesInput[15]}), .b ({new_AGEMA_signal_2731, SubBytesInput[9]}), .c ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_2734, SubBytesInput[12]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_2733, SubBytesInput[11]}), .b ({new_AGEMA_signal_2731, SubBytesInput[9]}), .c ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_2736, SubBytesInput[14]}), .b ({new_AGEMA_signal_2735, SubBytesInput[13]}), .c ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_2722, SubBytesInput[8]}), .b ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_3127, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_2722, SubBytesInput[8]}), .b ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_2736, SubBytesInput[14]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3058, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_2735, SubBytesInput[13]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3059, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_3092, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3058, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3129, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3058, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3093, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3059, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_2734, SubBytesInput[12]}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .c ({new_AGEMA_signal_3060, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3060, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_2731, SubBytesInput[9]}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .c ({new_AGEMA_signal_3061, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3061, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_3132, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_3175, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_3176, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3133, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3059, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3097, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_2745, SubBytesInput[23]}), .b ({new_AGEMA_signal_2742, SubBytesInput[20]}), .c ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_2745, SubBytesInput[23]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_2745, SubBytesInput[23]}), .b ({new_AGEMA_signal_2739, SubBytesInput[17]}), .c ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_2742, SubBytesInput[20]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_2741, SubBytesInput[19]}), .b ({new_AGEMA_signal_2739, SubBytesInput[17]}), .c ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_2744, SubBytesInput[22]}), .b ({new_AGEMA_signal_2743, SubBytesInput[21]}), .c ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_2738, SubBytesInput[16]}), .b ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_3140, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_2738, SubBytesInput[16]}), .b ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_2744, SubBytesInput[22]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3068, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_2743, SubBytesInput[21]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3069, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_3100, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3068, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3142, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3068, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3101, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3069, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_2742, SubBytesInput[20]}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .c ({new_AGEMA_signal_3070, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3070, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_2739, SubBytesInput[17]}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .c ({new_AGEMA_signal_3071, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3071, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_3145, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_3184, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_3185, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3146, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3069, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3105, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_2753, SubBytesInput[31]}), .b ({new_AGEMA_signal_2750, SubBytesInput[28]}), .c ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_2753, SubBytesInput[31]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_2753, SubBytesInput[31]}), .b ({new_AGEMA_signal_2747, SubBytesInput[25]}), .c ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_2750, SubBytesInput[28]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_2749, SubBytesInput[27]}), .b ({new_AGEMA_signal_2747, SubBytesInput[25]}), .c ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_2752, SubBytesInput[30]}), .b ({new_AGEMA_signal_2751, SubBytesInput[29]}), .c ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_2746, SubBytesInput[24]}), .b ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_3153, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_2746, SubBytesInput[24]}), .b ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_2752, SubBytesInput[30]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3078, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_2751, SubBytesInput[29]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3079, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_3108, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3078, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3155, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3078, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3109, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3079, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_2750, SubBytesInput[28]}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .c ({new_AGEMA_signal_3080, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3080, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_2747, SubBytesInput[25]}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .c ({new_AGEMA_signal_3081, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3081, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_3158, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_3193, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_3194, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3159, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3079, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3113, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    INV_X1 MuxMCOut_U3 ( .A (LastRoundorDone), .ZN (MuxMCOut_n6) ) ;
    INV_X1 MuxMCOut_U2 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n5) ) ;
    INV_X1 MuxMCOut_U1 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n4) ) ;
    INV_X1 MuxRound_U7 ( .A (AKSRnotDone), .ZN (MuxRound_n19) ) ;
    INV_X1 MuxRound_U6 ( .A (MuxRound_n19), .ZN (MuxRound_n16) ) ;
    INV_X1 MuxRound_U5 ( .A (MuxRound_n19), .ZN (MuxRound_n14) ) ;
    INV_X1 MuxRound_U4 ( .A (MuxRound_n19), .ZN (MuxRound_n13) ) ;
    INV_X1 MuxRound_U3 ( .A (MuxRound_n19), .ZN (MuxRound_n15) ) ;
    INV_X1 MuxRound_U2 ( .A (MuxRound_n19), .ZN (MuxRound_n18) ) ;
    INV_X1 MuxRound_U1 ( .A (MuxRound_n19), .ZN (MuxRound_n17) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_32_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .a ({new_AGEMA_signal_2604, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_2754, RoundOutput[32]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_33_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .a ({new_AGEMA_signal_2607, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_2755, RoundOutput[33]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_34_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .a ({new_AGEMA_signal_2610, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_2756, RoundOutput[34]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_35_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .a ({new_AGEMA_signal_2613, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_2757, RoundOutput[35]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_36_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .a ({new_AGEMA_signal_2616, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_2758, RoundOutput[36]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_37_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .a ({new_AGEMA_signal_2619, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_2759, RoundOutput[37]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_38_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .a ({new_AGEMA_signal_2625, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_2760, RoundOutput[38]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_39_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .a ({new_AGEMA_signal_2628, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_2761, RoundOutput[39]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_40_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .a ({new_AGEMA_signal_2355, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_2762, RoundOutput[40]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_41_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .a ({new_AGEMA_signal_2358, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_2763, RoundOutput[41]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_42_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .a ({new_AGEMA_signal_2361, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_2764, RoundOutput[42]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_43_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .a ({new_AGEMA_signal_2364, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_2765, RoundOutput[43]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_44_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .a ({new_AGEMA_signal_2367, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_2766, RoundOutput[44]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_45_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .a ({new_AGEMA_signal_2370, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_2767, RoundOutput[45]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_46_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .a ({new_AGEMA_signal_2376, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_2768, RoundOutput[46]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_47_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .a ({new_AGEMA_signal_2379, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_2769, RoundOutput[47]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_48_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .a ({new_AGEMA_signal_2445, ShiftRowsOutput[48]}), .c ({new_AGEMA_signal_2770, RoundOutput[48]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_49_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .a ({new_AGEMA_signal_2448, ShiftRowsOutput[49]}), .c ({new_AGEMA_signal_2771, RoundOutput[49]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_50_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .a ({new_AGEMA_signal_2451, ShiftRowsOutput[50]}), .c ({new_AGEMA_signal_2772, RoundOutput[50]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_51_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .a ({new_AGEMA_signal_2454, ShiftRowsOutput[51]}), .c ({new_AGEMA_signal_2773, RoundOutput[51]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_52_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .a ({new_AGEMA_signal_2460, ShiftRowsOutput[52]}), .c ({new_AGEMA_signal_2774, RoundOutput[52]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_53_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .a ({new_AGEMA_signal_2463, ShiftRowsOutput[53]}), .c ({new_AGEMA_signal_2775, RoundOutput[53]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_54_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .a ({new_AGEMA_signal_2466, ShiftRowsOutput[54]}), .c ({new_AGEMA_signal_2776, RoundOutput[54]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_55_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .a ({new_AGEMA_signal_2469, ShiftRowsOutput[55]}), .c ({new_AGEMA_signal_2777, RoundOutput[55]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_56_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_2577, ShiftRowsOutput[56]}), .c ({new_AGEMA_signal_2778, RoundOutput[56]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_57_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_2580, ShiftRowsOutput[57]}), .c ({new_AGEMA_signal_2779, RoundOutput[57]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_58_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_2583, ShiftRowsOutput[58]}), .c ({new_AGEMA_signal_2780, RoundOutput[58]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_59_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_2586, ShiftRowsOutput[59]}), .c ({new_AGEMA_signal_2781, RoundOutput[59]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_60_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_2592, ShiftRowsOutput[60]}), .c ({new_AGEMA_signal_2782, RoundOutput[60]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_61_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_2595, ShiftRowsOutput[61]}), .c ({new_AGEMA_signal_2783, RoundOutput[61]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_62_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_2598, ShiftRowsOutput[62]}), .c ({new_AGEMA_signal_2784, RoundOutput[62]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_63_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_2601, ShiftRowsOutput[63]}), .c ({new_AGEMA_signal_2785, RoundOutput[63]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_64_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .a ({new_AGEMA_signal_2709, ShiftRowsOutput[64]}), .c ({new_AGEMA_signal_2786, RoundOutput[64]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_65_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .a ({new_AGEMA_signal_2712, ShiftRowsOutput[65]}), .c ({new_AGEMA_signal_2787, RoundOutput[65]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_66_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .a ({new_AGEMA_signal_2715, ShiftRowsOutput[66]}), .c ({new_AGEMA_signal_2788, RoundOutput[66]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_67_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .a ({new_AGEMA_signal_2718, ShiftRowsOutput[67]}), .c ({new_AGEMA_signal_2789, RoundOutput[67]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_68_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .a ({new_AGEMA_signal_2343, ShiftRowsOutput[68]}), .c ({new_AGEMA_signal_2790, RoundOutput[68]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_69_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .a ({new_AGEMA_signal_2346, ShiftRowsOutput[69]}), .c ({new_AGEMA_signal_2791, RoundOutput[69]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_70_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .a ({new_AGEMA_signal_2349, ShiftRowsOutput[70]}), .c ({new_AGEMA_signal_2792, RoundOutput[70]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_71_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .a ({new_AGEMA_signal_2352, ShiftRowsOutput[71]}), .c ({new_AGEMA_signal_2793, RoundOutput[71]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_72_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .a ({new_AGEMA_signal_2688, ShiftRowsOutput[72]}), .c ({new_AGEMA_signal_2794, RoundOutput[72]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_73_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .a ({new_AGEMA_signal_2721, ShiftRowsOutput[73]}), .c ({new_AGEMA_signal_2795, RoundOutput[73]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_74_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .a ({new_AGEMA_signal_2373, ShiftRowsOutput[74]}), .c ({new_AGEMA_signal_2796, RoundOutput[74]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_75_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .a ({new_AGEMA_signal_2406, ShiftRowsOutput[75]}), .c ({new_AGEMA_signal_2797, RoundOutput[75]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_76_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .a ({new_AGEMA_signal_2433, ShiftRowsOutput[76]}), .c ({new_AGEMA_signal_2798, RoundOutput[76]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_77_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .a ({new_AGEMA_signal_2436, ShiftRowsOutput[77]}), .c ({new_AGEMA_signal_2799, RoundOutput[77]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_78_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .a ({new_AGEMA_signal_2439, ShiftRowsOutput[78]}), .c ({new_AGEMA_signal_2800, RoundOutput[78]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_79_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .a ({new_AGEMA_signal_2442, ShiftRowsOutput[79]}), .c ({new_AGEMA_signal_2801, RoundOutput[79]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_80_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .a ({new_AGEMA_signal_2550, ShiftRowsOutput[80]}), .c ({new_AGEMA_signal_2802, RoundOutput[80]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_81_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .a ({new_AGEMA_signal_2553, ShiftRowsOutput[81]}), .c ({new_AGEMA_signal_2803, RoundOutput[81]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_82_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .a ({new_AGEMA_signal_2559, ShiftRowsOutput[82]}), .c ({new_AGEMA_signal_2804, RoundOutput[82]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_83_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .a ({new_AGEMA_signal_2562, ShiftRowsOutput[83]}), .c ({new_AGEMA_signal_2805, RoundOutput[83]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_84_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .a ({new_AGEMA_signal_2565, ShiftRowsOutput[84]}), .c ({new_AGEMA_signal_2806, RoundOutput[84]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_85_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .a ({new_AGEMA_signal_2568, ShiftRowsOutput[85]}), .c ({new_AGEMA_signal_2807, RoundOutput[85]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_86_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .a ({new_AGEMA_signal_2571, ShiftRowsOutput[86]}), .c ({new_AGEMA_signal_2808, RoundOutput[86]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_87_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .a ({new_AGEMA_signal_2574, ShiftRowsOutput[87]}), .c ({new_AGEMA_signal_2809, RoundOutput[87]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_88_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_2682, ShiftRowsOutput[88]}), .c ({new_AGEMA_signal_2810, RoundOutput[88]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_89_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_2685, ShiftRowsOutput[89]}), .c ({new_AGEMA_signal_2811, RoundOutput[89]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_90_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_2691, ShiftRowsOutput[90]}), .c ({new_AGEMA_signal_2812, RoundOutput[90]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_91_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_2694, ShiftRowsOutput[91]}), .c ({new_AGEMA_signal_2813, RoundOutput[91]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_92_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_2697, ShiftRowsOutput[92]}), .c ({new_AGEMA_signal_2814, RoundOutput[92]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_93_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_2700, ShiftRowsOutput[93]}), .c ({new_AGEMA_signal_2815, RoundOutput[93]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_94_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_2703, ShiftRowsOutput[94]}), .c ({new_AGEMA_signal_2816, RoundOutput[94]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_95_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_2706, ShiftRowsOutput[95]}), .c ({new_AGEMA_signal_2817, RoundOutput[95]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_96_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .a ({new_AGEMA_signal_2340, ShiftRowsOutput[96]}), .c ({new_AGEMA_signal_2818, RoundOutput[96]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_97_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .a ({new_AGEMA_signal_2457, ShiftRowsOutput[97]}), .c ({new_AGEMA_signal_2819, RoundOutput[97]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_98_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .a ({new_AGEMA_signal_2490, ShiftRowsOutput[98]}), .c ({new_AGEMA_signal_2820, RoundOutput[98]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_99_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .a ({new_AGEMA_signal_2523, ShiftRowsOutput[99]}), .c ({new_AGEMA_signal_2821, RoundOutput[99]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_100_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .a ({new_AGEMA_signal_2556, ShiftRowsOutput[100]}), .c ({new_AGEMA_signal_2822, RoundOutput[100]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_101_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .a ({new_AGEMA_signal_2589, ShiftRowsOutput[101]}), .c ({new_AGEMA_signal_2823, RoundOutput[101]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_102_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .a ({new_AGEMA_signal_2622, ShiftRowsOutput[102]}), .c ({new_AGEMA_signal_2824, RoundOutput[102]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_103_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .a ({new_AGEMA_signal_2655, ShiftRowsOutput[103]}), .c ({new_AGEMA_signal_2825, RoundOutput[103]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_104_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .a ({new_AGEMA_signal_2526, ShiftRowsOutput[104]}), .c ({new_AGEMA_signal_2826, RoundOutput[104]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_105_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .a ({new_AGEMA_signal_2529, ShiftRowsOutput[105]}), .c ({new_AGEMA_signal_2827, RoundOutput[105]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_106_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .a ({new_AGEMA_signal_2532, ShiftRowsOutput[106]}), .c ({new_AGEMA_signal_2828, RoundOutput[106]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_107_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .a ({new_AGEMA_signal_2535, ShiftRowsOutput[107]}), .c ({new_AGEMA_signal_2829, RoundOutput[107]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_108_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .a ({new_AGEMA_signal_2538, ShiftRowsOutput[108]}), .c ({new_AGEMA_signal_2830, RoundOutput[108]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_109_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .a ({new_AGEMA_signal_2541, ShiftRowsOutput[109]}), .c ({new_AGEMA_signal_2831, RoundOutput[109]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_110_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .a ({new_AGEMA_signal_2544, ShiftRowsOutput[110]}), .c ({new_AGEMA_signal_2832, RoundOutput[110]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_111_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .a ({new_AGEMA_signal_2547, ShiftRowsOutput[111]}), .c ({new_AGEMA_signal_2833, RoundOutput[111]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_112_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .a ({new_AGEMA_signal_2658, ShiftRowsOutput[112]}), .c ({new_AGEMA_signal_2834, RoundOutput[112]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_113_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .a ({new_AGEMA_signal_2661, ShiftRowsOutput[113]}), .c ({new_AGEMA_signal_2835, RoundOutput[113]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_114_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .a ({new_AGEMA_signal_2664, ShiftRowsOutput[114]}), .c ({new_AGEMA_signal_2836, RoundOutput[114]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_115_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .a ({new_AGEMA_signal_2667, ShiftRowsOutput[115]}), .c ({new_AGEMA_signal_2837, RoundOutput[115]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_116_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .a ({new_AGEMA_signal_2670, ShiftRowsOutput[116]}), .c ({new_AGEMA_signal_2838, RoundOutput[116]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_117_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .a ({new_AGEMA_signal_2673, ShiftRowsOutput[117]}), .c ({new_AGEMA_signal_2839, RoundOutput[117]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_118_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .a ({new_AGEMA_signal_2676, ShiftRowsOutput[118]}), .c ({new_AGEMA_signal_2840, RoundOutput[118]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_119_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .a ({new_AGEMA_signal_2679, ShiftRowsOutput[119]}), .c ({new_AGEMA_signal_2841, RoundOutput[119]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_120_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2409, ShiftRowsOutput[120]}), .c ({new_AGEMA_signal_2842, RoundOutput[120]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_121_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2412, ShiftRowsOutput[121]}), .c ({new_AGEMA_signal_2843, RoundOutput[121]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_122_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2415, ShiftRowsOutput[122]}), .c ({new_AGEMA_signal_2844, RoundOutput[122]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_123_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2418, ShiftRowsOutput[123]}), .c ({new_AGEMA_signal_2845, RoundOutput[123]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_124_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2421, ShiftRowsOutput[124]}), .c ({new_AGEMA_signal_2846, RoundOutput[124]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_125_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2424, ShiftRowsOutput[125]}), .c ({new_AGEMA_signal_2847, RoundOutput[125]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_126_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2427, ShiftRowsOutput[126]}), .c ({new_AGEMA_signal_2848, RoundOutput[126]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_127_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2430, ShiftRowsOutput[127]}), .c ({new_AGEMA_signal_2849, RoundOutput[127]}) ) ;
    INV_X1 MuxKeyExpansion_U8 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n14) ) ;
    INV_X1 MuxKeyExpansion_U7 ( .A (AKSRnotDone), .ZN (MuxKeyExpansion_n21) ) ;
    INV_X1 MuxKeyExpansion_U6 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n16) ) ;
    INV_X1 MuxKeyExpansion_U5 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n17) ) ;
    INV_X1 MuxKeyExpansion_U4 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n18) ) ;
    INV_X1 MuxKeyExpansion_U3 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n19) ) ;
    INV_X1 MuxKeyExpansion_U2 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n20) ) ;
    INV_X1 MuxKeyExpansion_U1 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n15) ) ;
    NOR2_X1 RoundCounterIns_U11 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_n45) ) ;
    XNOR2_X1 RoundCounterIns_U10 ( .A (RoundCounter[0]), .B (AKSRnotDone), .ZN (RoundCounterIns_n10) ) ;
    NOR2_X1 RoundCounterIns_U9 ( .A1 (reset), .A2 (RoundCounterIns_n9), .ZN (RoundCounterIns_n44) ) ;
    XOR2_X1 RoundCounterIns_U8 ( .A (RoundCounter[1]), .B (RoundCounterIns_n8), .Z (RoundCounterIns_n9) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (reset), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n42) ) ;
    XOR2_X1 RoundCounterIns_U6 ( .A (RoundCounter[3]), .B (RoundCounterIns_n6), .Z (RoundCounterIns_n7) ) ;
    NAND2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounter[2]), .ZN (RoundCounterIns_n6) ) ;
    NOR2_X1 RoundCounterIns_U4 ( .A1 (reset), .A2 (RoundCounterIns_n4), .ZN (RoundCounterIns_n1) ) ;
    XNOR2_X1 RoundCounterIns_U3 ( .A (RoundCounter[2]), .B (RoundCounterIns_n5), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (RoundCounterIns_n2), .A2 (RoundCounterIns_n8), .ZN (RoundCounterIns_n5) ) ;
    NAND2_X1 RoundCounterIns_U1 ( .A1 (AKSRnotDone), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_n8) ) ;
    INV_X1 RoundCounterIns_count_reg_1__U1 ( .A (RoundCounter[1]), .ZN (RoundCounterIns_n2) ) ;
    NOR2_X1 InRoundCounterIns_U13 ( .A1 (reset), .A2 (InRoundCounterIns_n12), .ZN (InRoundCounterIns_n41) ) ;
    XOR2_X1 InRoundCounterIns_U12 ( .A (InRoundCounter[0]), .B (InRoundCounterIns_n11), .Z (InRoundCounterIns_n12) ) ;
    NAND2_X1 InRoundCounterIns_U11 ( .A1 (InRoundCounterIns_n10), .A2 (1'b1), .ZN (InRoundCounterIns_n11) ) ;
    NAND2_X1 InRoundCounterIns_U10 ( .A1 (InRoundCounterIns_n9), .A2 (InRoundCounter[2]), .ZN (InRoundCounterIns_n10) ) ;
    NAND2_X1 InRoundCounterIns_U9 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (InRoundCounterIns_n9) ) ;
    NOR2_X1 InRoundCounterIns_U8 ( .A1 (reset), .A2 (InRoundCounterIns_n8), .ZN (InRoundCounterIns_n40) ) ;
    MUX2_X1 InRoundCounterIns_U7 ( .S (InRoundCounter[1]), .A (InRoundCounterIns_n7), .B (InRoundCounterIns_n5), .Z (InRoundCounterIns_n8) ) ;
    NOR2_X1 InRoundCounterIns_U6 ( .A1 (reset), .A2 (InRoundCounterIns_n4), .ZN (InRoundCounterIns_n39) ) ;
    NOR2_X1 InRoundCounterIns_U5 ( .A1 (InRoundCounterIns_n3), .A2 (InRoundCounterIns_n2), .ZN (InRoundCounterIns_n4) ) ;
    NOR2_X1 InRoundCounterIns_U4 ( .A1 (InRoundCounterIns_n1), .A2 (InRoundCounterIns_n7), .ZN (InRoundCounterIns_n2) ) ;
    NAND2_X1 InRoundCounterIns_U3 ( .A1 (InRoundCounterIns_n5), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n7) ) ;
    AND2_X1 InRoundCounterIns_U2 ( .A1 (InRoundCounter[0]), .A2 (1'b1), .ZN (InRoundCounterIns_n5) ) ;
    NOR2_X1 InRoundCounterIns_U1 ( .A1 (1'b1), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n3) ) ;
    INV_X1 InRoundCounterIns_count_reg_1__U1 ( .A (InRoundCounter[1]), .ZN (InRoundCounterIns_n1) ) ;
    INV_X1 InRoundCounterIns_count_reg_2__U1 ( .A (InRoundCounter[2]), .ZN (InRoundCounterIns_n6) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_3084, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_3121, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_3119, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_3114, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_3168, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_3116, SubBytesIns_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_3121, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_3169, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_3122, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_3122, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_3121, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_3170, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_3123, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_3124, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_3120, SubBytesIns_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_3123, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_3171, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_3172, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_3172, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_3123, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_3202, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3085, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_3125, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_3089, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_3126, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_3126, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_3125, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_3173, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_3174, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_3174, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_3125, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_3203, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_3169, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_3168, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_3204, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_3170, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_3166, SubBytesIns_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_3205, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_3171, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_3124, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_3206, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_3202, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_3203, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_3222, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_3204, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_3173, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_3205, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_3203, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_3206, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_3173, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_3222, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_3167, SubBytesIns_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_3254, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_3240, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_3092, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_3134, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_3132, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_3127, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_3177, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_3129, SubBytesIns_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_3134, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_3178, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_3135, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_3135, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_3134, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_3179, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_3136, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_3137, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_3133, SubBytesIns_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_3136, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_3180, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_3181, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_3181, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_3136, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_3207, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3093, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_3138, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_3097, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_3139, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_3139, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_3138, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_3182, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_3183, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_3183, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_3138, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_3208, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_3178, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_3177, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_3209, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_3179, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_3175, SubBytesIns_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_3210, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_3180, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_3137, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_3211, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_3207, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_3208, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_3226, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_3209, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_3182, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_3210, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_3208, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_3211, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_3182, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_3226, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_3176, SubBytesIns_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_3259, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_3244, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_3100, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_3147, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_3145, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_3140, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_3186, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_3142, SubBytesIns_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_3147, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_3187, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_3148, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_3148, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_3147, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_3188, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_3149, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_3150, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_3146, SubBytesIns_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_3149, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_3189, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_3190, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_3190, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_3149, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_3212, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3101, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_3151, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_3105, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_3152, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_3152, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_3151, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_3191, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_3192, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_3192, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_3151, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_3213, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_3187, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_3186, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_3214, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_3188, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_3184, SubBytesIns_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_3215, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_3189, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_3150, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_3216, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_3212, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_3213, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_3230, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_3214, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_3191, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_3215, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_3213, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_3216, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_3191, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_3230, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_3185, SubBytesIns_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_3264, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_3248, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_3108, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_3160, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_3158, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_3153, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_3195, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_3155, SubBytesIns_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_3160, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_3196, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_3161, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_3161, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_3160, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_3197, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_3162, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_3163, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_3159, SubBytesIns_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_3162, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_3198, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_3199, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_3199, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_3162, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_3217, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3109, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_3164, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_3113, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r (Fresh[34]), .c ({new_AGEMA_signal_3165, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_3165, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_3164, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_3200, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r (Fresh[35]), .c ({new_AGEMA_signal_3201, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_3201, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_3164, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_3218, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_3196, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_3195, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_3219, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_3197, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_3193, SubBytesIns_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_3220, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_3198, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_3163, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_3221, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_3217, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_3218, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_3234, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_3219, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_3200, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_3220, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_3218, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_3221, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_3200, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_3234, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_3194, SubBytesIns_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_3269, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_3252, SubBytesIns_Inst_Sbox_3_M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r (Fresh[36]), .c ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3255, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3256, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r (Fresh[37]), .c ({new_AGEMA_signal_3257, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_3240, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3258, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r (Fresh[38]), .c ({new_AGEMA_signal_3241, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_3254, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3278, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r (Fresh[39]), .c ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3260, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3261, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r (Fresh[40]), .c ({new_AGEMA_signal_3262, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_3244, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3263, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r (Fresh[41]), .c ({new_AGEMA_signal_3245, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_3259, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3283, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r (Fresh[42]), .c ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3265, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3266, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r (Fresh[43]), .c ({new_AGEMA_signal_3267, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_3248, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3268, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r (Fresh[44]), .c ({new_AGEMA_signal_3249, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_3264, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3288, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r (Fresh[45]), .c ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3270, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3271, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r (Fresh[46]), .c ({new_AGEMA_signal_3272, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_3252, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3273, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r (Fresh[47]), .c ({new_AGEMA_signal_3253, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_3269, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3293, SubBytesIns_Inst_Sbox_3_M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_3256, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_3240, SubBytesIns_Inst_Sbox_0_M27}), .clk (clk), .r (Fresh[48]), .c ({new_AGEMA_signal_3274, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_3255, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_3254, SubBytesIns_Inst_Sbox_0_M24}), .clk (clk), .r (Fresh[49]), .c ({new_AGEMA_signal_3275, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_3240, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_3257, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r (Fresh[50]), .c ({new_AGEMA_signal_3276, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_3254, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_3241, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r (Fresh[51]), .c ({new_AGEMA_signal_3277, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_3274, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_3276, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_3258, SubBytesIns_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_3275, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_3277, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_3278, SubBytesIns_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_3312, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_3313, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_3358, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_3261, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_3244, SubBytesIns_Inst_Sbox_1_M27}), .clk (clk), .r (Fresh[52]), .c ({new_AGEMA_signal_3279, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_3260, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_3259, SubBytesIns_Inst_Sbox_1_M24}), .clk (clk), .r (Fresh[53]), .c ({new_AGEMA_signal_3280, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_3244, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_3262, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r (Fresh[54]), .c ({new_AGEMA_signal_3281, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_3259, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_3245, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r (Fresh[55]), .c ({new_AGEMA_signal_3282, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_3279, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_3281, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_3263, SubBytesIns_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_3280, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_3282, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_3283, SubBytesIns_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_3324, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_3325, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_3370, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_3266, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_3248, SubBytesIns_Inst_Sbox_2_M27}), .clk (clk), .r (Fresh[56]), .c ({new_AGEMA_signal_3284, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_3265, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_3264, SubBytesIns_Inst_Sbox_2_M24}), .clk (clk), .r (Fresh[57]), .c ({new_AGEMA_signal_3285, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_3248, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_3267, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r (Fresh[58]), .c ({new_AGEMA_signal_3286, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_3264, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_3249, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r (Fresh[59]), .c ({new_AGEMA_signal_3287, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_3284, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_3286, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_3268, SubBytesIns_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_3285, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_3287, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_3288, SubBytesIns_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_3336, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_3337, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_3382, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_3271, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_3252, SubBytesIns_Inst_Sbox_3_M27}), .clk (clk), .r (Fresh[60]), .c ({new_AGEMA_signal_3289, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_3270, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_3269, SubBytesIns_Inst_Sbox_3_M24}), .clk (clk), .r (Fresh[61]), .c ({new_AGEMA_signal_3290, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_3252, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_3272, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r (Fresh[62]), .c ({new_AGEMA_signal_3291, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_3269, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_3253, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r (Fresh[63]), .c ({new_AGEMA_signal_3292, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_3289, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_3291, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_3273, SubBytesIns_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_3290, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_3292, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_3293, SubBytesIns_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_3348, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_3349, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_3394, SubBytesIns_Inst_Sbox_3_M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4035, RoundOutput[0]}), .a ({plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_4156, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4195, RoundOutput[1]}), .a ({plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_4273, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4036, RoundOutput[2]}), .a ({plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_4158, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4196, RoundOutput[3]}), .a ({plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_4275, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4197, RoundOutput[4]}), .a ({plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_4277, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4037, RoundOutput[5]}), .a ({plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_4160, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4038, RoundOutput[6]}), .a ({plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_4162, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4039, RoundOutput[7]}), .a ({plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_4164, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4040, RoundOutput[8]}), .a ({plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_4166, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4198, RoundOutput[9]}), .a ({plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_4279, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4041, RoundOutput[10]}), .a ({plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_4168, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4199, RoundOutput[11]}), .a ({plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_4281, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4200, RoundOutput[12]}), .a ({plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_4283, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4042, RoundOutput[13]}), .a ({plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_4170, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4043, RoundOutput[14]}), .a ({plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_4172, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4044, RoundOutput[15]}), .a ({plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_4174, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4045, RoundOutput[16]}), .a ({plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_4176, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4201, RoundOutput[17]}), .a ({plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_4285, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4046, RoundOutput[18]}), .a ({plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_4178, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4202, RoundOutput[19]}), .a ({plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_4287, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4203, RoundOutput[20]}), .a ({plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_4289, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4047, RoundOutput[21]}), .a ({plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_4180, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4048, RoundOutput[22]}), .a ({plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_4182, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4049, RoundOutput[23]}), .a ({plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_4184, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4050, RoundOutput[24]}), .a ({plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_4186, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4204, RoundOutput[25]}), .a ({plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_4291, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4051, RoundOutput[26]}), .a ({plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_4188, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4205, RoundOutput[27]}), .a ({plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_4293, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4206, RoundOutput[28]}), .a ({plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_4295, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4052, RoundOutput[29]}), .a ({plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_4190, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4053, RoundOutput[30]}), .a ({plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_4192, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4054, RoundOutput[31]}), .a ({plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_4194, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_3313, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r (Fresh[64]), .c ({new_AGEMA_signal_3359, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_3114, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r (Fresh[65]), .c ({new_AGEMA_signal_3314, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .clk (clk), .r (Fresh[66]), .c ({new_AGEMA_signal_3315, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_3312, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r (Fresh[67]), .c ({new_AGEMA_signal_3360, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r (Fresh[68]), .c ({new_AGEMA_signal_3316, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r (Fresh[69]), .c ({new_AGEMA_signal_3317, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_3085, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r (Fresh[70]), .c ({new_AGEMA_signal_3361, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_3358, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_3089, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r (Fresh[71]), .c ({new_AGEMA_signal_3406, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r (Fresh[72]), .c ({new_AGEMA_signal_3362, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_3313, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_3084, SubBytesIns_Inst_Sbox_0_T13}), .clk (clk), .r (Fresh[73]), .c ({new_AGEMA_signal_3363, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_3119, SubBytesIns_Inst_Sbox_0_T23}), .clk (clk), .r (Fresh[74]), .c ({new_AGEMA_signal_3318, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}), .clk (clk), .r (Fresh[75]), .c ({new_AGEMA_signal_3319, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_3312, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .clk (clk), .r (Fresh[76]), .c ({new_AGEMA_signal_3364, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}), .clk (clk), .r (Fresh[77]), .c ({new_AGEMA_signal_3320, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}), .clk (clk), .r (Fresh[78]), .c ({new_AGEMA_signal_3321, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .clk (clk), .r (Fresh[79]), .c ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_3358, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}), .clk (clk), .r (Fresh[80]), .c ({new_AGEMA_signal_3407, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .clk (clk), .r (Fresh[81]), .c ({new_AGEMA_signal_3366, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_3407, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_3316, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_3318, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_3359, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_3315, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_3408, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_3314, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_3363, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_3409, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_3362, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_3364, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_3410, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_3360, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_3411, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_3407, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_3411, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_3359, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_3409, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_3448, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_3317, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_3320, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_3368, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_3361, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_3406, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_3449, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_3406, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_3410, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_3450, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_3321, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_3408, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_3451, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_3315, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_3317, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_3369, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_3316, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_3482, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_3361, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_3412, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_3363, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_3413, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_3318, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_3483, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_3319, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_3414, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_3364, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_3368, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_3415, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_3366, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_3410, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_3452, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_3484, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_3448, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_3485, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_3409, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_3369, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_3453, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_3415, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_3408, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_3454, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_3413, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_3449, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_3486, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3450, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_3487, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_3448, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_3449, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_3488, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_3368, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_3450, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_3489, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_3451, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_3412, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_3490, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_3451, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_3414, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_3491, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3486, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_3483, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_3488, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_3452, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_3490, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3485, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_3484, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_3453, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_3530, SubBytesOutput[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_3487, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_3491, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_3531, SubBytesOutput[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_3482, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_3489, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3454, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_3492, SubBytesOutput[0]}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_3325, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r (Fresh[82]), .c ({new_AGEMA_signal_3371, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_3127, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r (Fresh[83]), .c ({new_AGEMA_signal_3326, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .clk (clk), .r (Fresh[84]), .c ({new_AGEMA_signal_3327, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_3324, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r (Fresh[85]), .c ({new_AGEMA_signal_3372, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r (Fresh[86]), .c ({new_AGEMA_signal_3328, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r (Fresh[87]), .c ({new_AGEMA_signal_3329, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_3093, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r (Fresh[88]), .c ({new_AGEMA_signal_3373, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_3370, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_3097, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r (Fresh[89]), .c ({new_AGEMA_signal_3416, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r (Fresh[90]), .c ({new_AGEMA_signal_3374, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_3325, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_3092, SubBytesIns_Inst_Sbox_1_T13}), .clk (clk), .r (Fresh[91]), .c ({new_AGEMA_signal_3375, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_3132, SubBytesIns_Inst_Sbox_1_T23}), .clk (clk), .r (Fresh[92]), .c ({new_AGEMA_signal_3330, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}), .clk (clk), .r (Fresh[93]), .c ({new_AGEMA_signal_3331, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_3324, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .clk (clk), .r (Fresh[94]), .c ({new_AGEMA_signal_3376, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}), .clk (clk), .r (Fresh[95]), .c ({new_AGEMA_signal_3332, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}), .clk (clk), .r (Fresh[96]), .c ({new_AGEMA_signal_3333, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .clk (clk), .r (Fresh[97]), .c ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_3370, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}), .clk (clk), .r (Fresh[98]), .c ({new_AGEMA_signal_3417, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .clk (clk), .r (Fresh[99]), .c ({new_AGEMA_signal_3378, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_3417, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_3328, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_3330, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_3371, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_3327, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_3418, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_3326, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_3375, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_3419, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_3374, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_3376, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_3420, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_3372, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_3421, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_3417, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_3421, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_3371, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_3419, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_3457, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_3329, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_3332, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_3380, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_3373, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_3416, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_3458, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_3416, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_3420, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_3459, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_3333, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_3418, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_3460, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_3327, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_3329, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_3381, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_3328, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_3493, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_3373, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_3422, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_3375, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_3423, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_3330, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_3494, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_3331, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_3424, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_3376, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_3380, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_3425, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_3378, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_3420, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_3461, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_3495, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_3457, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_3496, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_3419, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_3381, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_3462, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_3425, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_3418, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_3463, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_3423, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_3458, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_3497, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3459, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_3498, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_3457, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_3458, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_3499, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_3380, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_3459, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_3500, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_3460, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_3422, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_3501, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_3460, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_3424, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_3502, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3497, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_3494, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_3499, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_3461, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_3501, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3496, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_3495, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_3462, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_3498, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_3502, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_3493, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_3500, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3463, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_3337, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r (Fresh[100]), .c ({new_AGEMA_signal_3383, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_3140, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r (Fresh[101]), .c ({new_AGEMA_signal_3338, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .clk (clk), .r (Fresh[102]), .c ({new_AGEMA_signal_3339, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_3336, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r (Fresh[103]), .c ({new_AGEMA_signal_3384, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r (Fresh[104]), .c ({new_AGEMA_signal_3340, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r (Fresh[105]), .c ({new_AGEMA_signal_3341, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_3101, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r (Fresh[106]), .c ({new_AGEMA_signal_3385, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_3382, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_3105, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r (Fresh[107]), .c ({new_AGEMA_signal_3426, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r (Fresh[108]), .c ({new_AGEMA_signal_3386, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_3337, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_3100, SubBytesIns_Inst_Sbox_2_T13}), .clk (clk), .r (Fresh[109]), .c ({new_AGEMA_signal_3387, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_3145, SubBytesIns_Inst_Sbox_2_T23}), .clk (clk), .r (Fresh[110]), .c ({new_AGEMA_signal_3342, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}), .clk (clk), .r (Fresh[111]), .c ({new_AGEMA_signal_3343, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_3336, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .clk (clk), .r (Fresh[112]), .c ({new_AGEMA_signal_3388, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}), .clk (clk), .r (Fresh[113]), .c ({new_AGEMA_signal_3344, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}), .clk (clk), .r (Fresh[114]), .c ({new_AGEMA_signal_3345, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .clk (clk), .r (Fresh[115]), .c ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_3382, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}), .clk (clk), .r (Fresh[116]), .c ({new_AGEMA_signal_3427, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .clk (clk), .r (Fresh[117]), .c ({new_AGEMA_signal_3390, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_3427, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_3340, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_3342, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_3383, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_3339, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_3428, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_3338, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_3387, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_3429, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_3386, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_3388, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_3430, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_3384, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_3431, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_3427, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_3431, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_3383, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_3429, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_3466, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_3341, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_3344, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_3392, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_3385, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_3426, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_3467, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_3426, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_3430, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_3468, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_3345, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_3428, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_3469, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_3339, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_3341, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_3393, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_3340, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_3504, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_3385, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_3432, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_3387, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_3433, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_3342, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_3505, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_3343, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_3434, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_3388, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_3392, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_3435, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_3390, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_3430, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_3470, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_3506, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_3466, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_3507, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_3429, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_3393, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_3471, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_3435, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_3428, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_3472, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_3433, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_3467, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_3508, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3468, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_3509, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_3466, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_3467, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_3510, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_3392, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_3468, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_3511, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_3469, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_3432, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_3512, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_3469, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_3434, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_3513, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3508, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_3505, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_3510, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_3470, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_3512, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3507, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_3506, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_3471, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_3509, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_3513, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_3504, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_3511, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3472, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_3349, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r (Fresh[118]), .c ({new_AGEMA_signal_3395, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_3153, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r (Fresh[119]), .c ({new_AGEMA_signal_3350, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .clk (clk), .r (Fresh[120]), .c ({new_AGEMA_signal_3351, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_3348, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r (Fresh[121]), .c ({new_AGEMA_signal_3396, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r (Fresh[122]), .c ({new_AGEMA_signal_3352, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r (Fresh[123]), .c ({new_AGEMA_signal_3353, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_3109, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r (Fresh[124]), .c ({new_AGEMA_signal_3397, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_3394, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_3113, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r (Fresh[125]), .c ({new_AGEMA_signal_3436, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r (Fresh[126]), .c ({new_AGEMA_signal_3398, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_3349, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_3108, SubBytesIns_Inst_Sbox_3_T13}), .clk (clk), .r (Fresh[127]), .c ({new_AGEMA_signal_3399, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_3158, SubBytesIns_Inst_Sbox_3_T23}), .clk (clk), .r (Fresh[128]), .c ({new_AGEMA_signal_3354, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}), .clk (clk), .r (Fresh[129]), .c ({new_AGEMA_signal_3355, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_3348, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .clk (clk), .r (Fresh[130]), .c ({new_AGEMA_signal_3400, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}), .clk (clk), .r (Fresh[131]), .c ({new_AGEMA_signal_3356, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}), .clk (clk), .r (Fresh[132]), .c ({new_AGEMA_signal_3357, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .clk (clk), .r (Fresh[133]), .c ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_3394, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}), .clk (clk), .r (Fresh[134]), .c ({new_AGEMA_signal_3437, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .clk (clk), .r (Fresh[135]), .c ({new_AGEMA_signal_3402, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_3437, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_3352, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_3354, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_3395, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_3351, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_3438, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_3350, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_3399, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_3439, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_3398, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_3400, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_3440, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_3396, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_3441, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_3437, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_3441, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_3395, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_3439, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_3475, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_3353, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_3356, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_3404, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_3397, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_3436, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_3476, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_3436, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_3440, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_3477, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_3357, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_3438, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_3478, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_3351, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_3353, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_3405, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_3352, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_3515, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_3397, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_3442, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_3399, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_3443, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_3354, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_3516, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_3355, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_3444, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_3400, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_3404, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_3445, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_3402, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_3440, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_3479, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_3517, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_3475, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_3518, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_3439, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_3405, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_3480, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_3445, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_3438, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_3481, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_3443, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_3476, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_3519, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3477, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_3520, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_3475, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_3476, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_3521, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_3404, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_3477, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_3522, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_3478, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_3442, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_3523, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_3478, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_3444, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_3524, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3519, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_3516, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_3521, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_3479, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_3523, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3518, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_3517, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_3480, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_3520, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_3524, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_3515, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_3522, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3481, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U96 ( .a ({new_AGEMA_signal_3720, MixColumnsIns_n64}), .b ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_3866, MixColumnsOutput[9]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U95 ( .a ({new_AGEMA_signal_3646, MixColumnsIns_n63}), .b ({new_AGEMA_signal_3642, MixColumnsIns_n62}), .c ({new_AGEMA_signal_3720, MixColumnsIns_n64}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U94 ( .a ({new_AGEMA_signal_3625, MixColumnsIns_n61}), .b ({new_AGEMA_signal_3567, MixColumnsIns_n60}), .c ({new_AGEMA_signal_3721, MixColumnsOutput[8]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U93 ( .a ({new_AGEMA_signal_3577, MixColumnsIns_n59}), .b ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3625, MixColumnsIns_n61}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U92 ( .a ({new_AGEMA_signal_3626, MixColumnsIns_n58}), .b ({new_AGEMA_signal_3558, MixColumnsIns_n57}), .c ({new_AGEMA_signal_3722, MixColumnsOutput[7]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U91 ( .a ({new_AGEMA_signal_3569, MixColumnsIns_n56}), .b ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_3626, MixColumnsIns_n58}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U90 ( .a ({new_AGEMA_signal_3627, MixColumnsIns_n55}), .b ({new_AGEMA_signal_3559, MixColumnsIns_n54}), .c ({new_AGEMA_signal_3723, MixColumnsOutput[6]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U89 ( .a ({new_AGEMA_signal_3571, MixColumnsIns_n53}), .b ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3627, MixColumnsIns_n55}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U88 ( .a ({new_AGEMA_signal_3628, MixColumnsIns_n52}), .b ({new_AGEMA_signal_3560, MixColumnsIns_n51}), .c ({new_AGEMA_signal_3724, MixColumnsOutput[5]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U87 ( .a ({new_AGEMA_signal_3573, MixColumnsIns_n50}), .b ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3628, MixColumnsIns_n52}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U86 ( .a ({new_AGEMA_signal_3725, MixColumnsIns_n49}), .b ({new_AGEMA_signal_3633, MixColumnsIns_n48}), .c ({new_AGEMA_signal_3867, MixColumnsOutput[4]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U85 ( .a ({new_AGEMA_signal_3652, MixColumnsIns_n47}), .b ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_3725, MixColumnsIns_n49}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U84 ( .a ({new_AGEMA_signal_3726, MixColumnsIns_n46}), .b ({new_AGEMA_signal_3634, MixColumnsIns_n45}), .c ({new_AGEMA_signal_3868, MixColumnsOutput[3]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U83 ( .a ({new_AGEMA_signal_3654, MixColumnsIns_n44}), .b ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_3726, MixColumnsIns_n46}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U82 ( .a ({new_AGEMA_signal_3629, MixColumnsIns_n43}), .b ({new_AGEMA_signal_3558, MixColumnsIns_n57}), .c ({new_AGEMA_signal_3727, MixColumnsOutput[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U81 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3558, MixColumnsIns_n57}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U80 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3562, MixColumnsIns_n42}), .c ({new_AGEMA_signal_3629, MixColumnsIns_n43}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U79 ( .a ({new_AGEMA_signal_3630, MixColumnsIns_n41}), .b ({new_AGEMA_signal_3559, MixColumnsIns_n54}), .c ({new_AGEMA_signal_3728, MixColumnsOutput[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U78 ( .a ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .b ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3559, MixColumnsIns_n54}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U77 ( .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_3563, MixColumnsIns_n40}), .c ({new_AGEMA_signal_3630, MixColumnsIns_n41}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U76 ( .a ({new_AGEMA_signal_3631, MixColumnsIns_n39}), .b ({new_AGEMA_signal_3561, MixColumnsIns_n38}), .c ({new_AGEMA_signal_3729, MixColumnsOutput[2]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U75 ( .a ({new_AGEMA_signal_3575, MixColumnsIns_n37}), .b ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3631, MixColumnsIns_n39}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U74 ( .a ({new_AGEMA_signal_3632, MixColumnsIns_n36}), .b ({new_AGEMA_signal_3560, MixColumnsIns_n51}), .c ({new_AGEMA_signal_3730, MixColumnsOutput[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U73 ( .a ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .b ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_3560, MixColumnsIns_n51}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U72 ( .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_3564, MixColumnsIns_n35}), .c ({new_AGEMA_signal_3632, MixColumnsIns_n36}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U71 ( .a ({new_AGEMA_signal_3731, MixColumnsIns_n34}), .b ({new_AGEMA_signal_3633, MixColumnsIns_n48}), .c ({new_AGEMA_signal_3869, MixColumnsOutput[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U70 ( .a ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .b ({new_AGEMA_signal_3578, MixColumnsIns_DoubleBytes[28]}), .c ({new_AGEMA_signal_3633, MixColumnsIns_n48}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U69 ( .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_3640, MixColumnsIns_n33}), .c ({new_AGEMA_signal_3731, MixColumnsIns_n34}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U68 ( .a ({new_AGEMA_signal_3732, MixColumnsIns_n32}), .b ({new_AGEMA_signal_3634, MixColumnsIns_n45}), .c ({new_AGEMA_signal_3870, MixColumnsOutput[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U67 ( .a ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .b ({new_AGEMA_signal_3579, MixColumnsIns_DoubleBytes[27]}), .c ({new_AGEMA_signal_3634, MixColumnsIns_n45}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U66 ( .a ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .b ({new_AGEMA_signal_3643, MixColumnsIns_n31}), .c ({new_AGEMA_signal_3732, MixColumnsIns_n32}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U65 ( .a ({new_AGEMA_signal_3635, MixColumnsIns_n30}), .b ({new_AGEMA_signal_3561, MixColumnsIns_n38}), .c ({new_AGEMA_signal_3733, MixColumnsOutput[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U64 ( .a ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .b ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_3561, MixColumnsIns_n38}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U63 ( .a ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .b ({new_AGEMA_signal_3565, MixColumnsIns_n29}), .c ({new_AGEMA_signal_3635, MixColumnsIns_n30}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U62 ( .a ({new_AGEMA_signal_3734, MixColumnsIns_n28}), .b ({new_AGEMA_signal_3641, MixColumnsIns_n27}), .c ({new_AGEMA_signal_3871, MixColumnsOutput[25]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U61 ( .a ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_3645, MixColumnsIns_n26}), .c ({new_AGEMA_signal_3734, MixColumnsIns_n28}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U60 ( .a ({new_AGEMA_signal_3636, MixColumnsIns_n25}), .b ({new_AGEMA_signal_3566, MixColumnsIns_n24}), .c ({new_AGEMA_signal_3735, MixColumnsOutput[24]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U59 ( .a ({new_AGEMA_signal_3576, MixColumnsIns_n23}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3636, MixColumnsIns_n25}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U58 ( .a ({new_AGEMA_signal_3637, MixColumnsIns_n22}), .b ({new_AGEMA_signal_3562, MixColumnsIns_n42}), .c ({new_AGEMA_signal_3736, MixColumnsOutput[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U57 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3562, MixColumnsIns_n42}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U56 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3568, MixColumnsIns_n21}), .c ({new_AGEMA_signal_3637, MixColumnsIns_n22}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U55 ( .a ({new_AGEMA_signal_3638, MixColumnsIns_n20}), .b ({new_AGEMA_signal_3563, MixColumnsIns_n40}), .c ({new_AGEMA_signal_3737, MixColumnsOutput[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U54 ( .a ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .b ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3563, MixColumnsIns_n40}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U53 ( .a ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .b ({new_AGEMA_signal_3570, MixColumnsIns_n19}), .c ({new_AGEMA_signal_3638, MixColumnsIns_n20}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U52 ( .a ({new_AGEMA_signal_3639, MixColumnsIns_n18}), .b ({new_AGEMA_signal_3564, MixColumnsIns_n35}), .c ({new_AGEMA_signal_3738, MixColumnsOutput[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U51 ( .a ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .b ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_3564, MixColumnsIns_n35}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U50 ( .a ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .b ({new_AGEMA_signal_3572, MixColumnsIns_n17}), .c ({new_AGEMA_signal_3639, MixColumnsIns_n18}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U49 ( .a ({new_AGEMA_signal_3739, MixColumnsIns_n16}), .b ({new_AGEMA_signal_3640, MixColumnsIns_n33}), .c ({new_AGEMA_signal_3872, MixColumnsOutput[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U48 ( .a ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .b ({new_AGEMA_signal_3581, MixColumnsIns_DoubleBytes[20]}), .c ({new_AGEMA_signal_3640, MixColumnsIns_n33}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U47 ( .a ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .b ({new_AGEMA_signal_3651, MixColumnsIns_n15}), .c ({new_AGEMA_signal_3739, MixColumnsIns_n16}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U46 ( .a ({new_AGEMA_signal_3740, MixColumnsIns_n14}), .b ({new_AGEMA_signal_3641, MixColumnsIns_n27}), .c ({new_AGEMA_signal_3873, MixColumnsOutput[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U45 ( .a ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .b ({new_AGEMA_signal_3580, MixColumnsIns_DoubleBytes[25]}), .c ({new_AGEMA_signal_3641, MixColumnsIns_n27}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U44 ( .a ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .b ({new_AGEMA_signal_3642, MixColumnsIns_n62}), .c ({new_AGEMA_signal_3740, MixColumnsIns_n14}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U43 ( .a ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .b ({new_AGEMA_signal_3589, MixColumnsIns_DoubleBytes[1]}), .c ({new_AGEMA_signal_3642, MixColumnsIns_n62}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U42 ( .a ({new_AGEMA_signal_3741, MixColumnsIns_n13}), .b ({new_AGEMA_signal_3643, MixColumnsIns_n31}), .c ({new_AGEMA_signal_3874, MixColumnsOutput[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U41 ( .a ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .b ({new_AGEMA_signal_3582, MixColumnsIns_DoubleBytes[19]}), .c ({new_AGEMA_signal_3643, MixColumnsIns_n31}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U40 ( .a ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .b ({new_AGEMA_signal_3653, MixColumnsIns_n12}), .c ({new_AGEMA_signal_3741, MixColumnsIns_n13}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U39 ( .a ({new_AGEMA_signal_3644, MixColumnsIns_n11}), .b ({new_AGEMA_signal_3565, MixColumnsIns_n29}), .c ({new_AGEMA_signal_3742, MixColumnsOutput[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U38 ( .a ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .b ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_3565, MixColumnsIns_n29}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U37 ( .a ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .b ({new_AGEMA_signal_3574, MixColumnsIns_n10}), .c ({new_AGEMA_signal_3644, MixColumnsIns_n11}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U36 ( .a ({new_AGEMA_signal_3743, MixColumnsIns_n9}), .b ({new_AGEMA_signal_3645, MixColumnsIns_n26}), .c ({new_AGEMA_signal_3875, MixColumnsOutput[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U35 ( .a ({new_AGEMA_signal_3583, MixColumnsIns_DoubleBytes[17]}), .b ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_3645, MixColumnsIns_n26}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U34 ( .a ({new_AGEMA_signal_3646, MixColumnsIns_n63}), .b ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_3743, MixColumnsIns_n9}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U33 ( .a ({new_AGEMA_signal_3586, MixColumnsIns_DoubleBytes[9]}), .b ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_3646, MixColumnsIns_n63}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U32 ( .a ({new_AGEMA_signal_3647, MixColumnsIns_n8}), .b ({new_AGEMA_signal_3566, MixColumnsIns_n24}), .c ({new_AGEMA_signal_3744, MixColumnsOutput[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U31 ( .a ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .b ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3566, MixColumnsIns_n24}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U30 ( .a ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .b ({new_AGEMA_signal_3567, MixColumnsIns_n60}), .c ({new_AGEMA_signal_3647, MixColumnsIns_n8}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U29 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3567, MixColumnsIns_n60}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U28 ( .a ({new_AGEMA_signal_3648, MixColumnsIns_n7}), .b ({new_AGEMA_signal_3568, MixColumnsIns_n21}), .c ({new_AGEMA_signal_3745, MixColumnsOutput[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U27 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3568, MixColumnsIns_n21}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U26 ( .a ({new_AGEMA_signal_3569, MixColumnsIns_n56}), .b ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3648, MixColumnsIns_n7}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U25 ( .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3569, MixColumnsIns_n56}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U24 ( .a ({new_AGEMA_signal_3649, MixColumnsIns_n6}), .b ({new_AGEMA_signal_3570, MixColumnsIns_n19}), .c ({new_AGEMA_signal_3746, MixColumnsOutput[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U23 ( .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3570, MixColumnsIns_n19}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U22 ( .a ({new_AGEMA_signal_3571, MixColumnsIns_n53}), .b ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3649, MixColumnsIns_n6}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U21 ( .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3571, MixColumnsIns_n53}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U20 ( .a ({new_AGEMA_signal_3650, MixColumnsIns_n5}), .b ({new_AGEMA_signal_3572, MixColumnsIns_n17}), .c ({new_AGEMA_signal_3747, MixColumnsOutput[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U19 ( .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_3572, MixColumnsIns_n17}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U18 ( .a ({new_AGEMA_signal_3573, MixColumnsIns_n50}), .b ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3650, MixColumnsIns_n5}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U17 ( .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3573, MixColumnsIns_n50}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U16 ( .a ({new_AGEMA_signal_3748, MixColumnsIns_n4}), .b ({new_AGEMA_signal_3651, MixColumnsIns_n15}), .c ({new_AGEMA_signal_3876, MixColumnsOutput[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U15 ( .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_3584, MixColumnsIns_DoubleBytes[12]}), .c ({new_AGEMA_signal_3651, MixColumnsIns_n15}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U14 ( .a ({new_AGEMA_signal_3652, MixColumnsIns_n47}), .b ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_3748, MixColumnsIns_n4}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U13 ( .a ({new_AGEMA_signal_3587, MixColumnsIns_DoubleBytes[4]}), .b ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_3652, MixColumnsIns_n47}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U12 ( .a ({new_AGEMA_signal_3749, MixColumnsIns_n3}), .b ({new_AGEMA_signal_3653, MixColumnsIns_n12}), .c ({new_AGEMA_signal_3877, MixColumnsOutput[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U11 ( .a ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .b ({new_AGEMA_signal_3585, MixColumnsIns_DoubleBytes[11]}), .c ({new_AGEMA_signal_3653, MixColumnsIns_n12}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U10 ( .a ({new_AGEMA_signal_3654, MixColumnsIns_n44}), .b ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_3749, MixColumnsIns_n3}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U9 ( .a ({new_AGEMA_signal_3588, MixColumnsIns_DoubleBytes[3]}), .b ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_3654, MixColumnsIns_n44}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U8 ( .a ({new_AGEMA_signal_3655, MixColumnsIns_n2}), .b ({new_AGEMA_signal_3574, MixColumnsIns_n10}), .c ({new_AGEMA_signal_3750, MixColumnsOutput[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U7 ( .a ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .b ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_3574, MixColumnsIns_n10}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U6 ( .a ({new_AGEMA_signal_3575, MixColumnsIns_n37}), .b ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3655, MixColumnsIns_n2}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U5 ( .a ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3575, MixColumnsIns_n37}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U4 ( .a ({new_AGEMA_signal_3656, MixColumnsIns_n1}), .b ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3751, MixColumnsOutput[0]}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U3 ( .a ({new_AGEMA_signal_3577, MixColumnsIns_n59}), .b ({new_AGEMA_signal_3576, MixColumnsIns_n23}), .c ({new_AGEMA_signal_3656, MixColumnsIns_n1}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U2 ( .a ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .b ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3576, MixColumnsIns_n23}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_U1 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3577, MixColumnsIns_n59}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_3578, MixColumnsIns_DoubleBytes[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3579, MixColumnsIns_DoubleBytes[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3580, MixColumnsIns_DoubleBytes[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_3581, MixColumnsIns_DoubleBytes[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3582, MixColumnsIns_DoubleBytes[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3583, MixColumnsIns_DoubleBytes[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_3584, MixColumnsIns_DoubleBytes[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3585, MixColumnsIns_DoubleBytes[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3586, MixColumnsIns_DoubleBytes[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .c ({new_AGEMA_signal_3587, MixColumnsIns_DoubleBytes[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .c ({new_AGEMA_signal_3588, MixColumnsIns_DoubleBytes[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) MixColumnsIns_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3589, MixColumnsIns_DoubleBytes[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_0_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3751, MixColumnsOutput[0]}), .a ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3878, ColumnOutput[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_1_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_3873, MixColumnsOutput[1]}), .a ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_4023, ColumnOutput[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_2_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_3729, MixColumnsOutput[2]}), .a ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .c ({new_AGEMA_signal_3879, ColumnOutput[2]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_3_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_3868, MixColumnsOutput[3]}), .a ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .c ({new_AGEMA_signal_4024, ColumnOutput[3]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_4_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_3867, MixColumnsOutput[4]}), .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_4025, ColumnOutput[4]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_5_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_3724, MixColumnsOutput[5]}), .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_3880, ColumnOutput[5]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_6_U1 ( .s (LastRoundorDone), .b ({new_AGEMA_signal_3723, MixColumnsOutput[6]}), .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_3881, ColumnOutput[6]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_7_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3722, MixColumnsOutput[7]}), .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_3882, ColumnOutput[7]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_8_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3721, MixColumnsOutput[8]}), .a ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3883, ColumnOutput[8]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_9_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3866, MixColumnsOutput[9]}), .a ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4026, ColumnOutput[9]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_10_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3750, MixColumnsOutput[10]}), .a ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3884, ColumnOutput[10]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_11_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3877, MixColumnsOutput[11]}), .a ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_4027, ColumnOutput[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_12_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3876, MixColumnsOutput[12]}), .a ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_4028, ColumnOutput[12]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_13_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3747, MixColumnsOutput[13]}), .a ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3885, ColumnOutput[13]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_14_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3746, MixColumnsOutput[14]}), .a ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3886, ColumnOutput[14]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_15_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3745, MixColumnsOutput[15]}), .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_3887, ColumnOutput[15]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_16_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3744, MixColumnsOutput[16]}), .a ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3888, ColumnOutput[16]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_17_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3875, MixColumnsOutput[17]}), .a ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_4029, ColumnOutput[17]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_18_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3742, MixColumnsOutput[18]}), .a ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3889, ColumnOutput[18]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_19_U1 ( .s (MuxMCOut_n5), .b ({new_AGEMA_signal_3874, MixColumnsOutput[19]}), .a ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_4030, ColumnOutput[19]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_20_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3872, MixColumnsOutput[20]}), .a ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_4031, ColumnOutput[20]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_21_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3738, MixColumnsOutput[21]}), .a ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3890, ColumnOutput[21]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_22_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3737, MixColumnsOutput[22]}), .a ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3891, ColumnOutput[22]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_23_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3736, MixColumnsOutput[23]}), .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3892, ColumnOutput[23]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_24_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3735, MixColumnsOutput[24]}), .a ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3893, ColumnOutput[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_25_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3871, MixColumnsOutput[25]}), .a ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_4032, ColumnOutput[25]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_26_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3733, MixColumnsOutput[26]}), .a ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3894, ColumnOutput[26]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_27_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3870, MixColumnsOutput[27]}), .a ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4033, ColumnOutput[27]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_28_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3869, MixColumnsOutput[28]}), .a ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4034, ColumnOutput[28]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_29_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3730, MixColumnsOutput[29]}), .a ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3895, ColumnOutput[29]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_30_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3728, MixColumnsOutput[30]}), .a ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3896, ColumnOutput[30]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxMCOut_mux_inst_31_U1 ( .s (MuxMCOut_n4), .b ({new_AGEMA_signal_3727, MixColumnsOutput[31]}), .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3897, ColumnOutput[31]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_0_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3878, ColumnOutput[0]}), .a ({new_AGEMA_signal_2499, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_4035, RoundOutput[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_1_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_4023, ColumnOutput[1]}), .a ({new_AGEMA_signal_2502, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_4195, RoundOutput[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_2_U1 ( .s (MuxRound_n14), .b ({new_AGEMA_signal_3879, ColumnOutput[2]}), .a ({new_AGEMA_signal_2505, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_4036, RoundOutput[2]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_3_U1 ( .s (MuxRound_n15), .b ({new_AGEMA_signal_4024, ColumnOutput[3]}), .a ({new_AGEMA_signal_2508, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_4196, RoundOutput[3]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_4_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_4025, ColumnOutput[4]}), .a ({new_AGEMA_signal_2511, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_4197, RoundOutput[4]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_5_U1 ( .s (MuxRound_n17), .b ({new_AGEMA_signal_3880, ColumnOutput[5]}), .a ({new_AGEMA_signal_2514, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_4037, RoundOutput[5]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_6_U1 ( .s (MuxRound_n18), .b ({new_AGEMA_signal_3881, ColumnOutput[6]}), .a ({new_AGEMA_signal_2517, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_4038, RoundOutput[6]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_7_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_3882, ColumnOutput[7]}), .a ({new_AGEMA_signal_2520, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_4039, RoundOutput[7]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_8_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_3883, ColumnOutput[8]}), .a ({new_AGEMA_signal_2631, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_4040, RoundOutput[8]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_9_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_4026, ColumnOutput[9]}), .a ({new_AGEMA_signal_2634, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_4198, RoundOutput[9]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_10_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3884, ColumnOutput[10]}), .a ({new_AGEMA_signal_2637, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_4041, RoundOutput[10]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_11_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_4027, ColumnOutput[11]}), .a ({new_AGEMA_signal_2640, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_4199, RoundOutput[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_12_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_4028, ColumnOutput[12]}), .a ({new_AGEMA_signal_2643, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_4200, RoundOutput[12]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_13_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3885, ColumnOutput[13]}), .a ({new_AGEMA_signal_2646, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_4042, RoundOutput[13]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_14_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3886, ColumnOutput[14]}), .a ({new_AGEMA_signal_2649, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_4043, RoundOutput[14]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_15_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3887, ColumnOutput[15]}), .a ({new_AGEMA_signal_2652, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_4044, RoundOutput[15]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_16_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3888, ColumnOutput[16]}), .a ({new_AGEMA_signal_2382, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_4045, RoundOutput[16]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_17_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_4029, ColumnOutput[17]}), .a ({new_AGEMA_signal_2385, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_4201, RoundOutput[17]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_18_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_3889, ColumnOutput[18]}), .a ({new_AGEMA_signal_2388, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_4046, RoundOutput[18]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_19_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_4030, ColumnOutput[19]}), .a ({new_AGEMA_signal_2391, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_4202, RoundOutput[19]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_20_U1 ( .s (MuxRound_n14), .b ({new_AGEMA_signal_4031, ColumnOutput[20]}), .a ({new_AGEMA_signal_2394, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_4203, RoundOutput[20]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_21_U1 ( .s (MuxRound_n15), .b ({new_AGEMA_signal_3890, ColumnOutput[21]}), .a ({new_AGEMA_signal_2397, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_4047, RoundOutput[21]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_22_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_3891, ColumnOutput[22]}), .a ({new_AGEMA_signal_2400, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_4048, RoundOutput[22]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_23_U1 ( .s (MuxRound_n17), .b ({new_AGEMA_signal_3892, ColumnOutput[23]}), .a ({new_AGEMA_signal_2403, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_4049, RoundOutput[23]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_24_U1 ( .s (MuxRound_n18), .b ({new_AGEMA_signal_3893, ColumnOutput[24]}), .a ({new_AGEMA_signal_2472, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_4050, RoundOutput[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_25_U1 ( .s (MuxRound_n16), .b ({new_AGEMA_signal_4032, ColumnOutput[25]}), .a ({new_AGEMA_signal_2475, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_4204, RoundOutput[25]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_26_U1 ( .s (MuxRound_n17), .b ({new_AGEMA_signal_3894, ColumnOutput[26]}), .a ({new_AGEMA_signal_2478, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_4051, RoundOutput[26]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_27_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_4033, ColumnOutput[27]}), .a ({new_AGEMA_signal_2481, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_4205, RoundOutput[27]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_28_U1 ( .s (AKSRnotDone), .b ({new_AGEMA_signal_4034, ColumnOutput[28]}), .a ({new_AGEMA_signal_2484, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_4206, RoundOutput[28]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_29_U1 ( .s (MuxRound_n13), .b ({new_AGEMA_signal_3895, ColumnOutput[29]}), .a ({new_AGEMA_signal_2487, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_4052, RoundOutput[29]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_30_U1 ( .s (MuxRound_n14), .b ({new_AGEMA_signal_3896, ColumnOutput[30]}), .a ({new_AGEMA_signal_2493, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_4053, RoundOutput[30]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxRound_mux_inst_31_U1 ( .s (MuxRound_n15), .b ({new_AGEMA_signal_3897, ColumnOutput[31]}), .a ({new_AGEMA_signal_2496, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_4054, RoundOutput[31]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3991, RoundKeyOutput[0]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_4056, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4126, RoundKeyOutput[1]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_4208, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4127, RoundKeyOutput[2]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_4210, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4128, RoundKeyOutput[3]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_4212, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4129, RoundKeyOutput[4]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_4214, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4130, RoundKeyOutput[5]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_4216, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4131, RoundKeyOutput[6]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_4218, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4132, RoundKeyOutput[7]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_4220, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3992, RoundKeyOutput[8]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_4058, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4133, RoundKeyOutput[9]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_4222, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4134, RoundKeyOutput[10]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_4224, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4135, RoundKeyOutput[11]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_4226, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4136, RoundKeyOutput[12]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_4228, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4137, RoundKeyOutput[13]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_4230, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4138, RoundKeyOutput[14]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_4232, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4139, RoundKeyOutput[15]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_4234, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3993, RoundKeyOutput[16]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_4060, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4140, RoundKeyOutput[17]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_4236, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4141, RoundKeyOutput[18]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_4238, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4142, RoundKeyOutput[19]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_4240, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4143, RoundKeyOutput[20]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_4242, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4144, RoundKeyOutput[21]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_4244, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4145, RoundKeyOutput[22]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_4246, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4146, RoundKeyOutput[23]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_4248, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4147, RoundKeyOutput[24]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_4250, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4265, RoundKeyOutput[25]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_4297, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4266, RoundKeyOutput[26]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_4299, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4267, RoundKeyOutput[27]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_4301, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4268, RoundKeyOutput[28]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_4303, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4269, RoundKeyOutput[29]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_4305, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4270, RoundKeyOutput[30]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_4307, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4271, RoundKeyOutput[31]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_4309, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3834, RoundKeyOutput[32]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_3899, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3994, RoundKeyOutput[33]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_4062, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3995, RoundKeyOutput[34]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_4064, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3996, RoundKeyOutput[35]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_4066, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3997, RoundKeyOutput[36]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_4068, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3998, RoundKeyOutput[37]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_4070, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3999, RoundKeyOutput[38]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_4072, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4000, RoundKeyOutput[39]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_4074, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3835, RoundKeyOutput[40]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_3901, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4001, RoundKeyOutput[41]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_4076, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4002, RoundKeyOutput[42]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_4078, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4003, RoundKeyOutput[43]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_4080, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4004, RoundKeyOutput[44]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_4082, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4005, RoundKeyOutput[45]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_4084, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4006, RoundKeyOutput[46]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_4086, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4007, RoundKeyOutput[47]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_4088, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3836, RoundKeyOutput[48]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_3903, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4008, RoundKeyOutput[49]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_4090, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4009, RoundKeyOutput[50]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_4092, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4010, RoundKeyOutput[51]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_4094, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4011, RoundKeyOutput[52]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_4096, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4012, RoundKeyOutput[53]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_4098, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4013, RoundKeyOutput[54]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_4100, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4014, RoundKeyOutput[55]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_4102, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4015, RoundKeyOutput[56]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_4104, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4148, RoundKeyOutput[57]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_4252, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4149, RoundKeyOutput[58]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_4254, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4150, RoundKeyOutput[59]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_4256, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4151, RoundKeyOutput[60]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_4258, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4152, RoundKeyOutput[61]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_4260, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4153, RoundKeyOutput[62]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_4262, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4154, RoundKeyOutput[63]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_4264, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3695, RoundKeyOutput[64]}), .a ({key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_3753, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3837, RoundKeyOutput[65]}), .a ({key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_3905, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3838, RoundKeyOutput[66]}), .a ({key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_3907, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3839, RoundKeyOutput[67]}), .a ({key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_3909, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3840, RoundKeyOutput[68]}), .a ({key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_3911, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3841, RoundKeyOutput[69]}), .a ({key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_3913, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3842, RoundKeyOutput[70]}), .a ({key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_3915, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3843, RoundKeyOutput[71]}), .a ({key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_3917, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3696, RoundKeyOutput[72]}), .a ({key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_3755, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3844, RoundKeyOutput[73]}), .a ({key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_3919, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3845, RoundKeyOutput[74]}), .a ({key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_3921, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3846, RoundKeyOutput[75]}), .a ({key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_3923, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3847, RoundKeyOutput[76]}), .a ({key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_3925, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3848, RoundKeyOutput[77]}), .a ({key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_3927, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3849, RoundKeyOutput[78]}), .a ({key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_3929, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3850, RoundKeyOutput[79]}), .a ({key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_3931, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3697, RoundKeyOutput[80]}), .a ({key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_3757, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3851, RoundKeyOutput[81]}), .a ({key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_3933, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3852, RoundKeyOutput[82]}), .a ({key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_3935, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3853, RoundKeyOutput[83]}), .a ({key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_3937, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3854, RoundKeyOutput[84]}), .a ({key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_3939, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3855, RoundKeyOutput[85]}), .a ({key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_3941, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3856, RoundKeyOutput[86]}), .a ({key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_3943, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3857, RoundKeyOutput[87]}), .a ({key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_3945, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3858, RoundKeyOutput[88]}), .a ({key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_3947, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4016, RoundKeyOutput[89]}), .a ({key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_4106, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4017, RoundKeyOutput[90]}), .a ({key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_4108, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4018, RoundKeyOutput[91]}), .a ({key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_4110, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4019, RoundKeyOutput[92]}), .a ({key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_4112, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4020, RoundKeyOutput[93]}), .a ({key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_4114, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4021, RoundKeyOutput[94]}), .a ({key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_4116, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_4022, RoundKeyOutput[95]}), .a ({key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_4118, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3622, RoundKeyOutput[96]}), .a ({key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_3658, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3698, RoundKeyOutput[97]}), .a ({key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_3759, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3699, RoundKeyOutput[98]}), .a ({key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_3761, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3700, RoundKeyOutput[99]}), .a ({key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_3763, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3701, RoundKeyOutput[100]}), .a ({key_s1[100], key_s0[100]}), .c ({new_AGEMA_signal_3765, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3702, RoundKeyOutput[101]}), .a ({key_s1[101], key_s0[101]}), .c ({new_AGEMA_signal_3767, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3703, RoundKeyOutput[102]}), .a ({key_s1[102], key_s0[102]}), .c ({new_AGEMA_signal_3769, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3704, RoundKeyOutput[103]}), .a ({key_s1[103], key_s0[103]}), .c ({new_AGEMA_signal_3771, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3623, RoundKeyOutput[104]}), .a ({key_s1[104], key_s0[104]}), .c ({new_AGEMA_signal_3660, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3705, RoundKeyOutput[105]}), .a ({key_s1[105], key_s0[105]}), .c ({new_AGEMA_signal_3773, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3706, RoundKeyOutput[106]}), .a ({key_s1[106], key_s0[106]}), .c ({new_AGEMA_signal_3775, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3707, RoundKeyOutput[107]}), .a ({key_s1[107], key_s0[107]}), .c ({new_AGEMA_signal_3777, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3708, RoundKeyOutput[108]}), .a ({key_s1[108], key_s0[108]}), .c ({new_AGEMA_signal_3779, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3709, RoundKeyOutput[109]}), .a ({key_s1[109], key_s0[109]}), .c ({new_AGEMA_signal_3781, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3710, RoundKeyOutput[110]}), .a ({key_s1[110], key_s0[110]}), .c ({new_AGEMA_signal_3783, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3711, RoundKeyOutput[111]}), .a ({key_s1[111], key_s0[111]}), .c ({new_AGEMA_signal_3785, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3624, RoundKeyOutput[112]}), .a ({key_s1[112], key_s0[112]}), .c ({new_AGEMA_signal_3662, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3712, RoundKeyOutput[113]}), .a ({key_s1[113], key_s0[113]}), .c ({new_AGEMA_signal_3787, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3713, RoundKeyOutput[114]}), .a ({key_s1[114], key_s0[114]}), .c ({new_AGEMA_signal_3789, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3714, RoundKeyOutput[115]}), .a ({key_s1[115], key_s0[115]}), .c ({new_AGEMA_signal_3791, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3715, RoundKeyOutput[116]}), .a ({key_s1[116], key_s0[116]}), .c ({new_AGEMA_signal_3793, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3716, RoundKeyOutput[117]}), .a ({key_s1[117], key_s0[117]}), .c ({new_AGEMA_signal_3795, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3717, RoundKeyOutput[118]}), .a ({key_s1[118], key_s0[118]}), .c ({new_AGEMA_signal_3797, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3718, RoundKeyOutput[119]}), .a ({key_s1[119], key_s0[119]}), .c ({new_AGEMA_signal_3799, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3719, RoundKeyOutput[120]}), .a ({key_s1[120], key_s0[120]}), .c ({new_AGEMA_signal_3801, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3859, RoundKeyOutput[121]}), .a ({key_s1[121], key_s0[121]}), .c ({new_AGEMA_signal_3949, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3860, RoundKeyOutput[122]}), .a ({key_s1[122], key_s0[122]}), .c ({new_AGEMA_signal_3951, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3861, RoundKeyOutput[123]}), .a ({key_s1[123], key_s0[123]}), .c ({new_AGEMA_signal_3953, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3862, RoundKeyOutput[124]}), .a ({key_s1[124], key_s0[124]}), .c ({new_AGEMA_signal_3955, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3863, RoundKeyOutput[125]}), .a ({key_s1[125], key_s0[125]}), .c ({new_AGEMA_signal_3957, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3864, RoundKeyOutput[126]}), .a ({key_s1[126], key_s0[126]}), .c ({new_AGEMA_signal_3959, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_3865, RoundKeyOutput[127]}), .a ({key_s1[127], key_s0[127]}), .c ({new_AGEMA_signal_3961, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_2720, KSSubBytesInput[9]}), .b ({new_AGEMA_signal_3803, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_3962, KeyExpansionOutput[9]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_2687, KSSubBytesInput[8]}), .b ({new_AGEMA_signal_3664, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_3802, KeyExpansionOutput[8]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_2654, KSSubBytesInput[23]}), .b ({new_AGEMA_signal_3804, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_3963, KeyExpansionOutput[7]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_2621, KSSubBytesInput[22]}), .b ({new_AGEMA_signal_3805, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_3964, KeyExpansionOutput[6]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_2588, KSSubBytesInput[21]}), .b ({new_AGEMA_signal_3806, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_3965, KeyExpansionOutput[5]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_2555, KSSubBytesInput[20]}), .b ({new_AGEMA_signal_3807, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_3966, KeyExpansionOutput[4]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_2528, RoundKey[41]}), .b ({new_AGEMA_signal_3663, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_3803, KeyExpansionOutput[41]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_2633, RoundKey[73]}), .b ({new_AGEMA_signal_3609, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_3663, KeyExpansionOutput[73]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_2525, RoundKey[40]}), .b ({new_AGEMA_signal_3590, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_3664, KeyExpansionOutput[40]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_2630, RoundKey[72]}), .b ({new_AGEMA_signal_3555, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_3590, KeyExpansionOutput[72]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_2522, KSSubBytesInput[19]}), .b ({new_AGEMA_signal_3808, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_3967, KeyExpansionOutput[3]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_2519, RoundKey[39]}), .b ({new_AGEMA_signal_3665, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_3804, KeyExpansionOutput[39]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_2627, RoundKey[71]}), .b ({new_AGEMA_signal_3610, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_3665, KeyExpansionOutput[71]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_2516, RoundKey[38]}), .b ({new_AGEMA_signal_3666, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_3805, KeyExpansionOutput[38]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_2624, RoundKey[70]}), .b ({new_AGEMA_signal_3611, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_3666, KeyExpansionOutput[70]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_2513, RoundKey[37]}), .b ({new_AGEMA_signal_3667, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_3806, KeyExpansionOutput[37]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_2618, RoundKey[69]}), .b ({new_AGEMA_signal_3612, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_3667, KeyExpansionOutput[69]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_2510, RoundKey[36]}), .b ({new_AGEMA_signal_3668, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_3807, KeyExpansionOutput[36]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_2615, RoundKey[68]}), .b ({new_AGEMA_signal_3613, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_3668, KeyExpansionOutput[68]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_2507, RoundKey[35]}), .b ({new_AGEMA_signal_3669, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_3808, KeyExpansionOutput[35]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_2612, RoundKey[67]}), .b ({new_AGEMA_signal_3591, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_3669, KeyExpansionOutput[67]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_2717, RoundKey[99]}), .b ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_3591, KeyExpansionOutput[99]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_2495, KSSubBytesInput[31]}), .b ({new_AGEMA_signal_3968, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_4119, KeyExpansionOutput[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_2600, RoundKey[63]}), .b ({new_AGEMA_signal_3809, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_3968, KeyExpansionOutput[63]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_2705, RoundKey[95]}), .b ({new_AGEMA_signal_3685, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_3809, KeyExpansionOutput[95]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_2492, KSSubBytesInput[30]}), .b ({new_AGEMA_signal_3969, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_4120, KeyExpansionOutput[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_2597, RoundKey[62]}), .b ({new_AGEMA_signal_3810, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_3969, KeyExpansionOutput[62]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_2702, RoundKey[94]}), .b ({new_AGEMA_signal_3686, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_3810, KeyExpansionOutput[94]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_2489, KSSubBytesInput[18]}), .b ({new_AGEMA_signal_3811, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_3970, KeyExpansionOutput[2]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_2504, RoundKey[34]}), .b ({new_AGEMA_signal_3670, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_3811, KeyExpansionOutput[34]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_2609, RoundKey[66]}), .b ({new_AGEMA_signal_3592, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_3670, KeyExpansionOutput[66]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_2714, RoundKey[98]}), .b ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3592, KeyExpansionOutput[98]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_2486, KSSubBytesInput[29]}), .b ({new_AGEMA_signal_3971, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_4121, KeyExpansionOutput[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_2594, RoundKey[61]}), .b ({new_AGEMA_signal_3812, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_3971, KeyExpansionOutput[61]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_2699, RoundKey[93]}), .b ({new_AGEMA_signal_3687, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_3812, KeyExpansionOutput[93]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_2483, KSSubBytesInput[28]}), .b ({new_AGEMA_signal_3972, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_4122, KeyExpansionOutput[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_2591, RoundKey[60]}), .b ({new_AGEMA_signal_3813, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_3972, KeyExpansionOutput[60]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_2696, RoundKey[92]}), .b ({new_AGEMA_signal_3688, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_3813, KeyExpansionOutput[92]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_2480, KSSubBytesInput[27]}), .b ({new_AGEMA_signal_3973, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_4123, KeyExpansionOutput[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_2585, RoundKey[59]}), .b ({new_AGEMA_signal_3814, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_3973, KeyExpansionOutput[59]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_2693, RoundKey[91]}), .b ({new_AGEMA_signal_3689, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_3814, KeyExpansionOutput[91]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_2477, KSSubBytesInput[26]}), .b ({new_AGEMA_signal_3974, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_4124, KeyExpansionOutput[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_2582, RoundKey[58]}), .b ({new_AGEMA_signal_3815, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_3974, KeyExpansionOutput[58]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_2690, RoundKey[90]}), .b ({new_AGEMA_signal_3690, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_3815, KeyExpansionOutput[90]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_2474, KSSubBytesInput[25]}), .b ({new_AGEMA_signal_3975, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_4125, KeyExpansionOutput[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_2579, RoundKey[57]}), .b ({new_AGEMA_signal_3816, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_3975, KeyExpansionOutput[57]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_2684, RoundKey[89]}), .b ({new_AGEMA_signal_3691, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_3816, KeyExpansionOutput[89]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_2471, KSSubBytesInput[24]}), .b ({new_AGEMA_signal_3817, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_3976, KeyExpansionOutput[24]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_2576, RoundKey[56]}), .b ({new_AGEMA_signal_3671, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_3817, KeyExpansionOutput[56]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_2681, RoundKey[88]}), .b ({new_AGEMA_signal_3595, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_3671, KeyExpansionOutput[88]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_2468, KSSubBytesInput[7]}), .b ({new_AGEMA_signal_3818, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_3977, KeyExpansionOutput[23]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_2573, RoundKey[55]}), .b ({new_AGEMA_signal_3672, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_3818, KeyExpansionOutput[55]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_2678, RoundKey[87]}), .b ({new_AGEMA_signal_3596, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_3672, KeyExpansionOutput[87]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_2465, KSSubBytesInput[6]}), .b ({new_AGEMA_signal_3819, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_3978, KeyExpansionOutput[22]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_2570, RoundKey[54]}), .b ({new_AGEMA_signal_3673, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_3819, KeyExpansionOutput[54]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_2675, RoundKey[86]}), .b ({new_AGEMA_signal_3597, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_3673, KeyExpansionOutput[86]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_2462, KSSubBytesInput[5]}), .b ({new_AGEMA_signal_3820, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_3979, KeyExpansionOutput[21]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_2567, RoundKey[53]}), .b ({new_AGEMA_signal_3674, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_3820, KeyExpansionOutput[53]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_2672, RoundKey[85]}), .b ({new_AGEMA_signal_3598, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_3674, KeyExpansionOutput[85]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_2459, KSSubBytesInput[4]}), .b ({new_AGEMA_signal_3821, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_3980, KeyExpansionOutput[20]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_2564, RoundKey[52]}), .b ({new_AGEMA_signal_3675, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_3821, KeyExpansionOutput[52]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_2669, RoundKey[84]}), .b ({new_AGEMA_signal_3599, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_3675, KeyExpansionOutput[84]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_2456, KSSubBytesInput[17]}), .b ({new_AGEMA_signal_3822, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_3981, KeyExpansionOutput[1]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_2501, RoundKey[33]}), .b ({new_AGEMA_signal_3676, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_3822, KeyExpansionOutput[33]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_2606, RoundKey[65]}), .b ({new_AGEMA_signal_3593, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_3676, KeyExpansionOutput[65]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_2711, RoundKey[97]}), .b ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_3593, KeyExpansionOutput[97]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_2453, KSSubBytesInput[3]}), .b ({new_AGEMA_signal_3823, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_3982, KeyExpansionOutput[19]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_2561, RoundKey[51]}), .b ({new_AGEMA_signal_3677, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_3823, KeyExpansionOutput[51]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_2666, RoundKey[83]}), .b ({new_AGEMA_signal_3600, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_3677, KeyExpansionOutput[83]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_2450, KSSubBytesInput[2]}), .b ({new_AGEMA_signal_3824, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_3983, KeyExpansionOutput[18]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_2558, RoundKey[50]}), .b ({new_AGEMA_signal_3678, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_3824, KeyExpansionOutput[50]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_2663, RoundKey[82]}), .b ({new_AGEMA_signal_3601, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_3678, KeyExpansionOutput[82]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_2447, KSSubBytesInput[1]}), .b ({new_AGEMA_signal_3825, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_3984, KeyExpansionOutput[17]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_2552, RoundKey[49]}), .b ({new_AGEMA_signal_3679, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_3825, KeyExpansionOutput[49]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_2660, RoundKey[81]}), .b ({new_AGEMA_signal_3602, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_3679, KeyExpansionOutput[81]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_2444, KSSubBytesInput[0]}), .b ({new_AGEMA_signal_3680, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_3826, KeyExpansionOutput[16]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_2549, RoundKey[48]}), .b ({new_AGEMA_signal_3594, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_3680, KeyExpansionOutput[48]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_2657, RoundKey[80]}), .b ({new_AGEMA_signal_3554, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_3594, KeyExpansionOutput[80]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_2441, KSSubBytesInput[15]}), .b ({new_AGEMA_signal_3827, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_3985, KeyExpansionOutput[15]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_2546, RoundKey[47]}), .b ({new_AGEMA_signal_3681, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_3827, KeyExpansionOutput[47]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_2651, RoundKey[79]}), .b ({new_AGEMA_signal_3603, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_3681, KeyExpansionOutput[79]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_2438, KSSubBytesInput[14]}), .b ({new_AGEMA_signal_3828, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_3986, KeyExpansionOutput[14]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_2543, RoundKey[46]}), .b ({new_AGEMA_signal_3682, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_3828, KeyExpansionOutput[46]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_2648, RoundKey[78]}), .b ({new_AGEMA_signal_3604, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_3682, KeyExpansionOutput[78]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_2435, KSSubBytesInput[13]}), .b ({new_AGEMA_signal_3829, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_3987, KeyExpansionOutput[13]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_2540, RoundKey[45]}), .b ({new_AGEMA_signal_3683, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_3829, KeyExpansionOutput[45]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_2645, RoundKey[77]}), .b ({new_AGEMA_signal_3605, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_3683, KeyExpansionOutput[77]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_2432, KSSubBytesInput[12]}), .b ({new_AGEMA_signal_3830, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_3988, KeyExpansionOutput[12]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_2537, RoundKey[44]}), .b ({new_AGEMA_signal_3684, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_3830, KeyExpansionOutput[44]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_2642, RoundKey[76]}), .b ({new_AGEMA_signal_3606, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_3684, KeyExpansionOutput[76]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_2429, RoundKey[127]}), .b ({new_AGEMA_signal_3615, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_3685, KeyExpansionOutput[127]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_2426, RoundKey[126]}), .b ({new_AGEMA_signal_3616, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_3686, KeyExpansionOutput[126]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_2423, RoundKey[125]}), .b ({new_AGEMA_signal_3617, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_3687, KeyExpansionOutput[125]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_2420, RoundKey[124]}), .b ({new_AGEMA_signal_3618, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_3688, KeyExpansionOutput[124]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_2417, RoundKey[123]}), .b ({new_AGEMA_signal_3619, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_3689, KeyExpansionOutput[123]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_2414, RoundKey[122]}), .b ({new_AGEMA_signal_3620, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_3690, KeyExpansionOutput[122]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_2411, RoundKey[121]}), .b ({new_AGEMA_signal_3621, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_3691, KeyExpansionOutput[121]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_2408, RoundKey[120]}), .b ({new_AGEMA_signal_3557, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_3595, KeyExpansionOutput[120]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_2405, KSSubBytesInput[11]}), .b ({new_AGEMA_signal_3831, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_3989, KeyExpansionOutput[11]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_2534, RoundKey[43]}), .b ({new_AGEMA_signal_3692, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_3831, KeyExpansionOutput[43]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_2639, RoundKey[75]}), .b ({new_AGEMA_signal_3607, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_3692, KeyExpansionOutput[75]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_2402, RoundKey[119]}), .b ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_3596, KeyExpansionOutput[119]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_2399, RoundKey[118]}), .b ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3597, KeyExpansionOutput[118]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_2396, RoundKey[117]}), .b ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3598, KeyExpansionOutput[117]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_2393, RoundKey[116]}), .b ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_3599, KeyExpansionOutput[116]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_2390, RoundKey[115]}), .b ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_3600, KeyExpansionOutput[115]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_2387, RoundKey[114]}), .b ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3601, KeyExpansionOutput[114]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_2384, RoundKey[113]}), .b ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_3602, KeyExpansionOutput[113]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_2381, RoundKey[112]}), .b ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3554, KeyExpansionOutput[112]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_2378, RoundKey[111]}), .b ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3603, KeyExpansionOutput[111]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_2375, RoundKey[110]}), .b ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3604, KeyExpansionOutput[110]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_2372, KSSubBytesInput[10]}), .b ({new_AGEMA_signal_3832, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_3990, KeyExpansionOutput[10]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_2531, RoundKey[42]}), .b ({new_AGEMA_signal_3693, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_3832, KeyExpansionOutput[42]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_2636, RoundKey[74]}), .b ({new_AGEMA_signal_3608, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_3693, KeyExpansionOutput[74]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_2369, RoundKey[109]}), .b ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3605, KeyExpansionOutput[109]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_2366, RoundKey[108]}), .b ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_3606, KeyExpansionOutput[108]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_2363, RoundKey[107]}), .b ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_3607, KeyExpansionOutput[107]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_2360, RoundKey[106]}), .b ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3608, KeyExpansionOutput[106]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_2357, RoundKey[105]}), .b ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_3609, KeyExpansionOutput[105]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_2354, RoundKey[104]}), .b ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3555, KeyExpansionOutput[104]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_2351, RoundKey[103]}), .b ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3610, KeyExpansionOutput[103]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_2348, RoundKey[102]}), .b ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3611, KeyExpansionOutput[102]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_2345, RoundKey[101]}), .b ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3612, KeyExpansionOutput[101]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_2342, RoundKey[100]}), .b ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_3613, KeyExpansionOutput[100]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_2339, KSSubBytesInput[16]}), .b ({new_AGEMA_signal_3694, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_3833, KeyExpansionOutput[0]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_2498, RoundKey[32]}), .b ({new_AGEMA_signal_3614, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_3694, KeyExpansionOutput[32]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_2603, RoundKey[64]}), .b ({new_AGEMA_signal_3556, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_3614, KeyExpansionOutput[64]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_2708, RoundKey[96]}), .b ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3556, KeyExpansionOutput[96]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({1'b0, Rcon[7]}), .b ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_3615, KeyExpansionIns_tmp[31]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({1'b0, Rcon[6]}), .b ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_3616, KeyExpansionIns_tmp[30]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({1'b0, Rcon[5]}), .b ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_3617, KeyExpansionIns_tmp[29]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({1'b0, Rcon[4]}), .b ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_3618, KeyExpansionIns_tmp[28]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({1'b0, Rcon[3]}), .b ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .c ({new_AGEMA_signal_3619, KeyExpansionIns_tmp[27]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({1'b0, Rcon[2]}), .b ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .c ({new_AGEMA_signal_3620, KeyExpansionIns_tmp[26]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({1'b0, Rcon[1]}), .b ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_3621, KeyExpansionIns_tmp[25]}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({1'b0, Rcon[0]}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3557, KeyExpansionIns_tmp[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_0_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2339, KSSubBytesInput[16]}), .a ({new_AGEMA_signal_3833, KeyExpansionOutput[0]}), .c ({new_AGEMA_signal_3991, RoundKeyOutput[0]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_1_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2456, KSSubBytesInput[17]}), .a ({new_AGEMA_signal_3981, KeyExpansionOutput[1]}), .c ({new_AGEMA_signal_4126, RoundKeyOutput[1]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_2_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2489, KSSubBytesInput[18]}), .a ({new_AGEMA_signal_3970, KeyExpansionOutput[2]}), .c ({new_AGEMA_signal_4127, RoundKeyOutput[2]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_3_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2522, KSSubBytesInput[19]}), .a ({new_AGEMA_signal_3967, KeyExpansionOutput[3]}), .c ({new_AGEMA_signal_4128, RoundKeyOutput[3]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_4_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2555, KSSubBytesInput[20]}), .a ({new_AGEMA_signal_3966, KeyExpansionOutput[4]}), .c ({new_AGEMA_signal_4129, RoundKeyOutput[4]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_5_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2588, KSSubBytesInput[21]}), .a ({new_AGEMA_signal_3965, KeyExpansionOutput[5]}), .c ({new_AGEMA_signal_4130, RoundKeyOutput[5]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_6_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2621, KSSubBytesInput[22]}), .a ({new_AGEMA_signal_3964, KeyExpansionOutput[6]}), .c ({new_AGEMA_signal_4131, RoundKeyOutput[6]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_7_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2654, KSSubBytesInput[23]}), .a ({new_AGEMA_signal_3963, KeyExpansionOutput[7]}), .c ({new_AGEMA_signal_4132, RoundKeyOutput[7]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_8_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2687, KSSubBytesInput[8]}), .a ({new_AGEMA_signal_3802, KeyExpansionOutput[8]}), .c ({new_AGEMA_signal_3992, RoundKeyOutput[8]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_9_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2720, KSSubBytesInput[9]}), .a ({new_AGEMA_signal_3962, KeyExpansionOutput[9]}), .c ({new_AGEMA_signal_4133, RoundKeyOutput[9]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_10_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2372, KSSubBytesInput[10]}), .a ({new_AGEMA_signal_3990, KeyExpansionOutput[10]}), .c ({new_AGEMA_signal_4134, RoundKeyOutput[10]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_11_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2405, KSSubBytesInput[11]}), .a ({new_AGEMA_signal_3989, KeyExpansionOutput[11]}), .c ({new_AGEMA_signal_4135, RoundKeyOutput[11]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_12_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2432, KSSubBytesInput[12]}), .a ({new_AGEMA_signal_3988, KeyExpansionOutput[12]}), .c ({new_AGEMA_signal_4136, RoundKeyOutput[12]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_13_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2435, KSSubBytesInput[13]}), .a ({new_AGEMA_signal_3987, KeyExpansionOutput[13]}), .c ({new_AGEMA_signal_4137, RoundKeyOutput[13]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_14_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2438, KSSubBytesInput[14]}), .a ({new_AGEMA_signal_3986, KeyExpansionOutput[14]}), .c ({new_AGEMA_signal_4138, RoundKeyOutput[14]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_15_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2441, KSSubBytesInput[15]}), .a ({new_AGEMA_signal_3985, KeyExpansionOutput[15]}), .c ({new_AGEMA_signal_4139, RoundKeyOutput[15]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_16_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2444, KSSubBytesInput[0]}), .a ({new_AGEMA_signal_3826, KeyExpansionOutput[16]}), .c ({new_AGEMA_signal_3993, RoundKeyOutput[16]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_17_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2447, KSSubBytesInput[1]}), .a ({new_AGEMA_signal_3984, KeyExpansionOutput[17]}), .c ({new_AGEMA_signal_4140, RoundKeyOutput[17]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_18_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2450, KSSubBytesInput[2]}), .a ({new_AGEMA_signal_3983, KeyExpansionOutput[18]}), .c ({new_AGEMA_signal_4141, RoundKeyOutput[18]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_19_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2453, KSSubBytesInput[3]}), .a ({new_AGEMA_signal_3982, KeyExpansionOutput[19]}), .c ({new_AGEMA_signal_4142, RoundKeyOutput[19]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_20_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2459, KSSubBytesInput[4]}), .a ({new_AGEMA_signal_3980, KeyExpansionOutput[20]}), .c ({new_AGEMA_signal_4143, RoundKeyOutput[20]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_21_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2462, KSSubBytesInput[5]}), .a ({new_AGEMA_signal_3979, KeyExpansionOutput[21]}), .c ({new_AGEMA_signal_4144, RoundKeyOutput[21]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_22_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2465, KSSubBytesInput[6]}), .a ({new_AGEMA_signal_3978, KeyExpansionOutput[22]}), .c ({new_AGEMA_signal_4145, RoundKeyOutput[22]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_23_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2468, KSSubBytesInput[7]}), .a ({new_AGEMA_signal_3977, KeyExpansionOutput[23]}), .c ({new_AGEMA_signal_4146, RoundKeyOutput[23]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_24_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2471, KSSubBytesInput[24]}), .a ({new_AGEMA_signal_3976, KeyExpansionOutput[24]}), .c ({new_AGEMA_signal_4147, RoundKeyOutput[24]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_25_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2474, KSSubBytesInput[25]}), .a ({new_AGEMA_signal_4125, KeyExpansionOutput[25]}), .c ({new_AGEMA_signal_4265, RoundKeyOutput[25]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_26_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2477, KSSubBytesInput[26]}), .a ({new_AGEMA_signal_4124, KeyExpansionOutput[26]}), .c ({new_AGEMA_signal_4266, RoundKeyOutput[26]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_27_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2480, KSSubBytesInput[27]}), .a ({new_AGEMA_signal_4123, KeyExpansionOutput[27]}), .c ({new_AGEMA_signal_4267, RoundKeyOutput[27]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_28_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2483, KSSubBytesInput[28]}), .a ({new_AGEMA_signal_4122, KeyExpansionOutput[28]}), .c ({new_AGEMA_signal_4268, RoundKeyOutput[28]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_29_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2486, KSSubBytesInput[29]}), .a ({new_AGEMA_signal_4121, KeyExpansionOutput[29]}), .c ({new_AGEMA_signal_4269, RoundKeyOutput[29]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_30_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2492, KSSubBytesInput[30]}), .a ({new_AGEMA_signal_4120, KeyExpansionOutput[30]}), .c ({new_AGEMA_signal_4270, RoundKeyOutput[30]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_31_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2495, KSSubBytesInput[31]}), .a ({new_AGEMA_signal_4119, KeyExpansionOutput[31]}), .c ({new_AGEMA_signal_4271, RoundKeyOutput[31]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_32_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2498, RoundKey[32]}), .a ({new_AGEMA_signal_3694, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_3834, RoundKeyOutput[32]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_33_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2501, RoundKey[33]}), .a ({new_AGEMA_signal_3822, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_3994, RoundKeyOutput[33]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_34_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2504, RoundKey[34]}), .a ({new_AGEMA_signal_3811, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_3995, RoundKeyOutput[34]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_35_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2507, RoundKey[35]}), .a ({new_AGEMA_signal_3808, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_3996, RoundKeyOutput[35]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_36_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2510, RoundKey[36]}), .a ({new_AGEMA_signal_3807, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_3997, RoundKeyOutput[36]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_37_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2513, RoundKey[37]}), .a ({new_AGEMA_signal_3806, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_3998, RoundKeyOutput[37]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_38_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2516, RoundKey[38]}), .a ({new_AGEMA_signal_3805, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_3999, RoundKeyOutput[38]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_39_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2519, RoundKey[39]}), .a ({new_AGEMA_signal_3804, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_4000, RoundKeyOutput[39]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_40_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2525, RoundKey[40]}), .a ({new_AGEMA_signal_3664, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_3835, RoundKeyOutput[40]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_41_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2528, RoundKey[41]}), .a ({new_AGEMA_signal_3803, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_4001, RoundKeyOutput[41]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_42_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2531, RoundKey[42]}), .a ({new_AGEMA_signal_3832, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_4002, RoundKeyOutput[42]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_43_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2534, RoundKey[43]}), .a ({new_AGEMA_signal_3831, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_4003, RoundKeyOutput[43]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_44_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2537, RoundKey[44]}), .a ({new_AGEMA_signal_3830, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_4004, RoundKeyOutput[44]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_45_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2540, RoundKey[45]}), .a ({new_AGEMA_signal_3829, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_4005, RoundKeyOutput[45]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_46_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2543, RoundKey[46]}), .a ({new_AGEMA_signal_3828, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_4006, RoundKeyOutput[46]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_47_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2546, RoundKey[47]}), .a ({new_AGEMA_signal_3827, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_4007, RoundKeyOutput[47]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_48_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2549, RoundKey[48]}), .a ({new_AGEMA_signal_3680, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_3836, RoundKeyOutput[48]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_49_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2552, RoundKey[49]}), .a ({new_AGEMA_signal_3825, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_4008, RoundKeyOutput[49]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_50_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2558, RoundKey[50]}), .a ({new_AGEMA_signal_3824, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_4009, RoundKeyOutput[50]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_51_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2561, RoundKey[51]}), .a ({new_AGEMA_signal_3823, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_4010, RoundKeyOutput[51]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_52_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2564, RoundKey[52]}), .a ({new_AGEMA_signal_3821, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_4011, RoundKeyOutput[52]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_53_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2567, RoundKey[53]}), .a ({new_AGEMA_signal_3820, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_4012, RoundKeyOutput[53]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_54_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2570, RoundKey[54]}), .a ({new_AGEMA_signal_3819, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_4013, RoundKeyOutput[54]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_55_U1 ( .s (MuxKeyExpansion_n20), .b ({new_AGEMA_signal_2573, RoundKey[55]}), .a ({new_AGEMA_signal_3818, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_4014, RoundKeyOutput[55]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_56_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2576, RoundKey[56]}), .a ({new_AGEMA_signal_3817, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_4015, RoundKeyOutput[56]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_57_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2579, RoundKey[57]}), .a ({new_AGEMA_signal_3975, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_4148, RoundKeyOutput[57]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_58_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2582, RoundKey[58]}), .a ({new_AGEMA_signal_3974, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_4149, RoundKeyOutput[58]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_59_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2585, RoundKey[59]}), .a ({new_AGEMA_signal_3973, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_4150, RoundKeyOutput[59]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_60_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2591, RoundKey[60]}), .a ({new_AGEMA_signal_3972, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_4151, RoundKeyOutput[60]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_61_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2594, RoundKey[61]}), .a ({new_AGEMA_signal_3971, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_4152, RoundKeyOutput[61]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_62_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2597, RoundKey[62]}), .a ({new_AGEMA_signal_3969, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_4153, RoundKeyOutput[62]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_63_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2600, RoundKey[63]}), .a ({new_AGEMA_signal_3968, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_4154, RoundKeyOutput[63]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_64_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2603, RoundKey[64]}), .a ({new_AGEMA_signal_3614, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_3695, RoundKeyOutput[64]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_65_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2606, RoundKey[65]}), .a ({new_AGEMA_signal_3676, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_3837, RoundKeyOutput[65]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_66_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2609, RoundKey[66]}), .a ({new_AGEMA_signal_3670, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_3838, RoundKeyOutput[66]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_67_U1 ( .s (MuxKeyExpansion_n19), .b ({new_AGEMA_signal_2612, RoundKey[67]}), .a ({new_AGEMA_signal_3669, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_3839, RoundKeyOutput[67]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_68_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2615, RoundKey[68]}), .a ({new_AGEMA_signal_3668, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_3840, RoundKeyOutput[68]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_69_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2618, RoundKey[69]}), .a ({new_AGEMA_signal_3667, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_3841, RoundKeyOutput[69]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_70_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2624, RoundKey[70]}), .a ({new_AGEMA_signal_3666, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_3842, RoundKeyOutput[70]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_71_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2627, RoundKey[71]}), .a ({new_AGEMA_signal_3665, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_3843, RoundKeyOutput[71]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_72_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2630, RoundKey[72]}), .a ({new_AGEMA_signal_3590, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_3696, RoundKeyOutput[72]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_73_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2633, RoundKey[73]}), .a ({new_AGEMA_signal_3663, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_3844, RoundKeyOutput[73]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_74_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2636, RoundKey[74]}), .a ({new_AGEMA_signal_3693, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_3845, RoundKeyOutput[74]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_75_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2639, RoundKey[75]}), .a ({new_AGEMA_signal_3692, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_3846, RoundKeyOutput[75]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_76_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2642, RoundKey[76]}), .a ({new_AGEMA_signal_3684, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_3847, RoundKeyOutput[76]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_77_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2645, RoundKey[77]}), .a ({new_AGEMA_signal_3683, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_3848, RoundKeyOutput[77]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_78_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2648, RoundKey[78]}), .a ({new_AGEMA_signal_3682, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_3849, RoundKeyOutput[78]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_79_U1 ( .s (MuxKeyExpansion_n18), .b ({new_AGEMA_signal_2651, RoundKey[79]}), .a ({new_AGEMA_signal_3681, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_3850, RoundKeyOutput[79]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_80_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2657, RoundKey[80]}), .a ({new_AGEMA_signal_3594, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_3697, RoundKeyOutput[80]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_81_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2660, RoundKey[81]}), .a ({new_AGEMA_signal_3679, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_3851, RoundKeyOutput[81]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_82_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2663, RoundKey[82]}), .a ({new_AGEMA_signal_3678, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_3852, RoundKeyOutput[82]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_83_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2666, RoundKey[83]}), .a ({new_AGEMA_signal_3677, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_3853, RoundKeyOutput[83]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_84_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2669, RoundKey[84]}), .a ({new_AGEMA_signal_3675, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_3854, RoundKeyOutput[84]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_85_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2672, RoundKey[85]}), .a ({new_AGEMA_signal_3674, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_3855, RoundKeyOutput[85]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_86_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2675, RoundKey[86]}), .a ({new_AGEMA_signal_3673, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_3856, RoundKeyOutput[86]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_87_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2678, RoundKey[87]}), .a ({new_AGEMA_signal_3672, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_3857, RoundKeyOutput[87]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_88_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2681, RoundKey[88]}), .a ({new_AGEMA_signal_3671, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_3858, RoundKeyOutput[88]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_89_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2684, RoundKey[89]}), .a ({new_AGEMA_signal_3816, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_4016, RoundKeyOutput[89]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_90_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2690, RoundKey[90]}), .a ({new_AGEMA_signal_3815, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_4017, RoundKeyOutput[90]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_91_U1 ( .s (MuxKeyExpansion_n17), .b ({new_AGEMA_signal_2693, RoundKey[91]}), .a ({new_AGEMA_signal_3814, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_4018, RoundKeyOutput[91]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_92_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2696, RoundKey[92]}), .a ({new_AGEMA_signal_3813, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_4019, RoundKeyOutput[92]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_93_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2699, RoundKey[93]}), .a ({new_AGEMA_signal_3812, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_4020, RoundKeyOutput[93]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_94_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2702, RoundKey[94]}), .a ({new_AGEMA_signal_3810, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_4021, RoundKeyOutput[94]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_95_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2705, RoundKey[95]}), .a ({new_AGEMA_signal_3809, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_4022, RoundKeyOutput[95]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_96_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2708, RoundKey[96]}), .a ({new_AGEMA_signal_3556, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_3622, RoundKeyOutput[96]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_97_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2711, RoundKey[97]}), .a ({new_AGEMA_signal_3593, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_3698, RoundKeyOutput[97]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_98_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2714, RoundKey[98]}), .a ({new_AGEMA_signal_3592, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_3699, RoundKeyOutput[98]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_99_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2717, RoundKey[99]}), .a ({new_AGEMA_signal_3591, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_3700, RoundKeyOutput[99]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_100_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2342, RoundKey[100]}), .a ({new_AGEMA_signal_3613, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_3701, RoundKeyOutput[100]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_101_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2345, RoundKey[101]}), .a ({new_AGEMA_signal_3612, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_3702, RoundKeyOutput[101]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_102_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2348, RoundKey[102]}), .a ({new_AGEMA_signal_3611, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_3703, RoundKeyOutput[102]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_103_U1 ( .s (MuxKeyExpansion_n16), .b ({new_AGEMA_signal_2351, RoundKey[103]}), .a ({new_AGEMA_signal_3610, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_3704, RoundKeyOutput[103]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_104_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2354, RoundKey[104]}), .a ({new_AGEMA_signal_3555, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_3623, RoundKeyOutput[104]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_105_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2357, RoundKey[105]}), .a ({new_AGEMA_signal_3609, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_3705, RoundKeyOutput[105]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_106_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2360, RoundKey[106]}), .a ({new_AGEMA_signal_3608, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_3706, RoundKeyOutput[106]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_107_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2363, RoundKey[107]}), .a ({new_AGEMA_signal_3607, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_3707, RoundKeyOutput[107]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_108_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2366, RoundKey[108]}), .a ({new_AGEMA_signal_3606, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_3708, RoundKeyOutput[108]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_109_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2369, RoundKey[109]}), .a ({new_AGEMA_signal_3605, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_3709, RoundKeyOutput[109]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_110_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2375, RoundKey[110]}), .a ({new_AGEMA_signal_3604, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_3710, RoundKeyOutput[110]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_111_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2378, RoundKey[111]}), .a ({new_AGEMA_signal_3603, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_3711, RoundKeyOutput[111]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_112_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2381, RoundKey[112]}), .a ({new_AGEMA_signal_3554, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_3624, RoundKeyOutput[112]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_113_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2384, RoundKey[113]}), .a ({new_AGEMA_signal_3602, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_3712, RoundKeyOutput[113]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_114_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2387, RoundKey[114]}), .a ({new_AGEMA_signal_3601, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_3713, RoundKeyOutput[114]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_115_U1 ( .s (MuxKeyExpansion_n15), .b ({new_AGEMA_signal_2390, RoundKey[115]}), .a ({new_AGEMA_signal_3600, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_3714, RoundKeyOutput[115]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_116_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2393, RoundKey[116]}), .a ({new_AGEMA_signal_3599, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_3715, RoundKeyOutput[116]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_117_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2396, RoundKey[117]}), .a ({new_AGEMA_signal_3598, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_3716, RoundKeyOutput[117]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_118_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2399, RoundKey[118]}), .a ({new_AGEMA_signal_3597, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_3717, RoundKeyOutput[118]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_119_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2402, RoundKey[119]}), .a ({new_AGEMA_signal_3596, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_3718, RoundKeyOutput[119]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_120_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2408, RoundKey[120]}), .a ({new_AGEMA_signal_3595, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_3719, RoundKeyOutput[120]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_121_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2411, RoundKey[121]}), .a ({new_AGEMA_signal_3691, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_3859, RoundKeyOutput[121]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_122_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2414, RoundKey[122]}), .a ({new_AGEMA_signal_3690, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_3860, RoundKeyOutput[122]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_123_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2417, RoundKey[123]}), .a ({new_AGEMA_signal_3689, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_3861, RoundKeyOutput[123]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_124_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2420, RoundKey[124]}), .a ({new_AGEMA_signal_3688, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_3862, RoundKeyOutput[124]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_125_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2423, RoundKey[125]}), .a ({new_AGEMA_signal_3687, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_3863, RoundKeyOutput[125]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_126_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2426, RoundKey[126]}), .a ({new_AGEMA_signal_3686, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_3864, RoundKeyOutput[126]}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(0)) MuxKeyExpansion_mux_inst_127_U1 ( .s (MuxKeyExpansion_n14), .b ({new_AGEMA_signal_2429, RoundKey[127]}), .a ({new_AGEMA_signal_3685, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_3865, RoundKeyOutput[127]}) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4156, RoundReg_Inst_ff_SDE_0_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4273, RoundReg_Inst_ff_SDE_1_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4158, RoundReg_Inst_ff_SDE_2_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4275, RoundReg_Inst_ff_SDE_3_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4277, RoundReg_Inst_ff_SDE_4_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4160, RoundReg_Inst_ff_SDE_5_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4162, RoundReg_Inst_ff_SDE_6_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4164, RoundReg_Inst_ff_SDE_7_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4166, RoundReg_Inst_ff_SDE_8_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4279, RoundReg_Inst_ff_SDE_9_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4168, RoundReg_Inst_ff_SDE_10_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4281, RoundReg_Inst_ff_SDE_11_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4283, RoundReg_Inst_ff_SDE_12_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4170, RoundReg_Inst_ff_SDE_13_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4172, RoundReg_Inst_ff_SDE_14_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4174, RoundReg_Inst_ff_SDE_15_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4176, RoundReg_Inst_ff_SDE_16_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4285, RoundReg_Inst_ff_SDE_17_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4178, RoundReg_Inst_ff_SDE_18_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4287, RoundReg_Inst_ff_SDE_19_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4289, RoundReg_Inst_ff_SDE_20_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4180, RoundReg_Inst_ff_SDE_21_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4182, RoundReg_Inst_ff_SDE_22_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4184, RoundReg_Inst_ff_SDE_23_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4186, RoundReg_Inst_ff_SDE_24_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4291, RoundReg_Inst_ff_SDE_25_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4188, RoundReg_Inst_ff_SDE_26_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4293, RoundReg_Inst_ff_SDE_27_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4295, RoundReg_Inst_ff_SDE_28_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4190, RoundReg_Inst_ff_SDE_29_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4192, RoundReg_Inst_ff_SDE_30_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4194, RoundReg_Inst_ff_SDE_31_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2851, RoundReg_Inst_ff_SDE_32_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2853, RoundReg_Inst_ff_SDE_33_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2855, RoundReg_Inst_ff_SDE_34_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2857, RoundReg_Inst_ff_SDE_35_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2859, RoundReg_Inst_ff_SDE_36_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2861, RoundReg_Inst_ff_SDE_37_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2863, RoundReg_Inst_ff_SDE_38_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2865, RoundReg_Inst_ff_SDE_39_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2867, RoundReg_Inst_ff_SDE_40_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2869, RoundReg_Inst_ff_SDE_41_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2871, RoundReg_Inst_ff_SDE_42_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2873, RoundReg_Inst_ff_SDE_43_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2875, RoundReg_Inst_ff_SDE_44_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2877, RoundReg_Inst_ff_SDE_45_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2879, RoundReg_Inst_ff_SDE_46_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2881, RoundReg_Inst_ff_SDE_47_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2883, RoundReg_Inst_ff_SDE_48_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2885, RoundReg_Inst_ff_SDE_49_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2887, RoundReg_Inst_ff_SDE_50_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2889, RoundReg_Inst_ff_SDE_51_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2891, RoundReg_Inst_ff_SDE_52_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2893, RoundReg_Inst_ff_SDE_53_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2895, RoundReg_Inst_ff_SDE_54_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2897, RoundReg_Inst_ff_SDE_55_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2899, RoundReg_Inst_ff_SDE_56_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2901, RoundReg_Inst_ff_SDE_57_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2903, RoundReg_Inst_ff_SDE_58_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2905, RoundReg_Inst_ff_SDE_59_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2907, RoundReg_Inst_ff_SDE_60_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2909, RoundReg_Inst_ff_SDE_61_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2911, RoundReg_Inst_ff_SDE_62_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2913, RoundReg_Inst_ff_SDE_63_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2915, RoundReg_Inst_ff_SDE_64_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2917, RoundReg_Inst_ff_SDE_65_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2919, RoundReg_Inst_ff_SDE_66_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2921, RoundReg_Inst_ff_SDE_67_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2923, RoundReg_Inst_ff_SDE_68_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2925, RoundReg_Inst_ff_SDE_69_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2927, RoundReg_Inst_ff_SDE_70_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2929, RoundReg_Inst_ff_SDE_71_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2931, RoundReg_Inst_ff_SDE_72_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2933, RoundReg_Inst_ff_SDE_73_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2935, RoundReg_Inst_ff_SDE_74_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2937, RoundReg_Inst_ff_SDE_75_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2939, RoundReg_Inst_ff_SDE_76_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2941, RoundReg_Inst_ff_SDE_77_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2943, RoundReg_Inst_ff_SDE_78_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2945, RoundReg_Inst_ff_SDE_79_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2947, RoundReg_Inst_ff_SDE_80_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2949, RoundReg_Inst_ff_SDE_81_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2951, RoundReg_Inst_ff_SDE_82_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2953, RoundReg_Inst_ff_SDE_83_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2955, RoundReg_Inst_ff_SDE_84_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2957, RoundReg_Inst_ff_SDE_85_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2959, RoundReg_Inst_ff_SDE_86_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2961, RoundReg_Inst_ff_SDE_87_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2963, RoundReg_Inst_ff_SDE_88_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2965, RoundReg_Inst_ff_SDE_89_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2967, RoundReg_Inst_ff_SDE_90_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2969, RoundReg_Inst_ff_SDE_91_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2971, RoundReg_Inst_ff_SDE_92_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2973, RoundReg_Inst_ff_SDE_93_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2975, RoundReg_Inst_ff_SDE_94_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2977, RoundReg_Inst_ff_SDE_95_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2979, RoundReg_Inst_ff_SDE_96_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2981, RoundReg_Inst_ff_SDE_97_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2983, RoundReg_Inst_ff_SDE_98_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2985, RoundReg_Inst_ff_SDE_99_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2987, RoundReg_Inst_ff_SDE_100_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2989, RoundReg_Inst_ff_SDE_101_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2991, RoundReg_Inst_ff_SDE_102_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2993, RoundReg_Inst_ff_SDE_103_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2995, RoundReg_Inst_ff_SDE_104_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2997, RoundReg_Inst_ff_SDE_105_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_2999, RoundReg_Inst_ff_SDE_106_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3001, RoundReg_Inst_ff_SDE_107_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3003, RoundReg_Inst_ff_SDE_108_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3005, RoundReg_Inst_ff_SDE_109_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3007, RoundReg_Inst_ff_SDE_110_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3009, RoundReg_Inst_ff_SDE_111_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3011, RoundReg_Inst_ff_SDE_112_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3013, RoundReg_Inst_ff_SDE_113_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3015, RoundReg_Inst_ff_SDE_114_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3017, RoundReg_Inst_ff_SDE_115_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3019, RoundReg_Inst_ff_SDE_116_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3021, RoundReg_Inst_ff_SDE_117_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3023, RoundReg_Inst_ff_SDE_118_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3025, RoundReg_Inst_ff_SDE_119_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3027, RoundReg_Inst_ff_SDE_120_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3029, RoundReg_Inst_ff_SDE_121_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3031, RoundReg_Inst_ff_SDE_122_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3033, RoundReg_Inst_ff_SDE_123_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3035, RoundReg_Inst_ff_SDE_124_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3037, RoundReg_Inst_ff_SDE_125_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3039, RoundReg_Inst_ff_SDE_126_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3041, RoundReg_Inst_ff_SDE_127_next_state}), .clk (clk_gated), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4056, KeyReg_Inst_ff_SDE_0_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2339, KSSubBytesInput[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4208, KeyReg_Inst_ff_SDE_1_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2456, KSSubBytesInput[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4210, KeyReg_Inst_ff_SDE_2_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2489, KSSubBytesInput[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4212, KeyReg_Inst_ff_SDE_3_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2522, KSSubBytesInput[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4214, KeyReg_Inst_ff_SDE_4_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2555, KSSubBytesInput[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4216, KeyReg_Inst_ff_SDE_5_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2588, KSSubBytesInput[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4218, KeyReg_Inst_ff_SDE_6_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2621, KSSubBytesInput[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4220, KeyReg_Inst_ff_SDE_7_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2654, KSSubBytesInput[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4058, KeyReg_Inst_ff_SDE_8_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2687, KSSubBytesInput[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4222, KeyReg_Inst_ff_SDE_9_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2720, KSSubBytesInput[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4224, KeyReg_Inst_ff_SDE_10_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2372, KSSubBytesInput[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4226, KeyReg_Inst_ff_SDE_11_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2405, KSSubBytesInput[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4228, KeyReg_Inst_ff_SDE_12_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2432, KSSubBytesInput[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4230, KeyReg_Inst_ff_SDE_13_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2435, KSSubBytesInput[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4232, KeyReg_Inst_ff_SDE_14_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2438, KSSubBytesInput[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4234, KeyReg_Inst_ff_SDE_15_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2441, KSSubBytesInput[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4060, KeyReg_Inst_ff_SDE_16_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2444, KSSubBytesInput[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4236, KeyReg_Inst_ff_SDE_17_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2447, KSSubBytesInput[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4238, KeyReg_Inst_ff_SDE_18_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2450, KSSubBytesInput[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4240, KeyReg_Inst_ff_SDE_19_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2453, KSSubBytesInput[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4242, KeyReg_Inst_ff_SDE_20_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2459, KSSubBytesInput[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4244, KeyReg_Inst_ff_SDE_21_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2462, KSSubBytesInput[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4246, KeyReg_Inst_ff_SDE_22_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2465, KSSubBytesInput[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4248, KeyReg_Inst_ff_SDE_23_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2468, KSSubBytesInput[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4250, KeyReg_Inst_ff_SDE_24_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2471, KSSubBytesInput[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4297, KeyReg_Inst_ff_SDE_25_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2474, KSSubBytesInput[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4299, KeyReg_Inst_ff_SDE_26_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2477, KSSubBytesInput[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4301, KeyReg_Inst_ff_SDE_27_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2480, KSSubBytesInput[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4303, KeyReg_Inst_ff_SDE_28_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2483, KSSubBytesInput[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4305, KeyReg_Inst_ff_SDE_29_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2486, KSSubBytesInput[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4307, KeyReg_Inst_ff_SDE_30_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2492, KSSubBytesInput[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4309, KeyReg_Inst_ff_SDE_31_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2495, KSSubBytesInput[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3899, KeyReg_Inst_ff_SDE_32_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2498, RoundKey[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4062, KeyReg_Inst_ff_SDE_33_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2501, RoundKey[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4064, KeyReg_Inst_ff_SDE_34_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2504, RoundKey[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4066, KeyReg_Inst_ff_SDE_35_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2507, RoundKey[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4068, KeyReg_Inst_ff_SDE_36_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2510, RoundKey[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4070, KeyReg_Inst_ff_SDE_37_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2513, RoundKey[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4072, KeyReg_Inst_ff_SDE_38_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2516, RoundKey[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4074, KeyReg_Inst_ff_SDE_39_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2519, RoundKey[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3901, KeyReg_Inst_ff_SDE_40_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2525, RoundKey[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4076, KeyReg_Inst_ff_SDE_41_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2528, RoundKey[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4078, KeyReg_Inst_ff_SDE_42_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2531, RoundKey[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4080, KeyReg_Inst_ff_SDE_43_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2534, RoundKey[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4082, KeyReg_Inst_ff_SDE_44_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2537, RoundKey[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4084, KeyReg_Inst_ff_SDE_45_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2540, RoundKey[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4086, KeyReg_Inst_ff_SDE_46_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2543, RoundKey[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4088, KeyReg_Inst_ff_SDE_47_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2546, RoundKey[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3903, KeyReg_Inst_ff_SDE_48_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2549, RoundKey[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4090, KeyReg_Inst_ff_SDE_49_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2552, RoundKey[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4092, KeyReg_Inst_ff_SDE_50_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2558, RoundKey[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4094, KeyReg_Inst_ff_SDE_51_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2561, RoundKey[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4096, KeyReg_Inst_ff_SDE_52_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2564, RoundKey[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4098, KeyReg_Inst_ff_SDE_53_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2567, RoundKey[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4100, KeyReg_Inst_ff_SDE_54_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2570, RoundKey[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4102, KeyReg_Inst_ff_SDE_55_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2573, RoundKey[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4104, KeyReg_Inst_ff_SDE_56_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2576, RoundKey[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4252, KeyReg_Inst_ff_SDE_57_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2579, RoundKey[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4254, KeyReg_Inst_ff_SDE_58_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2582, RoundKey[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4256, KeyReg_Inst_ff_SDE_59_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2585, RoundKey[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4258, KeyReg_Inst_ff_SDE_60_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2591, RoundKey[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4260, KeyReg_Inst_ff_SDE_61_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2594, RoundKey[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4262, KeyReg_Inst_ff_SDE_62_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2597, RoundKey[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4264, KeyReg_Inst_ff_SDE_63_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2600, RoundKey[63]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3753, KeyReg_Inst_ff_SDE_64_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2603, RoundKey[64]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3905, KeyReg_Inst_ff_SDE_65_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2606, RoundKey[65]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3907, KeyReg_Inst_ff_SDE_66_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2609, RoundKey[66]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3909, KeyReg_Inst_ff_SDE_67_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2612, RoundKey[67]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3911, KeyReg_Inst_ff_SDE_68_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2615, RoundKey[68]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3913, KeyReg_Inst_ff_SDE_69_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2618, RoundKey[69]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3915, KeyReg_Inst_ff_SDE_70_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2624, RoundKey[70]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3917, KeyReg_Inst_ff_SDE_71_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2627, RoundKey[71]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3755, KeyReg_Inst_ff_SDE_72_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2630, RoundKey[72]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3919, KeyReg_Inst_ff_SDE_73_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2633, RoundKey[73]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3921, KeyReg_Inst_ff_SDE_74_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2636, RoundKey[74]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3923, KeyReg_Inst_ff_SDE_75_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2639, RoundKey[75]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3925, KeyReg_Inst_ff_SDE_76_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2642, RoundKey[76]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3927, KeyReg_Inst_ff_SDE_77_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2645, RoundKey[77]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3929, KeyReg_Inst_ff_SDE_78_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2648, RoundKey[78]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3931, KeyReg_Inst_ff_SDE_79_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2651, RoundKey[79]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3757, KeyReg_Inst_ff_SDE_80_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2657, RoundKey[80]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3933, KeyReg_Inst_ff_SDE_81_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2660, RoundKey[81]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3935, KeyReg_Inst_ff_SDE_82_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2663, RoundKey[82]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3937, KeyReg_Inst_ff_SDE_83_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2666, RoundKey[83]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3939, KeyReg_Inst_ff_SDE_84_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2669, RoundKey[84]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3941, KeyReg_Inst_ff_SDE_85_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2672, RoundKey[85]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3943, KeyReg_Inst_ff_SDE_86_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2675, RoundKey[86]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3945, KeyReg_Inst_ff_SDE_87_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2678, RoundKey[87]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3947, KeyReg_Inst_ff_SDE_88_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2681, RoundKey[88]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4106, KeyReg_Inst_ff_SDE_89_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2684, RoundKey[89]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4108, KeyReg_Inst_ff_SDE_90_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2690, RoundKey[90]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4110, KeyReg_Inst_ff_SDE_91_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2693, RoundKey[91]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4112, KeyReg_Inst_ff_SDE_92_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2696, RoundKey[92]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4114, KeyReg_Inst_ff_SDE_93_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2699, RoundKey[93]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4116, KeyReg_Inst_ff_SDE_94_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2702, RoundKey[94]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4118, KeyReg_Inst_ff_SDE_95_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2705, RoundKey[95]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3658, KeyReg_Inst_ff_SDE_96_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2708, RoundKey[96]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3759, KeyReg_Inst_ff_SDE_97_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2711, RoundKey[97]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3761, KeyReg_Inst_ff_SDE_98_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2714, RoundKey[98]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3763, KeyReg_Inst_ff_SDE_99_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2717, RoundKey[99]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3765, KeyReg_Inst_ff_SDE_100_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2342, RoundKey[100]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3767, KeyReg_Inst_ff_SDE_101_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2345, RoundKey[101]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3769, KeyReg_Inst_ff_SDE_102_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2348, RoundKey[102]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3771, KeyReg_Inst_ff_SDE_103_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2351, RoundKey[103]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3660, KeyReg_Inst_ff_SDE_104_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2354, RoundKey[104]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3773, KeyReg_Inst_ff_SDE_105_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2357, RoundKey[105]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3775, KeyReg_Inst_ff_SDE_106_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2360, RoundKey[106]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3777, KeyReg_Inst_ff_SDE_107_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2363, RoundKey[107]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3779, KeyReg_Inst_ff_SDE_108_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2366, RoundKey[108]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3781, KeyReg_Inst_ff_SDE_109_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2369, RoundKey[109]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3783, KeyReg_Inst_ff_SDE_110_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2375, RoundKey[110]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3785, KeyReg_Inst_ff_SDE_111_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2378, RoundKey[111]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3662, KeyReg_Inst_ff_SDE_112_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2381, RoundKey[112]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3787, KeyReg_Inst_ff_SDE_113_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2384, RoundKey[113]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3789, KeyReg_Inst_ff_SDE_114_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2387, RoundKey[114]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3791, KeyReg_Inst_ff_SDE_115_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2390, RoundKey[115]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3793, KeyReg_Inst_ff_SDE_116_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2393, RoundKey[116]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3795, KeyReg_Inst_ff_SDE_117_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2396, RoundKey[117]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3797, KeyReg_Inst_ff_SDE_118_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2399, RoundKey[118]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3799, KeyReg_Inst_ff_SDE_119_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2402, RoundKey[119]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3801, KeyReg_Inst_ff_SDE_120_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2408, RoundKey[120]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3949, KeyReg_Inst_ff_SDE_121_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2411, RoundKey[121]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3951, KeyReg_Inst_ff_SDE_122_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2414, RoundKey[122]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3953, KeyReg_Inst_ff_SDE_123_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2417, RoundKey[123]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3955, KeyReg_Inst_ff_SDE_124_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2420, RoundKey[124]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3957, KeyReg_Inst_ff_SDE_125_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2423, RoundKey[125]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3959, KeyReg_Inst_ff_SDE_126_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2426, RoundKey[126]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3961, KeyReg_Inst_ff_SDE_127_next_state}), .clk (clk_gated), .Q ({new_AGEMA_signal_2429, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D (RoundCounterIns_n45), .CK (clk_gated), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D (RoundCounterIns_n44), .CK (clk_gated), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D (RoundCounterIns_n1), .CK (clk_gated), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D (RoundCounterIns_n42), .CK (clk_gated), .Q (RoundCounter[3]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_0__FF_FF ( .D (InRoundCounterIns_n41), .CK (clk_gated), .Q (InRoundCounter[0]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_1__FF_FF ( .D (InRoundCounterIns_n40), .CK (clk_gated), .Q (InRoundCounter[1]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_2__FF_FF ( .D (InRoundCounterIns_n39), .CK (clk_gated), .Q (InRoundCounter[2]), .QN () ) ;
endmodule
