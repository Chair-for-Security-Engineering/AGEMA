/* modified netlist. Source: module CRAFT in file Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module CRAFT_HPC2_ClockGating_d3 (plaintext_s0, key_s0, clk, rst, key_s1, key_s2, key_s3, plaintext_s1, plaintext_s2, plaintext_s3, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, ciphertext_s3, Synch);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] key_s3 ;
    input [63:0] plaintext_s1 ;
    input [63:0] plaintext_s2 ;
    input [63:0] plaintext_s3 ;
    input [1535:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    output [63:0] ciphertext_s2 ;
    output [63:0] ciphertext_s3 ;
    output Synch ;
    wire RoundConstant_4_ ;
    wire RoundConstant_0 ;
    wire done_internal ;
    wire MCInst_XOR_r0_Inst_0_n2 ;
    wire MCInst_XOR_r0_Inst_0_n1 ;
    wire MCInst_XOR_r1_Inst_0_n1 ;
    wire MCInst_XOR_r0_Inst_1_n2 ;
    wire MCInst_XOR_r0_Inst_1_n1 ;
    wire MCInst_XOR_r1_Inst_1_n1 ;
    wire MCInst_XOR_r0_Inst_2_n2 ;
    wire MCInst_XOR_r0_Inst_2_n1 ;
    wire MCInst_XOR_r1_Inst_2_n1 ;
    wire MCInst_XOR_r0_Inst_3_n2 ;
    wire MCInst_XOR_r0_Inst_3_n1 ;
    wire MCInst_XOR_r1_Inst_3_n1 ;
    wire MCInst_XOR_r0_Inst_4_n2 ;
    wire MCInst_XOR_r0_Inst_4_n1 ;
    wire MCInst_XOR_r1_Inst_4_n1 ;
    wire MCInst_XOR_r0_Inst_5_n2 ;
    wire MCInst_XOR_r0_Inst_5_n1 ;
    wire MCInst_XOR_r1_Inst_5_n1 ;
    wire MCInst_XOR_r0_Inst_6_n2 ;
    wire MCInst_XOR_r0_Inst_6_n1 ;
    wire MCInst_XOR_r1_Inst_6_n1 ;
    wire MCInst_XOR_r0_Inst_7_n2 ;
    wire MCInst_XOR_r0_Inst_7_n1 ;
    wire MCInst_XOR_r1_Inst_7_n1 ;
    wire MCInst_XOR_r0_Inst_8_n2 ;
    wire MCInst_XOR_r0_Inst_8_n1 ;
    wire MCInst_XOR_r1_Inst_8_n1 ;
    wire MCInst_XOR_r0_Inst_9_n2 ;
    wire MCInst_XOR_r0_Inst_9_n1 ;
    wire MCInst_XOR_r1_Inst_9_n1 ;
    wire MCInst_XOR_r0_Inst_10_n2 ;
    wire MCInst_XOR_r0_Inst_10_n1 ;
    wire MCInst_XOR_r1_Inst_10_n1 ;
    wire MCInst_XOR_r0_Inst_11_n2 ;
    wire MCInst_XOR_r0_Inst_11_n1 ;
    wire MCInst_XOR_r1_Inst_11_n1 ;
    wire MCInst_XOR_r0_Inst_12_n2 ;
    wire MCInst_XOR_r0_Inst_12_n1 ;
    wire MCInst_XOR_r1_Inst_12_n1 ;
    wire MCInst_XOR_r0_Inst_13_n2 ;
    wire MCInst_XOR_r0_Inst_13_n1 ;
    wire MCInst_XOR_r1_Inst_13_n1 ;
    wire MCInst_XOR_r0_Inst_14_n2 ;
    wire MCInst_XOR_r0_Inst_14_n1 ;
    wire MCInst_XOR_r1_Inst_14_n1 ;
    wire MCInst_XOR_r0_Inst_15_n2 ;
    wire MCInst_XOR_r0_Inst_15_n1 ;
    wire MCInst_XOR_r1_Inst_15_n1 ;
    wire AddKeyXOR1_XORInst_0_0_n1 ;
    wire AddKeyXOR1_XORInst_0_1_n1 ;
    wire AddKeyXOR1_XORInst_0_2_n1 ;
    wire AddKeyXOR1_XORInst_0_3_n1 ;
    wire AddKeyXOR1_XORInst_1_0_n1 ;
    wire AddKeyXOR1_XORInst_1_1_n1 ;
    wire AddKeyXOR1_XORInst_1_2_n1 ;
    wire AddKeyXOR1_XORInst_1_3_n1 ;
    wire AddKeyXOR1_XORInst_2_0_n1 ;
    wire AddKeyXOR1_XORInst_2_1_n1 ;
    wire AddKeyXOR1_XORInst_2_2_n1 ;
    wire AddKeyXOR1_XORInst_2_3_n1 ;
    wire AddKeyXOR1_XORInst_3_0_n1 ;
    wire AddKeyXOR1_XORInst_3_1_n1 ;
    wire AddKeyXOR1_XORInst_3_2_n1 ;
    wire AddKeyXOR1_XORInst_3_3_n1 ;
    wire AddKeyConstXOR_XORInst_0_0_n2 ;
    wire AddKeyConstXOR_XORInst_0_0_n1 ;
    wire AddKeyConstXOR_XORInst_0_1_n2 ;
    wire AddKeyConstXOR_XORInst_0_1_n1 ;
    wire AddKeyConstXOR_XORInst_0_2_n2 ;
    wire AddKeyConstXOR_XORInst_0_2_n1 ;
    wire AddKeyConstXOR_XORInst_0_3_n2 ;
    wire AddKeyConstXOR_XORInst_0_3_n1 ;
    wire AddKeyConstXOR_XORInst_1_0_n2 ;
    wire AddKeyConstXOR_XORInst_1_0_n1 ;
    wire AddKeyConstXOR_XORInst_1_1_n2 ;
    wire AddKeyConstXOR_XORInst_1_1_n1 ;
    wire AddKeyConstXOR_XORInst_1_2_n2 ;
    wire AddKeyConstXOR_XORInst_1_2_n1 ;
    wire AddKeyConstXOR_XORInst_1_3_n2 ;
    wire AddKeyConstXOR_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_0_0_n1 ;
    wire AddKeyXOR2_XORInst_0_1_n1 ;
    wire AddKeyXOR2_XORInst_0_2_n1 ;
    wire AddKeyXOR2_XORInst_0_3_n1 ;
    wire AddKeyXOR2_XORInst_1_0_n1 ;
    wire AddKeyXOR2_XORInst_1_1_n1 ;
    wire AddKeyXOR2_XORInst_1_2_n1 ;
    wire AddKeyXOR2_XORInst_1_3_n1 ;
    wire AddKeyXOR2_XORInst_2_0_n1 ;
    wire AddKeyXOR2_XORInst_2_1_n1 ;
    wire AddKeyXOR2_XORInst_2_2_n1 ;
    wire AddKeyXOR2_XORInst_2_3_n1 ;
    wire AddKeyXOR2_XORInst_3_0_n1 ;
    wire AddKeyXOR2_XORInst_3_1_n1 ;
    wire AddKeyXOR2_XORInst_3_2_n1 ;
    wire AddKeyXOR2_XORInst_3_3_n1 ;
    wire AddKeyXOR2_XORInst_4_0_n1 ;
    wire AddKeyXOR2_XORInst_4_1_n1 ;
    wire AddKeyXOR2_XORInst_4_2_n1 ;
    wire AddKeyXOR2_XORInst_4_3_n1 ;
    wire AddKeyXOR2_XORInst_5_0_n1 ;
    wire AddKeyXOR2_XORInst_5_1_n1 ;
    wire AddKeyXOR2_XORInst_5_2_n1 ;
    wire AddKeyXOR2_XORInst_5_3_n1 ;
    wire AddKeyXOR2_XORInst_6_0_n1 ;
    wire AddKeyXOR2_XORInst_6_1_n1 ;
    wire AddKeyXOR2_XORInst_6_2_n1 ;
    wire AddKeyXOR2_XORInst_6_3_n1 ;
    wire AddKeyXOR2_XORInst_7_0_n1 ;
    wire AddKeyXOR2_XORInst_7_1_n1 ;
    wire AddKeyXOR2_XORInst_7_2_n1 ;
    wire AddKeyXOR2_XORInst_7_3_n1 ;
    wire AddKeyXOR2_XORInst_8_0_n1 ;
    wire AddKeyXOR2_XORInst_8_1_n1 ;
    wire AddKeyXOR2_XORInst_8_2_n1 ;
    wire AddKeyXOR2_XORInst_8_3_n1 ;
    wire AddKeyXOR2_XORInst_9_0_n1 ;
    wire AddKeyXOR2_XORInst_9_1_n1 ;
    wire AddKeyXOR2_XORInst_9_2_n1 ;
    wire AddKeyXOR2_XORInst_9_3_n1 ;
    wire SubCellInst_SboxInst_0_n15 ;
    wire SubCellInst_SboxInst_0_n14 ;
    wire SubCellInst_SboxInst_0_n13 ;
    wire SubCellInst_SboxInst_0_n12 ;
    wire SubCellInst_SboxInst_0_n11 ;
    wire SubCellInst_SboxInst_0_n10 ;
    wire SubCellInst_SboxInst_0_n9 ;
    wire SubCellInst_SboxInst_0_n8 ;
    wire SubCellInst_SboxInst_0_n7 ;
    wire SubCellInst_SboxInst_0_n6 ;
    wire SubCellInst_SboxInst_0_n5 ;
    wire SubCellInst_SboxInst_0_n4 ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_n2 ;
    wire SubCellInst_SboxInst_0_n1 ;
    wire SubCellInst_SboxInst_1_n15 ;
    wire SubCellInst_SboxInst_1_n14 ;
    wire SubCellInst_SboxInst_1_n13 ;
    wire SubCellInst_SboxInst_1_n12 ;
    wire SubCellInst_SboxInst_1_n11 ;
    wire SubCellInst_SboxInst_1_n10 ;
    wire SubCellInst_SboxInst_1_n9 ;
    wire SubCellInst_SboxInst_1_n8 ;
    wire SubCellInst_SboxInst_1_n7 ;
    wire SubCellInst_SboxInst_1_n6 ;
    wire SubCellInst_SboxInst_1_n5 ;
    wire SubCellInst_SboxInst_1_n4 ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_n2 ;
    wire SubCellInst_SboxInst_1_n1 ;
    wire SubCellInst_SboxInst_2_n15 ;
    wire SubCellInst_SboxInst_2_n14 ;
    wire SubCellInst_SboxInst_2_n13 ;
    wire SubCellInst_SboxInst_2_n12 ;
    wire SubCellInst_SboxInst_2_n11 ;
    wire SubCellInst_SboxInst_2_n10 ;
    wire SubCellInst_SboxInst_2_n9 ;
    wire SubCellInst_SboxInst_2_n8 ;
    wire SubCellInst_SboxInst_2_n7 ;
    wire SubCellInst_SboxInst_2_n6 ;
    wire SubCellInst_SboxInst_2_n5 ;
    wire SubCellInst_SboxInst_2_n4 ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_n2 ;
    wire SubCellInst_SboxInst_2_n1 ;
    wire SubCellInst_SboxInst_3_n15 ;
    wire SubCellInst_SboxInst_3_n14 ;
    wire SubCellInst_SboxInst_3_n13 ;
    wire SubCellInst_SboxInst_3_n12 ;
    wire SubCellInst_SboxInst_3_n11 ;
    wire SubCellInst_SboxInst_3_n10 ;
    wire SubCellInst_SboxInst_3_n9 ;
    wire SubCellInst_SboxInst_3_n8 ;
    wire SubCellInst_SboxInst_3_n7 ;
    wire SubCellInst_SboxInst_3_n6 ;
    wire SubCellInst_SboxInst_3_n5 ;
    wire SubCellInst_SboxInst_3_n4 ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_n2 ;
    wire SubCellInst_SboxInst_3_n1 ;
    wire SubCellInst_SboxInst_4_n15 ;
    wire SubCellInst_SboxInst_4_n14 ;
    wire SubCellInst_SboxInst_4_n13 ;
    wire SubCellInst_SboxInst_4_n12 ;
    wire SubCellInst_SboxInst_4_n11 ;
    wire SubCellInst_SboxInst_4_n10 ;
    wire SubCellInst_SboxInst_4_n9 ;
    wire SubCellInst_SboxInst_4_n8 ;
    wire SubCellInst_SboxInst_4_n7 ;
    wire SubCellInst_SboxInst_4_n6 ;
    wire SubCellInst_SboxInst_4_n5 ;
    wire SubCellInst_SboxInst_4_n4 ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_n2 ;
    wire SubCellInst_SboxInst_4_n1 ;
    wire SubCellInst_SboxInst_5_n15 ;
    wire SubCellInst_SboxInst_5_n14 ;
    wire SubCellInst_SboxInst_5_n13 ;
    wire SubCellInst_SboxInst_5_n12 ;
    wire SubCellInst_SboxInst_5_n11 ;
    wire SubCellInst_SboxInst_5_n10 ;
    wire SubCellInst_SboxInst_5_n9 ;
    wire SubCellInst_SboxInst_5_n8 ;
    wire SubCellInst_SboxInst_5_n7 ;
    wire SubCellInst_SboxInst_5_n6 ;
    wire SubCellInst_SboxInst_5_n5 ;
    wire SubCellInst_SboxInst_5_n4 ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_n2 ;
    wire SubCellInst_SboxInst_5_n1 ;
    wire SubCellInst_SboxInst_6_n15 ;
    wire SubCellInst_SboxInst_6_n14 ;
    wire SubCellInst_SboxInst_6_n13 ;
    wire SubCellInst_SboxInst_6_n12 ;
    wire SubCellInst_SboxInst_6_n11 ;
    wire SubCellInst_SboxInst_6_n10 ;
    wire SubCellInst_SboxInst_6_n9 ;
    wire SubCellInst_SboxInst_6_n8 ;
    wire SubCellInst_SboxInst_6_n7 ;
    wire SubCellInst_SboxInst_6_n6 ;
    wire SubCellInst_SboxInst_6_n5 ;
    wire SubCellInst_SboxInst_6_n4 ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_n2 ;
    wire SubCellInst_SboxInst_6_n1 ;
    wire SubCellInst_SboxInst_7_n15 ;
    wire SubCellInst_SboxInst_7_n14 ;
    wire SubCellInst_SboxInst_7_n13 ;
    wire SubCellInst_SboxInst_7_n12 ;
    wire SubCellInst_SboxInst_7_n11 ;
    wire SubCellInst_SboxInst_7_n10 ;
    wire SubCellInst_SboxInst_7_n9 ;
    wire SubCellInst_SboxInst_7_n8 ;
    wire SubCellInst_SboxInst_7_n7 ;
    wire SubCellInst_SboxInst_7_n6 ;
    wire SubCellInst_SboxInst_7_n5 ;
    wire SubCellInst_SboxInst_7_n4 ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_n2 ;
    wire SubCellInst_SboxInst_7_n1 ;
    wire SubCellInst_SboxInst_8_n15 ;
    wire SubCellInst_SboxInst_8_n14 ;
    wire SubCellInst_SboxInst_8_n13 ;
    wire SubCellInst_SboxInst_8_n12 ;
    wire SubCellInst_SboxInst_8_n11 ;
    wire SubCellInst_SboxInst_8_n10 ;
    wire SubCellInst_SboxInst_8_n9 ;
    wire SubCellInst_SboxInst_8_n8 ;
    wire SubCellInst_SboxInst_8_n7 ;
    wire SubCellInst_SboxInst_8_n6 ;
    wire SubCellInst_SboxInst_8_n5 ;
    wire SubCellInst_SboxInst_8_n4 ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_n2 ;
    wire SubCellInst_SboxInst_8_n1 ;
    wire SubCellInst_SboxInst_9_n15 ;
    wire SubCellInst_SboxInst_9_n14 ;
    wire SubCellInst_SboxInst_9_n13 ;
    wire SubCellInst_SboxInst_9_n12 ;
    wire SubCellInst_SboxInst_9_n11 ;
    wire SubCellInst_SboxInst_9_n10 ;
    wire SubCellInst_SboxInst_9_n9 ;
    wire SubCellInst_SboxInst_9_n8 ;
    wire SubCellInst_SboxInst_9_n7 ;
    wire SubCellInst_SboxInst_9_n6 ;
    wire SubCellInst_SboxInst_9_n5 ;
    wire SubCellInst_SboxInst_9_n4 ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_n2 ;
    wire SubCellInst_SboxInst_9_n1 ;
    wire SubCellInst_SboxInst_10_n15 ;
    wire SubCellInst_SboxInst_10_n14 ;
    wire SubCellInst_SboxInst_10_n13 ;
    wire SubCellInst_SboxInst_10_n12 ;
    wire SubCellInst_SboxInst_10_n11 ;
    wire SubCellInst_SboxInst_10_n10 ;
    wire SubCellInst_SboxInst_10_n9 ;
    wire SubCellInst_SboxInst_10_n8 ;
    wire SubCellInst_SboxInst_10_n7 ;
    wire SubCellInst_SboxInst_10_n6 ;
    wire SubCellInst_SboxInst_10_n5 ;
    wire SubCellInst_SboxInst_10_n4 ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_n2 ;
    wire SubCellInst_SboxInst_10_n1 ;
    wire SubCellInst_SboxInst_11_n15 ;
    wire SubCellInst_SboxInst_11_n14 ;
    wire SubCellInst_SboxInst_11_n13 ;
    wire SubCellInst_SboxInst_11_n12 ;
    wire SubCellInst_SboxInst_11_n11 ;
    wire SubCellInst_SboxInst_11_n10 ;
    wire SubCellInst_SboxInst_11_n9 ;
    wire SubCellInst_SboxInst_11_n8 ;
    wire SubCellInst_SboxInst_11_n7 ;
    wire SubCellInst_SboxInst_11_n6 ;
    wire SubCellInst_SboxInst_11_n5 ;
    wire SubCellInst_SboxInst_11_n4 ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_n2 ;
    wire SubCellInst_SboxInst_11_n1 ;
    wire SubCellInst_SboxInst_12_n15 ;
    wire SubCellInst_SboxInst_12_n14 ;
    wire SubCellInst_SboxInst_12_n13 ;
    wire SubCellInst_SboxInst_12_n12 ;
    wire SubCellInst_SboxInst_12_n11 ;
    wire SubCellInst_SboxInst_12_n10 ;
    wire SubCellInst_SboxInst_12_n9 ;
    wire SubCellInst_SboxInst_12_n8 ;
    wire SubCellInst_SboxInst_12_n7 ;
    wire SubCellInst_SboxInst_12_n6 ;
    wire SubCellInst_SboxInst_12_n5 ;
    wire SubCellInst_SboxInst_12_n4 ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_n2 ;
    wire SubCellInst_SboxInst_12_n1 ;
    wire SubCellInst_SboxInst_13_n15 ;
    wire SubCellInst_SboxInst_13_n14 ;
    wire SubCellInst_SboxInst_13_n13 ;
    wire SubCellInst_SboxInst_13_n12 ;
    wire SubCellInst_SboxInst_13_n11 ;
    wire SubCellInst_SboxInst_13_n10 ;
    wire SubCellInst_SboxInst_13_n9 ;
    wire SubCellInst_SboxInst_13_n8 ;
    wire SubCellInst_SboxInst_13_n7 ;
    wire SubCellInst_SboxInst_13_n6 ;
    wire SubCellInst_SboxInst_13_n5 ;
    wire SubCellInst_SboxInst_13_n4 ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_n2 ;
    wire SubCellInst_SboxInst_13_n1 ;
    wire SubCellInst_SboxInst_14_n15 ;
    wire SubCellInst_SboxInst_14_n14 ;
    wire SubCellInst_SboxInst_14_n13 ;
    wire SubCellInst_SboxInst_14_n12 ;
    wire SubCellInst_SboxInst_14_n11 ;
    wire SubCellInst_SboxInst_14_n10 ;
    wire SubCellInst_SboxInst_14_n9 ;
    wire SubCellInst_SboxInst_14_n8 ;
    wire SubCellInst_SboxInst_14_n7 ;
    wire SubCellInst_SboxInst_14_n6 ;
    wire SubCellInst_SboxInst_14_n5 ;
    wire SubCellInst_SboxInst_14_n4 ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_n2 ;
    wire SubCellInst_SboxInst_14_n1 ;
    wire SubCellInst_SboxInst_15_n15 ;
    wire SubCellInst_SboxInst_15_n14 ;
    wire SubCellInst_SboxInst_15_n13 ;
    wire SubCellInst_SboxInst_15_n12 ;
    wire SubCellInst_SboxInst_15_n11 ;
    wire SubCellInst_SboxInst_15_n10 ;
    wire SubCellInst_SboxInst_15_n9 ;
    wire SubCellInst_SboxInst_15_n8 ;
    wire SubCellInst_SboxInst_15_n7 ;
    wire SubCellInst_SboxInst_15_n6 ;
    wire SubCellInst_SboxInst_15_n5 ;
    wire SubCellInst_SboxInst_15_n4 ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_n2 ;
    wire SubCellInst_SboxInst_15_n1 ;
    wire KeyMUX_n9 ;
    wire KeyMUX_n8 ;
    wire KeyMUX_n7 ;
    wire FSMSignalsInst_n5 ;
    wire FSMSignalsInst_n4 ;
    wire FSMSignalsInst_n3 ;
    wire FSMSignalsInst_n2 ;
    wire FSMSignalsInst_n1 ;
    wire selectsUpdateInst_n3 ;
    wire [63:0] Feedback ;
    wire [63:32] MCInput ;
    wire [63:0] MCOutput ;
    wire [63:0] SelectedKey ;
    wire [63:0] AddRoundKeyOutput ;
    wire [1:0] selects ;
    wire [6:0] FSMReg ;
    wire [6:0] FSMUpdate ;
    wire [1:0] selectsReg ;
    wire [1:0] selectsNext ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, SelectedKey[40]}), .b ({1'b0, 1'b0, 1'b0, RoundConstant_0}), .c ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, AddKeyConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, SelectedKey[41]}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[0]}), .c ({new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, AddKeyConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, SelectedKey[42]}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, AddKeyConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, SelectedKey[43]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, new_AGEMA_signal_3092, AddKeyConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, new_AGEMA_signal_2570, SelectedKey[44]}), .b ({1'b0, 1'b0, 1'b0, RoundConstant_4_}), .c ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, AddKeyConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, new_AGEMA_signal_2579, SelectedKey[45]}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, AddKeyConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, new_AGEMA_signal_2588, SelectedKey[46]}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, new_AGEMA_signal_3101, AddKeyConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, new_AGEMA_signal_2597, SelectedKey[47]}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[5]}), .c ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, AddKeyConstXOR_XORInst_1_3_n1}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U4 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, SubCellInst_SboxInst_0_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U2 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U1 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1042, new_AGEMA_signal_1041, new_AGEMA_signal_1040, SubCellInst_SboxInst_0_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U4 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, SubCellInst_SboxInst_1_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U2 ( .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_1_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U1 ( .a ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, new_AGEMA_signal_1064, SubCellInst_SboxInst_1_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U4 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, SubCellInst_SboxInst_2_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U2 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_2_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U1 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, SubCellInst_SboxInst_2_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U4 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, SubCellInst_SboxInst_3_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U2 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_3_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U1 ( .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, SubCellInst_SboxInst_3_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U4 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, SubCellInst_SboxInst_4_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U2 ( .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_4_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U1 ( .a ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, SubCellInst_SboxInst_4_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U4 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, SubCellInst_SboxInst_5_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U2 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_5_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U1 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, SubCellInst_SboxInst_5_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U4 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_6_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U2 ( .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_6_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U1 ( .a ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, SubCellInst_SboxInst_6_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U4 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_7_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U2 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_7_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U1 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, new_AGEMA_signal_1208, SubCellInst_SboxInst_7_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U4 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_8_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U2 ( .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_8_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U1 ( .a ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, SubCellInst_SboxInst_8_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U4 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_9_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U2 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_9_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U1 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, SubCellInst_SboxInst_9_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U4 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_10_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U2 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_10_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U1 ( .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, new_AGEMA_signal_1280, SubCellInst_SboxInst_10_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U4 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U2 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_11_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U1 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, SubCellInst_SboxInst_11_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U4 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_12_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U2 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_12_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U1 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, SubCellInst_SboxInst_12_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U4 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_13_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U2 ( .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_13_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U1 ( .a ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, new_AGEMA_signal_1352, SubCellInst_SboxInst_13_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U4 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, new_AGEMA_signal_1370, SubCellInst_SboxInst_14_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U2 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_14_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U1 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, SubCellInst_SboxInst_14_n9}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U4 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, SubCellInst_SboxInst_15_n7}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U2 ( .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_15_n8}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U1 ( .a ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, SubCellInst_SboxInst_15_n9}) ) ;
    INV_X1 KeyMUX_U3 ( .A (selects[0]), .ZN (KeyMUX_n9) ) ;
    INV_X1 KeyMUX_U2 ( .A (KeyMUX_n9), .ZN (KeyMUX_n8) ) ;
    INV_X1 KeyMUX_U1 ( .A (KeyMUX_n9), .ZN (KeyMUX_n7) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_0_U1 ( .s (selects[0]), .b ({key_s3[64], key_s2[64], key_s1[64], key_s0[64]}), .a ({key_s3[0], key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, SelectedKey[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_1_U1 ( .s (KeyMUX_n8), .b ({key_s3[65], key_s2[65], key_s1[65], key_s0[65]}), .a ({key_s3[1], key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, SelectedKey[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_2_U1 ( .s (selects[0]), .b ({key_s3[66], key_s2[66], key_s1[66], key_s0[66]}), .a ({key_s3[2], key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, SelectedKey[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_3_U1 ( .s (KeyMUX_n8), .b ({key_s3[67], key_s2[67], key_s1[67], key_s0[67]}), .a ({key_s3[3], key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, new_AGEMA_signal_2282, SelectedKey[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_4_U1 ( .s (KeyMUX_n8), .b ({key_s3[68], key_s2[68], key_s1[68], key_s0[68]}), .a ({key_s3[4], key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, SelectedKey[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_5_U1 ( .s (KeyMUX_n8), .b ({key_s3[69], key_s2[69], key_s1[69], key_s0[69]}), .a ({key_s3[5], key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, SelectedKey[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_6_U1 ( .s (KeyMUX_n8), .b ({key_s3[70], key_s2[70], key_s1[70], key_s0[70]}), .a ({key_s3[6], key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, SelectedKey[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_7_U1 ( .s (KeyMUX_n8), .b ({key_s3[71], key_s2[71], key_s1[71], key_s0[71]}), .a ({key_s3[7], key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, SelectedKey[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_8_U1 ( .s (KeyMUX_n8), .b ({key_s3[72], key_s2[72], key_s1[72], key_s0[72]}), .a ({key_s3[8], key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, SelectedKey[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_9_U1 ( .s (KeyMUX_n8), .b ({key_s3[73], key_s2[73], key_s1[73], key_s0[73]}), .a ({key_s3[9], key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, new_AGEMA_signal_2336, SelectedKey[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_10_U1 ( .s (KeyMUX_n8), .b ({key_s3[74], key_s2[74], key_s1[74], key_s0[74]}), .a ({key_s3[10], key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, SelectedKey[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_11_U1 ( .s (KeyMUX_n8), .b ({key_s3[75], key_s2[75], key_s1[75], key_s0[75]}), .a ({key_s3[11], key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, SelectedKey[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_12_U1 ( .s (KeyMUX_n8), .b ({key_s3[76], key_s2[76], key_s1[76], key_s0[76]}), .a ({key_s3[12], key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, SelectedKey[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_13_U1 ( .s (KeyMUX_n8), .b ({key_s3[77], key_s2[77], key_s1[77], key_s0[77]}), .a ({key_s3[13], key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, new_AGEMA_signal_2372, SelectedKey[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_14_U1 ( .s (KeyMUX_n8), .b ({key_s3[78], key_s2[78], key_s1[78], key_s0[78]}), .a ({key_s3[14], key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, SelectedKey[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_15_U1 ( .s (KeyMUX_n8), .b ({key_s3[79], key_s2[79], key_s1[79], key_s0[79]}), .a ({key_s3[15], key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, new_AGEMA_signal_2390, SelectedKey[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_16_U1 ( .s (KeyMUX_n8), .b ({key_s3[80], key_s2[80], key_s1[80], key_s0[80]}), .a ({key_s3[16], key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, SelectedKey[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_17_U1 ( .s (KeyMUX_n8), .b ({key_s3[81], key_s2[81], key_s1[81], key_s0[81]}), .a ({key_s3[17], key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, SelectedKey[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_18_U1 ( .s (KeyMUX_n8), .b ({key_s3[82], key_s2[82], key_s1[82], key_s0[82]}), .a ({key_s3[18], key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, SelectedKey[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_19_U1 ( .s (KeyMUX_n8), .b ({key_s3[83], key_s2[83], key_s1[83], key_s0[83]}), .a ({key_s3[19], key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, SelectedKey[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_20_U1 ( .s (KeyMUX_n8), .b ({key_s3[84], key_s2[84], key_s1[84], key_s0[84]}), .a ({key_s3[20], key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, SelectedKey[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_21_U1 ( .s (KeyMUX_n8), .b ({key_s3[85], key_s2[85], key_s1[85], key_s0[85]}), .a ({key_s3[21], key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, SelectedKey[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_22_U1 ( .s (selects[0]), .b ({key_s3[86], key_s2[86], key_s1[86], key_s0[86]}), .a ({key_s3[22], key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, SelectedKey[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_23_U1 ( .s (selects[0]), .b ({key_s3[87], key_s2[87], key_s1[87], key_s0[87]}), .a ({key_s3[23], key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, new_AGEMA_signal_1724, SelectedKey[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_24_U1 ( .s (selects[0]), .b ({key_s3[88], key_s2[88], key_s1[88], key_s0[88]}), .a ({key_s3[24], key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, new_AGEMA_signal_1733, SelectedKey[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_25_U1 ( .s (selects[0]), .b ({key_s3[89], key_s2[89], key_s1[89], key_s0[89]}), .a ({key_s3[25], key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, SelectedKey[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_26_U1 ( .s (selects[0]), .b ({key_s3[90], key_s2[90], key_s1[90], key_s0[90]}), .a ({key_s3[26], key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, SelectedKey[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_27_U1 ( .s (selects[0]), .b ({key_s3[91], key_s2[91], key_s1[91], key_s0[91]}), .a ({key_s3[27], key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, SelectedKey[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_28_U1 ( .s (KeyMUX_n7), .b ({key_s3[92], key_s2[92], key_s1[92], key_s0[92]}), .a ({key_s3[28], key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, SelectedKey[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_29_U1 ( .s (KeyMUX_n7), .b ({key_s3[93], key_s2[93], key_s1[93], key_s0[93]}), .a ({key_s3[29], key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, SelectedKey[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_30_U1 ( .s (KeyMUX_n7), .b ({key_s3[94], key_s2[94], key_s1[94], key_s0[94]}), .a ({key_s3[30], key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, SelectedKey[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_31_U1 ( .s (KeyMUX_n7), .b ({key_s3[95], key_s2[95], key_s1[95], key_s0[95]}), .a ({key_s3[31], key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, SelectedKey[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_32_U1 ( .s (KeyMUX_n7), .b ({key_s3[96], key_s2[96], key_s1[96], key_s0[96]}), .a ({key_s3[32], key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, SelectedKey[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_33_U1 ( .s (selects[0]), .b ({key_s3[97], key_s2[97], key_s1[97], key_s0[97]}), .a ({key_s3[33], key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, new_AGEMA_signal_1769, SelectedKey[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_34_U1 ( .s (KeyMUX_n7), .b ({key_s3[98], key_s2[98], key_s1[98], key_s0[98]}), .a ({key_s3[34], key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, SelectedKey[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_35_U1 ( .s (KeyMUX_n7), .b ({key_s3[99], key_s2[99], key_s1[99], key_s0[99]}), .a ({key_s3[35], key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, SelectedKey[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_36_U1 ( .s (selects[0]), .b ({key_s3[100], key_s2[100], key_s1[100], key_s0[100]}), .a ({key_s3[36], key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, new_AGEMA_signal_1778, SelectedKey[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_37_U1 ( .s (KeyMUX_n7), .b ({key_s3[101], key_s2[101], key_s1[101], key_s0[101]}), .a ({key_s3[37], key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, new_AGEMA_signal_2516, SelectedKey[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_38_U1 ( .s (KeyMUX_n7), .b ({key_s3[102], key_s2[102], key_s1[102], key_s0[102]}), .a ({key_s3[38], key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, new_AGEMA_signal_2525, SelectedKey[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_39_U1 ( .s (selects[0]), .b ({key_s3[103], key_s2[103], key_s1[103], key_s0[103]}), .a ({key_s3[39], key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, SelectedKey[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_40_U1 ( .s (KeyMUX_n7), .b ({key_s3[104], key_s2[104], key_s1[104], key_s0[104]}), .a ({key_s3[40], key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_2536, new_AGEMA_signal_2535, new_AGEMA_signal_2534, SelectedKey[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_41_U1 ( .s (KeyMUX_n7), .b ({key_s3[105], key_s2[105], key_s1[105], key_s0[105]}), .a ({key_s3[41], key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, new_AGEMA_signal_2543, SelectedKey[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_42_U1 ( .s (KeyMUX_n7), .b ({key_s3[106], key_s2[106], key_s1[106], key_s0[106]}), .a ({key_s3[42], key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_2554, new_AGEMA_signal_2553, new_AGEMA_signal_2552, SelectedKey[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_43_U1 ( .s (KeyMUX_n7), .b ({key_s3[107], key_s2[107], key_s1[107], key_s0[107]}), .a ({key_s3[43], key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, new_AGEMA_signal_2561, SelectedKey[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_44_U1 ( .s (KeyMUX_n7), .b ({key_s3[108], key_s2[108], key_s1[108], key_s0[108]}), .a ({key_s3[44], key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_2572, new_AGEMA_signal_2571, new_AGEMA_signal_2570, SelectedKey[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_45_U1 ( .s (KeyMUX_n7), .b ({key_s3[109], key_s2[109], key_s1[109], key_s0[109]}), .a ({key_s3[45], key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_2581, new_AGEMA_signal_2580, new_AGEMA_signal_2579, SelectedKey[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_46_U1 ( .s (KeyMUX_n7), .b ({key_s3[110], key_s2[110], key_s1[110], key_s0[110]}), .a ({key_s3[46], key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_2590, new_AGEMA_signal_2589, new_AGEMA_signal_2588, SelectedKey[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_47_U1 ( .s (KeyMUX_n7), .b ({key_s3[111], key_s2[111], key_s1[111], key_s0[111]}), .a ({key_s3[47], key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_2599, new_AGEMA_signal_2598, new_AGEMA_signal_2597, SelectedKey[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_48_U1 ( .s (KeyMUX_n7), .b ({key_s3[112], key_s2[112], key_s1[112], key_s0[112]}), .a ({key_s3[48], key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, SelectedKey[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_49_U1 ( .s (KeyMUX_n7), .b ({key_s3[113], key_s2[113], key_s1[113], key_s0[113]}), .a ({key_s3[49], key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, new_AGEMA_signal_2615, SelectedKey[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_50_U1 ( .s (KeyMUX_n7), .b ({key_s3[114], key_s2[114], key_s1[114], key_s0[114]}), .a ({key_s3[50], key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, new_AGEMA_signal_2624, SelectedKey[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_51_U1 ( .s (KeyMUX_n7), .b ({key_s3[115], key_s2[115], key_s1[115], key_s0[115]}), .a ({key_s3[51], key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, new_AGEMA_signal_2633, SelectedKey[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_52_U1 ( .s (KeyMUX_n7), .b ({key_s3[116], key_s2[116], key_s1[116], key_s0[116]}), .a ({key_s3[52], key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, SelectedKey[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_53_U1 ( .s (selects[0]), .b ({key_s3[117], key_s2[117], key_s1[117], key_s0[117]}), .a ({key_s3[53], key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, new_AGEMA_signal_1796, SelectedKey[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_54_U1 ( .s (selects[0]), .b ({key_s3[118], key_s2[118], key_s1[118], key_s0[118]}), .a ({key_s3[54], key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, new_AGEMA_signal_1805, SelectedKey[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_55_U1 ( .s (KeyMUX_n7), .b ({key_s3[119], key_s2[119], key_s1[119], key_s0[119]}), .a ({key_s3[55], key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, new_AGEMA_signal_2651, SelectedKey[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_56_U1 ( .s (selects[0]), .b ({key_s3[120], key_s2[120], key_s1[120], key_s0[120]}), .a ({key_s3[56], key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, SelectedKey[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_57_U1 ( .s (KeyMUX_n7), .b ({key_s3[121], key_s2[121], key_s1[121], key_s0[121]}), .a ({key_s3[57], key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, new_AGEMA_signal_2660, SelectedKey[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_58_U1 ( .s (KeyMUX_n7), .b ({key_s3[122], key_s2[122], key_s1[122], key_s0[122]}), .a ({key_s3[58], key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, new_AGEMA_signal_2669, SelectedKey[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_59_U1 ( .s (selects[0]), .b ({key_s3[123], key_s2[123], key_s1[123], key_s0[123]}), .a ({key_s3[59], key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, SelectedKey[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_60_U1 ( .s (KeyMUX_n7), .b ({key_s3[124], key_s2[124], key_s1[124], key_s0[124]}), .a ({key_s3[60], key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, SelectedKey[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_61_U1 ( .s (KeyMUX_n7), .b ({key_s3[125], key_s2[125], key_s1[125], key_s0[125]}), .a ({key_s3[61], key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, SelectedKey[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_62_U1 ( .s (selects[0]), .b ({key_s3[126], key_s2[126], key_s1[126], key_s0[126]}), .a ({key_s3[62], key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, SelectedKey[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyMUX_MUXInst_63_U1 ( .s (KeyMUX_n7), .b ({key_s3[127], key_s2[127], key_s1[127], key_s0[127]}), .a ({key_s3[63], key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, SelectedKey[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMReg[0]), .B (1'b1), .Z (RoundConstant_0) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMReg[1]), .B (1'b0), .Z (FSMUpdate[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMReg[2]), .B (1'b0), .Z (FSMUpdate[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMReg[3]), .B (1'b1), .Z (RoundConstant_4_) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMReg[4]), .B (1'b0), .Z (FSMUpdate[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMReg[5]), .B (1'b0), .Z (FSMUpdate[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_6_U1 ( .S (rst), .A (FSMReg[6]), .B (1'b0), .Z (FSMUpdate[5]) ) ;
    XOR2_X1 FSMUpdateInst_U2 ( .A (RoundConstant_4_), .B (FSMUpdate[3]), .Z (FSMUpdate[6]) ) ;
    XOR2_X1 FSMUpdateInst_U1 ( .A (FSMUpdate[0]), .B (RoundConstant_0), .Z (FSMUpdate[2]) ) ;
    AND2_X1 FSMSignalsInst_U6 ( .A1 (FSMUpdate[5]), .A2 (FSMSignalsInst_n5), .ZN (done_internal) ) ;
    NOR2_X1 FSMSignalsInst_U5 ( .A1 (FSMSignalsInst_n4), .A2 (FSMSignalsInst_n3), .ZN (FSMSignalsInst_n5) ) ;
    NAND2_X1 FSMSignalsInst_U4 ( .A1 (FSMSignalsInst_n2), .A2 (FSMSignalsInst_n1), .ZN (FSMSignalsInst_n3) ) ;
    NOR2_X1 FSMSignalsInst_U3 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMSignalsInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_U2 ( .A1 (FSMUpdate[0]), .A2 (RoundConstant_4_), .ZN (FSMSignalsInst_n2) ) ;
    NAND2_X1 FSMSignalsInst_U1 ( .A1 (RoundConstant_0), .A2 (FSMUpdate[1]), .ZN (FSMSignalsInst_n4) ) ;
    MUX2_X1 selectsMUX_MUXInst_0_U1 ( .S (rst), .A (selectsReg[0]), .B (1'b0), .Z (selects[0]) ) ;
    MUX2_X1 selectsMUX_MUXInst_1_U1 ( .S (rst), .A (selectsReg[1]), .B (1'b0), .Z (selects[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U3 ( .A (selectsUpdateInst_n3), .B (selects[1]), .ZN (selectsNext[1]) ) ;
    XNOR2_X1 selectsUpdateInst_U2 ( .A (selects[0]), .B (1'b0), .ZN (selectsUpdateInst_n3) ) ;
    INV_X1 selectsUpdateInst_U1 ( .A (selects[0]), .ZN (selectsNext[0]) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U14 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U13 ( .a ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n8}), .b ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, SubCellInst_SboxInst_0_n7}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, SubCellInst_SboxInst_0_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U10 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_1042, new_AGEMA_signal_1041, new_AGEMA_signal_1040, SubCellInst_SboxInst_0_n9}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_0_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U9 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, SubCellInst_SboxInst_0_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U5 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_1042, new_AGEMA_signal_1041, new_AGEMA_signal_1040, SubCellInst_SboxInst_0_n9}), .b ({new_AGEMA_signal_1039, new_AGEMA_signal_1038, new_AGEMA_signal_1037, SubCellInst_SboxInst_0_n8}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, SubCellInst_SboxInst_0_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U14 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U13 ( .a ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_1_n8}), .b ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, SubCellInst_SboxInst_1_n7}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, new_AGEMA_signal_1424, SubCellInst_SboxInst_1_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U10 ( .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, new_AGEMA_signal_1064, SubCellInst_SboxInst_1_n9}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_1_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U9 ( .a ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, SubCellInst_SboxInst_1_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U5 ( .a ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .b ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, SubCellInst_SboxInst_1_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, new_AGEMA_signal_1064, SubCellInst_SboxInst_1_n9}), .b ({new_AGEMA_signal_1063, new_AGEMA_signal_1062, new_AGEMA_signal_1061, SubCellInst_SboxInst_1_n8}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, SubCellInst_SboxInst_1_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U14 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, new_AGEMA_signal_1073, SubCellInst_SboxInst_2_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U13 ( .a ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_2_n8}), .b ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, SubCellInst_SboxInst_2_n7}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, SubCellInst_SboxInst_2_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U10 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, SubCellInst_SboxInst_2_n9}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_2_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U9 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, SubCellInst_SboxInst_2_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U5 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_2_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, SubCellInst_SboxInst_2_n9}), .b ({new_AGEMA_signal_1087, new_AGEMA_signal_1086, new_AGEMA_signal_1085, SubCellInst_SboxInst_2_n8}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, SubCellInst_SboxInst_2_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U14 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_3_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U13 ( .a ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_3_n8}), .b ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, SubCellInst_SboxInst_3_n7}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, new_AGEMA_signal_1460, SubCellInst_SboxInst_3_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U10 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, SubCellInst_SboxInst_3_n9}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_3_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U9 ( .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, SubCellInst_SboxInst_3_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U5 ( .a ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .b ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, SubCellInst_SboxInst_3_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, SubCellInst_SboxInst_3_n9}), .b ({new_AGEMA_signal_1111, new_AGEMA_signal_1110, new_AGEMA_signal_1109, SubCellInst_SboxInst_3_n8}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, SubCellInst_SboxInst_3_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U14 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, new_AGEMA_signal_1121, SubCellInst_SboxInst_4_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U13 ( .a ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_4_n8}), .b ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, SubCellInst_SboxInst_4_n7}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_1480, new_AGEMA_signal_1479, new_AGEMA_signal_1478, SubCellInst_SboxInst_4_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U10 ( .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, SubCellInst_SboxInst_4_n9}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, new_AGEMA_signal_1481, SubCellInst_SboxInst_4_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U9 ( .a ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1484, SubCellInst_SboxInst_4_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U5 ( .a ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .b ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_4_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, SubCellInst_SboxInst_4_n9}), .b ({new_AGEMA_signal_1135, new_AGEMA_signal_1134, new_AGEMA_signal_1133, SubCellInst_SboxInst_4_n8}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, SubCellInst_SboxInst_4_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U14 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_5_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U13 ( .a ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_5_n8}), .b ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, SubCellInst_SboxInst_5_n7}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, new_AGEMA_signal_1496, SubCellInst_SboxInst_5_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U10 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, SubCellInst_SboxInst_5_n9}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, SubCellInst_SboxInst_5_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U9 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, SubCellInst_SboxInst_5_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U5 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, SubCellInst_SboxInst_5_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, SubCellInst_SboxInst_5_n9}), .b ({new_AGEMA_signal_1159, new_AGEMA_signal_1158, new_AGEMA_signal_1157, SubCellInst_SboxInst_5_n8}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, new_AGEMA_signal_1508, SubCellInst_SboxInst_5_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U14 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, SubCellInst_SboxInst_6_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U13 ( .a ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_6_n8}), .b ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_6_n7}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, SubCellInst_SboxInst_6_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U10 ( .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, SubCellInst_SboxInst_6_n9}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, new_AGEMA_signal_1517, SubCellInst_SboxInst_6_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U9 ( .a ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, SubCellInst_SboxInst_6_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U5 ( .a ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .b ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_6_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, SubCellInst_SboxInst_6_n9}), .b ({new_AGEMA_signal_1183, new_AGEMA_signal_1182, new_AGEMA_signal_1181, SubCellInst_SboxInst_6_n8}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, SubCellInst_SboxInst_6_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U14 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_7_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U13 ( .a ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_7_n8}), .b ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_7_n7}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, SubCellInst_SboxInst_7_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U10 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, new_AGEMA_signal_1208, SubCellInst_SboxInst_7_n9}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, new_AGEMA_signal_1535, SubCellInst_SboxInst_7_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U9 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, SubCellInst_SboxInst_7_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U5 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, SubCellInst_SboxInst_7_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, new_AGEMA_signal_1208, SubCellInst_SboxInst_7_n9}), .b ({new_AGEMA_signal_1207, new_AGEMA_signal_1206, new_AGEMA_signal_1205, SubCellInst_SboxInst_7_n8}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, SubCellInst_SboxInst_7_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U14 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, new_AGEMA_signal_1217, SubCellInst_SboxInst_8_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U13 ( .a ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_8_n8}), .b ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_8_n7}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, SubCellInst_SboxInst_8_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U10 ( .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, SubCellInst_SboxInst_8_n9}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, new_AGEMA_signal_1553, SubCellInst_SboxInst_8_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U9 ( .a ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, SubCellInst_SboxInst_8_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U5 ( .a ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .b ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_8_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, SubCellInst_SboxInst_8_n9}), .b ({new_AGEMA_signal_1231, new_AGEMA_signal_1230, new_AGEMA_signal_1229, SubCellInst_SboxInst_8_n8}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, SubCellInst_SboxInst_8_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U14 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_9_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U13 ( .a ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_9_n8}), .b ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_9_n7}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, SubCellInst_SboxInst_9_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U10 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, SubCellInst_SboxInst_9_n9}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_9_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U9 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, SubCellInst_SboxInst_9_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U5 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, SubCellInst_SboxInst_9_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, SubCellInst_SboxInst_9_n9}), .b ({new_AGEMA_signal_1255, new_AGEMA_signal_1254, new_AGEMA_signal_1253, SubCellInst_SboxInst_9_n8}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, SubCellInst_SboxInst_9_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U14 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, SubCellInst_SboxInst_10_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U13 ( .a ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_10_n8}), .b ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_10_n7}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, SubCellInst_SboxInst_10_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U10 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, new_AGEMA_signal_1280, SubCellInst_SboxInst_10_n9}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, new_AGEMA_signal_1589, SubCellInst_SboxInst_10_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U9 ( .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, SubCellInst_SboxInst_10_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U5 ( .a ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .b ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_10_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, new_AGEMA_signal_1280, SubCellInst_SboxInst_10_n9}), .b ({new_AGEMA_signal_1279, new_AGEMA_signal_1278, new_AGEMA_signal_1277, SubCellInst_SboxInst_10_n8}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, SubCellInst_SboxInst_10_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U14 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_11_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U13 ( .a ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_11_n8}), .b ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n7}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, SubCellInst_SboxInst_11_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U10 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, SubCellInst_SboxInst_11_n9}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_11_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U9 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, SubCellInst_SboxInst_11_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U5 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_11_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, SubCellInst_SboxInst_11_n9}), .b ({new_AGEMA_signal_1303, new_AGEMA_signal_1302, new_AGEMA_signal_1301, SubCellInst_SboxInst_11_n8}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, SubCellInst_SboxInst_11_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U14 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_12_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U13 ( .a ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_12_n8}), .b ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_12_n7}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, SubCellInst_SboxInst_12_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U10 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, SubCellInst_SboxInst_12_n9}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_12_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U9 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, SubCellInst_SboxInst_12_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U5 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_12_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, SubCellInst_SboxInst_12_n9}), .b ({new_AGEMA_signal_1327, new_AGEMA_signal_1326, new_AGEMA_signal_1325, SubCellInst_SboxInst_12_n8}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, SubCellInst_SboxInst_12_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U14 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_13_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U13 ( .a ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_13_n8}), .b ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_13_n7}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, SubCellInst_SboxInst_13_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U10 ( .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, new_AGEMA_signal_1352, SubCellInst_SboxInst_13_n9}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, new_AGEMA_signal_1643, SubCellInst_SboxInst_13_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U9 ( .a ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, SubCellInst_SboxInst_13_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U5 ( .a ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .b ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_13_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, new_AGEMA_signal_1352, SubCellInst_SboxInst_13_n9}), .b ({new_AGEMA_signal_1351, new_AGEMA_signal_1350, new_AGEMA_signal_1349, SubCellInst_SboxInst_13_n8}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, SubCellInst_SboxInst_13_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U14 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_14_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U13 ( .a ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_14_n8}), .b ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, new_AGEMA_signal_1370, SubCellInst_SboxInst_14_n7}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, SubCellInst_SboxInst_14_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U10 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, SubCellInst_SboxInst_14_n9}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_14_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U9 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, SubCellInst_SboxInst_14_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U5 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_14_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, SubCellInst_SboxInst_14_n9}), .b ({new_AGEMA_signal_1375, new_AGEMA_signal_1374, new_AGEMA_signal_1373, SubCellInst_SboxInst_14_n8}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, SubCellInst_SboxInst_14_n13}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U14 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_15_n10}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U13 ( .a ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_15_n8}), .b ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, SubCellInst_SboxInst_15_n7}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1676, SubCellInst_SboxInst_15_n15}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U10 ( .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, SubCellInst_SboxInst_15_n9}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, SubCellInst_SboxInst_15_n4}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U9 ( .a ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, SubCellInst_SboxInst_15_n6}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U5 ( .a ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .b ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_15_n1}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, SubCellInst_SboxInst_15_n9}), .b ({new_AGEMA_signal_1399, new_AGEMA_signal_1398, new_AGEMA_signal_1397, SubCellInst_SboxInst_15_n8}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, SubCellInst_SboxInst_15_n13}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U18 ( .a ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, SubCellInst_SboxInst_0_n13}), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, SubCellInst_SboxInst_0_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U15 ( .a ({new_AGEMA_signal_1027, new_AGEMA_signal_1026, new_AGEMA_signal_1025, SubCellInst_SboxInst_0_n10}), .b ({new_AGEMA_signal_1042, new_AGEMA_signal_1041, new_AGEMA_signal_1040, SubCellInst_SboxInst_0_n9}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_0_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U11 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_1411, new_AGEMA_signal_1410, new_AGEMA_signal_1409, SubCellInst_SboxInst_0_n4}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_0_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U6 ( .a ({new_AGEMA_signal_1036, new_AGEMA_signal_1035, new_AGEMA_signal_1034, SubCellInst_SboxInst_0_n7}), .b ({new_AGEMA_signal_1033, new_AGEMA_signal_1032, new_AGEMA_signal_1031, SubCellInst_SboxInst_0_n1}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_0_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U18 ( .a ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, SubCellInst_SboxInst_1_n13}), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, new_AGEMA_signal_1853, SubCellInst_SboxInst_1_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U15 ( .a ({new_AGEMA_signal_1051, new_AGEMA_signal_1050, new_AGEMA_signal_1049, SubCellInst_SboxInst_1_n10}), .b ({new_AGEMA_signal_1066, new_AGEMA_signal_1065, new_AGEMA_signal_1064, SubCellInst_SboxInst_1_n9}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_1_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U11 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_1429, new_AGEMA_signal_1428, new_AGEMA_signal_1427, SubCellInst_SboxInst_1_n4}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, SubCellInst_SboxInst_1_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U6 ( .a ({new_AGEMA_signal_1060, new_AGEMA_signal_1059, new_AGEMA_signal_1058, SubCellInst_SboxInst_1_n7}), .b ({new_AGEMA_signal_1057, new_AGEMA_signal_1056, new_AGEMA_signal_1055, SubCellInst_SboxInst_1_n1}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_1_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U18 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, SubCellInst_SboxInst_2_n13}), .b ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_2_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U15 ( .a ({new_AGEMA_signal_1075, new_AGEMA_signal_1074, new_AGEMA_signal_1073, SubCellInst_SboxInst_2_n10}), .b ({new_AGEMA_signal_1090, new_AGEMA_signal_1089, new_AGEMA_signal_1088, SubCellInst_SboxInst_2_n9}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_2_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U11 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_1447, new_AGEMA_signal_1446, new_AGEMA_signal_1445, SubCellInst_SboxInst_2_n4}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, SubCellInst_SboxInst_2_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U6 ( .a ({new_AGEMA_signal_1084, new_AGEMA_signal_1083, new_AGEMA_signal_1082, SubCellInst_SboxInst_2_n7}), .b ({new_AGEMA_signal_1081, new_AGEMA_signal_1080, new_AGEMA_signal_1079, SubCellInst_SboxInst_2_n1}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_2_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U18 ( .a ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, SubCellInst_SboxInst_3_n13}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, new_AGEMA_signal_1883, SubCellInst_SboxInst_3_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U15 ( .a ({new_AGEMA_signal_1099, new_AGEMA_signal_1098, new_AGEMA_signal_1097, SubCellInst_SboxInst_3_n10}), .b ({new_AGEMA_signal_1114, new_AGEMA_signal_1113, new_AGEMA_signal_1112, SubCellInst_SboxInst_3_n9}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_3_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U11 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_1465, new_AGEMA_signal_1464, new_AGEMA_signal_1463, SubCellInst_SboxInst_3_n4}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1889, SubCellInst_SboxInst_3_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U6 ( .a ({new_AGEMA_signal_1108, new_AGEMA_signal_1107, new_AGEMA_signal_1106, SubCellInst_SboxInst_3_n7}), .b ({new_AGEMA_signal_1105, new_AGEMA_signal_1104, new_AGEMA_signal_1103, SubCellInst_SboxInst_3_n1}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, new_AGEMA_signal_1469, SubCellInst_SboxInst_3_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U18 ( .a ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, SubCellInst_SboxInst_4_n13}), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1898, SubCellInst_SboxInst_4_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U15 ( .a ({new_AGEMA_signal_1123, new_AGEMA_signal_1122, new_AGEMA_signal_1121, SubCellInst_SboxInst_4_n10}), .b ({new_AGEMA_signal_1138, new_AGEMA_signal_1137, new_AGEMA_signal_1136, SubCellInst_SboxInst_4_n9}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, SubCellInst_SboxInst_4_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U11 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_1483, new_AGEMA_signal_1482, new_AGEMA_signal_1481, SubCellInst_SboxInst_4_n4}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_4_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U6 ( .a ({new_AGEMA_signal_1132, new_AGEMA_signal_1131, new_AGEMA_signal_1130, SubCellInst_SboxInst_4_n7}), .b ({new_AGEMA_signal_1129, new_AGEMA_signal_1128, new_AGEMA_signal_1127, SubCellInst_SboxInst_4_n1}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1487, SubCellInst_SboxInst_4_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U18 ( .a ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, new_AGEMA_signal_1508, SubCellInst_SboxInst_5_n13}), .b ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, new_AGEMA_signal_1913, SubCellInst_SboxInst_5_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U15 ( .a ({new_AGEMA_signal_1147, new_AGEMA_signal_1146, new_AGEMA_signal_1145, SubCellInst_SboxInst_5_n10}), .b ({new_AGEMA_signal_1162, new_AGEMA_signal_1161, new_AGEMA_signal_1160, SubCellInst_SboxInst_5_n9}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, new_AGEMA_signal_1493, SubCellInst_SboxInst_5_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U11 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_1501, new_AGEMA_signal_1500, new_AGEMA_signal_1499, SubCellInst_SboxInst_5_n4}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, SubCellInst_SboxInst_5_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U6 ( .a ({new_AGEMA_signal_1156, new_AGEMA_signal_1155, new_AGEMA_signal_1154, SubCellInst_SboxInst_5_n7}), .b ({new_AGEMA_signal_1153, new_AGEMA_signal_1152, new_AGEMA_signal_1151, SubCellInst_SboxInst_5_n1}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1505, SubCellInst_SboxInst_5_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U18 ( .a ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, SubCellInst_SboxInst_6_n13}), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_6_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U15 ( .a ({new_AGEMA_signal_1171, new_AGEMA_signal_1170, new_AGEMA_signal_1169, SubCellInst_SboxInst_6_n10}), .b ({new_AGEMA_signal_1186, new_AGEMA_signal_1185, new_AGEMA_signal_1184, SubCellInst_SboxInst_6_n9}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, SubCellInst_SboxInst_6_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U11 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1518, new_AGEMA_signal_1517, SubCellInst_SboxInst_6_n4}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_6_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U6 ( .a ({new_AGEMA_signal_1180, new_AGEMA_signal_1179, new_AGEMA_signal_1178, SubCellInst_SboxInst_6_n7}), .b ({new_AGEMA_signal_1177, new_AGEMA_signal_1176, new_AGEMA_signal_1175, SubCellInst_SboxInst_6_n1}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, SubCellInst_SboxInst_6_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U18 ( .a ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, SubCellInst_SboxInst_7_n13}), .b ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, SubCellInst_SboxInst_7_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U15 ( .a ({new_AGEMA_signal_1195, new_AGEMA_signal_1194, new_AGEMA_signal_1193, SubCellInst_SboxInst_7_n10}), .b ({new_AGEMA_signal_1210, new_AGEMA_signal_1209, new_AGEMA_signal_1208, SubCellInst_SboxInst_7_n9}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1529, SubCellInst_SboxInst_7_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U11 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_1537, new_AGEMA_signal_1536, new_AGEMA_signal_1535, SubCellInst_SboxInst_7_n4}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, new_AGEMA_signal_1949, SubCellInst_SboxInst_7_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U6 ( .a ({new_AGEMA_signal_1204, new_AGEMA_signal_1203, new_AGEMA_signal_1202, SubCellInst_SboxInst_7_n7}), .b ({new_AGEMA_signal_1201, new_AGEMA_signal_1200, new_AGEMA_signal_1199, SubCellInst_SboxInst_7_n1}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1541, SubCellInst_SboxInst_7_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U18 ( .a ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, SubCellInst_SboxInst_8_n13}), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_8_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U15 ( .a ({new_AGEMA_signal_1219, new_AGEMA_signal_1218, new_AGEMA_signal_1217, SubCellInst_SboxInst_8_n10}), .b ({new_AGEMA_signal_1234, new_AGEMA_signal_1233, new_AGEMA_signal_1232, SubCellInst_SboxInst_8_n9}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, SubCellInst_SboxInst_8_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U11 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_1555, new_AGEMA_signal_1554, new_AGEMA_signal_1553, SubCellInst_SboxInst_8_n4}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_8_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U6 ( .a ({new_AGEMA_signal_1228, new_AGEMA_signal_1227, new_AGEMA_signal_1226, SubCellInst_SboxInst_8_n7}), .b ({new_AGEMA_signal_1225, new_AGEMA_signal_1224, new_AGEMA_signal_1223, SubCellInst_SboxInst_8_n1}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1559, SubCellInst_SboxInst_8_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U18 ( .a ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, SubCellInst_SboxInst_9_n13}), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, new_AGEMA_signal_1973, SubCellInst_SboxInst_9_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U15 ( .a ({new_AGEMA_signal_1243, new_AGEMA_signal_1242, new_AGEMA_signal_1241, SubCellInst_SboxInst_9_n10}), .b ({new_AGEMA_signal_1258, new_AGEMA_signal_1257, new_AGEMA_signal_1256, SubCellInst_SboxInst_9_n9}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1565, SubCellInst_SboxInst_9_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U11 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_1573, new_AGEMA_signal_1572, new_AGEMA_signal_1571, SubCellInst_SboxInst_9_n4}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, SubCellInst_SboxInst_9_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U6 ( .a ({new_AGEMA_signal_1252, new_AGEMA_signal_1251, new_AGEMA_signal_1250, SubCellInst_SboxInst_9_n7}), .b ({new_AGEMA_signal_1249, new_AGEMA_signal_1248, new_AGEMA_signal_1247, SubCellInst_SboxInst_9_n1}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_9_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U18 ( .a ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, SubCellInst_SboxInst_10_n13}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_10_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U15 ( .a ({new_AGEMA_signal_1267, new_AGEMA_signal_1266, new_AGEMA_signal_1265, SubCellInst_SboxInst_10_n10}), .b ({new_AGEMA_signal_1282, new_AGEMA_signal_1281, new_AGEMA_signal_1280, SubCellInst_SboxInst_10_n9}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, SubCellInst_SboxInst_10_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U11 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_1591, new_AGEMA_signal_1590, new_AGEMA_signal_1589, SubCellInst_SboxInst_10_n4}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U6 ( .a ({new_AGEMA_signal_1276, new_AGEMA_signal_1275, new_AGEMA_signal_1274, SubCellInst_SboxInst_10_n7}), .b ({new_AGEMA_signal_1273, new_AGEMA_signal_1272, new_AGEMA_signal_1271, SubCellInst_SboxInst_10_n1}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_10_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U18 ( .a ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, SubCellInst_SboxInst_11_n13}), .b ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, SubCellInst_SboxInst_11_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U15 ( .a ({new_AGEMA_signal_1291, new_AGEMA_signal_1290, new_AGEMA_signal_1289, SubCellInst_SboxInst_11_n10}), .b ({new_AGEMA_signal_1306, new_AGEMA_signal_1305, new_AGEMA_signal_1304, SubCellInst_SboxInst_11_n9}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_11_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U11 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_1609, new_AGEMA_signal_1608, new_AGEMA_signal_1607, SubCellInst_SboxInst_11_n4}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, SubCellInst_SboxInst_11_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U6 ( .a ({new_AGEMA_signal_1300, new_AGEMA_signal_1299, new_AGEMA_signal_1298, SubCellInst_SboxInst_11_n7}), .b ({new_AGEMA_signal_1297, new_AGEMA_signal_1296, new_AGEMA_signal_1295, SubCellInst_SboxInst_11_n1}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1613, SubCellInst_SboxInst_11_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U18 ( .a ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, SubCellInst_SboxInst_12_n13}), .b ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_12_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U15 ( .a ({new_AGEMA_signal_1315, new_AGEMA_signal_1314, new_AGEMA_signal_1313, SubCellInst_SboxInst_12_n10}), .b ({new_AGEMA_signal_1330, new_AGEMA_signal_1329, new_AGEMA_signal_1328, SubCellInst_SboxInst_12_n9}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, SubCellInst_SboxInst_12_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U11 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_1627, new_AGEMA_signal_1626, new_AGEMA_signal_1625, SubCellInst_SboxInst_12_n4}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_12_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U6 ( .a ({new_AGEMA_signal_1324, new_AGEMA_signal_1323, new_AGEMA_signal_1322, SubCellInst_SboxInst_12_n7}), .b ({new_AGEMA_signal_1321, new_AGEMA_signal_1320, new_AGEMA_signal_1319, SubCellInst_SboxInst_12_n1}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_12_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U18 ( .a ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, SubCellInst_SboxInst_13_n13}), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, SubCellInst_SboxInst_13_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U15 ( .a ({new_AGEMA_signal_1339, new_AGEMA_signal_1338, new_AGEMA_signal_1337, SubCellInst_SboxInst_13_n10}), .b ({new_AGEMA_signal_1354, new_AGEMA_signal_1353, new_AGEMA_signal_1352, SubCellInst_SboxInst_13_n9}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_13_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U11 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_1645, new_AGEMA_signal_1644, new_AGEMA_signal_1643, SubCellInst_SboxInst_13_n4}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, SubCellInst_SboxInst_13_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U6 ( .a ({new_AGEMA_signal_1348, new_AGEMA_signal_1347, new_AGEMA_signal_1346, SubCellInst_SboxInst_13_n7}), .b ({new_AGEMA_signal_1345, new_AGEMA_signal_1344, new_AGEMA_signal_1343, SubCellInst_SboxInst_13_n1}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1649, SubCellInst_SboxInst_13_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U18 ( .a ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, SubCellInst_SboxInst_14_n13}), .b ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, SubCellInst_SboxInst_14_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U15 ( .a ({new_AGEMA_signal_1363, new_AGEMA_signal_1362, new_AGEMA_signal_1361, SubCellInst_SboxInst_14_n10}), .b ({new_AGEMA_signal_1378, new_AGEMA_signal_1377, new_AGEMA_signal_1376, SubCellInst_SboxInst_14_n9}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_14_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U11 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_1663, new_AGEMA_signal_1662, new_AGEMA_signal_1661, SubCellInst_SboxInst_14_n4}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, SubCellInst_SboxInst_14_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U6 ( .a ({new_AGEMA_signal_1372, new_AGEMA_signal_1371, new_AGEMA_signal_1370, SubCellInst_SboxInst_14_n7}), .b ({new_AGEMA_signal_1369, new_AGEMA_signal_1368, new_AGEMA_signal_1367, SubCellInst_SboxInst_14_n1}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_14_n2}) ) ;
    or_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U18 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, SubCellInst_SboxInst_15_n13}), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, SubCellInst_SboxInst_15_n14}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U15 ( .a ({new_AGEMA_signal_1387, new_AGEMA_signal_1386, new_AGEMA_signal_1385, SubCellInst_SboxInst_15_n10}), .b ({new_AGEMA_signal_1402, new_AGEMA_signal_1401, new_AGEMA_signal_1400, SubCellInst_SboxInst_15_n9}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1673, SubCellInst_SboxInst_15_n11}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U11 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_1681, new_AGEMA_signal_1680, new_AGEMA_signal_1679, SubCellInst_SboxInst_15_n4}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, SubCellInst_SboxInst_15_n5}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U6 ( .a ({new_AGEMA_signal_1396, new_AGEMA_signal_1395, new_AGEMA_signal_1394, SubCellInst_SboxInst_15_n7}), .b ({new_AGEMA_signal_1393, new_AGEMA_signal_1392, new_AGEMA_signal_1391, SubCellInst_SboxInst_15_n1}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_15_n2}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, Feedback[1]}), .a ({plaintext_s3[1], plaintext_s2[1], plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, MCOutput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, Feedback[3]}), .a ({plaintext_s3[3], plaintext_s2[3], plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, MCOutput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, Feedback[5]}), .a ({plaintext_s3[5], plaintext_s2[5], plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, new_AGEMA_signal_2732, MCOutput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, Feedback[7]}), .a ({plaintext_s3[7], plaintext_s2[7], plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, new_AGEMA_signal_2105, Feedback[9]}), .a ({plaintext_s3[9], plaintext_s2[9], plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, Feedback[11]}), .a ({plaintext_s3[11], plaintext_s2[11], plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCOutput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, Feedback[13]}), .a ({plaintext_s3[13], plaintext_s2[13], plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCOutput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, new_AGEMA_signal_2111, Feedback[15]}), .a ({plaintext_s3[15], plaintext_s2[15], plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCOutput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, Feedback[17]}), .a ({plaintext_s3[17], plaintext_s2[17], plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, new_AGEMA_signal_2804, MCOutput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, Feedback[19]}), .a ({plaintext_s3[19], plaintext_s2[19], plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, MCOutput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, new_AGEMA_signal_2141, Feedback[21]}), .a ({plaintext_s3[21], plaintext_s2[21], plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, MCOutput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, Feedback[23]}), .a ({plaintext_s3[23], plaintext_s2[23], plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, MCOutput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, Feedback[25]}), .a ({plaintext_s3[25], plaintext_s2[25], plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, MCOutput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, Feedback[27]}), .a ({plaintext_s3[27], plaintext_s2[27], plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCOutput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, new_AGEMA_signal_2165, Feedback[29]}), .a ({plaintext_s3[29], plaintext_s2[29], plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCOutput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, Feedback[31]}), .a ({plaintext_s3[31], plaintext_s2[31], plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCOutput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, Feedback[33]}), .a ({plaintext_s3[33], plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, MCInput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, Feedback[35]}), .a ({plaintext_s3[35], plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_2914, new_AGEMA_signal_2913, new_AGEMA_signal_2912, MCInput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, Feedback[37]}), .a ({plaintext_s3[37], plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_2926, new_AGEMA_signal_2925, new_AGEMA_signal_2924, MCInput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, Feedback[39]}), .a ({plaintext_s3[39], plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_2938, new_AGEMA_signal_2937, new_AGEMA_signal_2936, MCInput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, new_AGEMA_signal_2201, Feedback[41]}), .a ({plaintext_s3[41], plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_2950, new_AGEMA_signal_2949, new_AGEMA_signal_2948, MCInput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, Feedback[43]}), .a ({plaintext_s3[43], plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_2962, new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCInput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, Feedback[45]}), .a ({plaintext_s3[45], plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, new_AGEMA_signal_2972, MCInput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, Feedback[47]}), .a ({plaintext_s3[47], plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, new_AGEMA_signal_2984, MCInput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, new_AGEMA_signal_2225, Feedback[49]}), .a ({plaintext_s3[49], plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, new_AGEMA_signal_2996, MCInput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, Feedback[51]}), .a ({plaintext_s3[51], plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, MCInput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, Feedback[53]}), .a ({plaintext_s3[53], plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, new_AGEMA_signal_3020, MCInput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, Feedback[55]}), .a ({plaintext_s3[55], plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, new_AGEMA_signal_3032, MCInput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, Feedback[57]}), .a ({plaintext_s3[57], plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, new_AGEMA_signal_3044, MCInput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, Feedback[59]}), .a ({plaintext_s3[59], plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, new_AGEMA_signal_3056, MCInput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, new_AGEMA_signal_2261, Feedback[61]}), .a ({plaintext_s3[61], plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_3070, new_AGEMA_signal_3069, new_AGEMA_signal_3068, MCInput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, Feedback[63]}), .a ({plaintext_s3[63], plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, MCInput[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_1_U3 ( .a ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, new_AGEMA_signal_3119, MCInst_XOR_r0_Inst_1_n2}), .b ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, MCInst_XOR_r0_Inst_1_n1}), .c ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, new_AGEMA_signal_3353, MCOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_1_U2 ( .a ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, new_AGEMA_signal_2804, MCOutput[17]}), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, MCOutput[1]}), .c ({new_AGEMA_signal_3118, new_AGEMA_signal_3117, new_AGEMA_signal_3116, MCInst_XOR_r0_Inst_1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2998, new_AGEMA_signal_2997, new_AGEMA_signal_2996, MCInput[49]}), .c ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, new_AGEMA_signal_3119, MCInst_XOR_r0_Inst_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_1_U2 ( .a ({new_AGEMA_signal_3124, new_AGEMA_signal_3123, new_AGEMA_signal_3122, MCInst_XOR_r1_Inst_1_n1}), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, MCOutput[1]}), .c ({new_AGEMA_signal_3358, new_AGEMA_signal_3357, new_AGEMA_signal_3356, MCOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2902, new_AGEMA_signal_2901, new_AGEMA_signal_2900, MCInput[33]}), .c ({new_AGEMA_signal_3124, new_AGEMA_signal_3123, new_AGEMA_signal_3122, MCInst_XOR_r1_Inst_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_3_U3 ( .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, new_AGEMA_signal_3137, MCInst_XOR_r0_Inst_3_n2}), .b ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, MCInst_XOR_r0_Inst_3_n1}), .c ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, new_AGEMA_signal_3365, MCOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_3_U2 ( .a ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, MCOutput[19]}), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, MCOutput[3]}), .c ({new_AGEMA_signal_3136, new_AGEMA_signal_3135, new_AGEMA_signal_3134, MCInst_XOR_r0_Inst_3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3010, new_AGEMA_signal_3009, new_AGEMA_signal_3008, MCInput[51]}), .c ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, new_AGEMA_signal_3137, MCInst_XOR_r0_Inst_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_3_U2 ( .a ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, new_AGEMA_signal_3140, MCInst_XOR_r1_Inst_3_n1}), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, MCOutput[3]}), .c ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, new_AGEMA_signal_3368, MCOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2914, new_AGEMA_signal_2913, new_AGEMA_signal_2912, MCInput[35]}), .c ({new_AGEMA_signal_3142, new_AGEMA_signal_3141, new_AGEMA_signal_3140, MCInst_XOR_r1_Inst_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_5_U3 ( .a ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, new_AGEMA_signal_3155, MCInst_XOR_r0_Inst_5_n2}), .b ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, new_AGEMA_signal_3152, MCInst_XOR_r0_Inst_5_n1}), .c ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, new_AGEMA_signal_3377, MCOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_5_U2 ( .a ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, MCOutput[21]}), .b ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, new_AGEMA_signal_2732, MCOutput[5]}), .c ({new_AGEMA_signal_3154, new_AGEMA_signal_3153, new_AGEMA_signal_3152, MCInst_XOR_r0_Inst_5_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_5_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3022, new_AGEMA_signal_3021, new_AGEMA_signal_3020, MCInput[53]}), .c ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, new_AGEMA_signal_3155, MCInst_XOR_r0_Inst_5_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_5_U2 ( .a ({new_AGEMA_signal_3160, new_AGEMA_signal_3159, new_AGEMA_signal_3158, MCInst_XOR_r1_Inst_5_n1}), .b ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, new_AGEMA_signal_2732, MCOutput[5]}), .c ({new_AGEMA_signal_3382, new_AGEMA_signal_3381, new_AGEMA_signal_3380, MCOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_5_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2926, new_AGEMA_signal_2925, new_AGEMA_signal_2924, MCInput[37]}), .c ({new_AGEMA_signal_3160, new_AGEMA_signal_3159, new_AGEMA_signal_3158, MCInst_XOR_r1_Inst_5_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_7_U3 ( .a ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, new_AGEMA_signal_3173, MCInst_XOR_r0_Inst_7_n2}), .b ({new_AGEMA_signal_3172, new_AGEMA_signal_3171, new_AGEMA_signal_3170, MCInst_XOR_r0_Inst_7_n1}), .c ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, new_AGEMA_signal_3389, MCOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_7_U2 ( .a ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, MCOutput[23]}), .b ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[7]}), .c ({new_AGEMA_signal_3172, new_AGEMA_signal_3171, new_AGEMA_signal_3170, MCInst_XOR_r0_Inst_7_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_7_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3034, new_AGEMA_signal_3033, new_AGEMA_signal_3032, MCInput[55]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, new_AGEMA_signal_3173, MCInst_XOR_r0_Inst_7_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_7_U2 ( .a ({new_AGEMA_signal_3178, new_AGEMA_signal_3177, new_AGEMA_signal_3176, MCInst_XOR_r1_Inst_7_n1}), .b ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[7]}), .c ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, MCOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_7_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2938, new_AGEMA_signal_2937, new_AGEMA_signal_2936, MCInput[39]}), .c ({new_AGEMA_signal_3178, new_AGEMA_signal_3177, new_AGEMA_signal_3176, MCInst_XOR_r1_Inst_7_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_9_U3 ( .a ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, new_AGEMA_signal_3191, MCInst_XOR_r0_Inst_9_n2}), .b ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, new_AGEMA_signal_3188, MCInst_XOR_r0_Inst_9_n1}), .c ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, MCOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_9_U2 ( .a ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, MCOutput[25]}), .b ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[9]}), .c ({new_AGEMA_signal_3190, new_AGEMA_signal_3189, new_AGEMA_signal_3188, MCInst_XOR_r0_Inst_9_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_9_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3046, new_AGEMA_signal_3045, new_AGEMA_signal_3044, MCInput[57]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, new_AGEMA_signal_3191, MCInst_XOR_r0_Inst_9_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_9_U2 ( .a ({new_AGEMA_signal_3196, new_AGEMA_signal_3195, new_AGEMA_signal_3194, MCInst_XOR_r1_Inst_9_n1}), .b ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[9]}), .c ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, new_AGEMA_signal_3404, MCOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_9_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2950, new_AGEMA_signal_2949, new_AGEMA_signal_2948, MCInput[41]}), .c ({new_AGEMA_signal_3196, new_AGEMA_signal_3195, new_AGEMA_signal_3194, MCInst_XOR_r1_Inst_9_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_11_U3 ( .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, new_AGEMA_signal_3209, MCInst_XOR_r0_Inst_11_n2}), .b ({new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, MCInst_XOR_r0_Inst_11_n1}), .c ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, new_AGEMA_signal_3413, MCOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_11_U2 ( .a ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCOutput[27]}), .b ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCOutput[11]}), .c ({new_AGEMA_signal_3208, new_AGEMA_signal_3207, new_AGEMA_signal_3206, MCInst_XOR_r0_Inst_11_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_11_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3058, new_AGEMA_signal_3057, new_AGEMA_signal_3056, MCInput[59]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, new_AGEMA_signal_3209, MCInst_XOR_r0_Inst_11_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_11_U2 ( .a ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, new_AGEMA_signal_3212, MCInst_XOR_r1_Inst_11_n1}), .b ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCOutput[11]}), .c ({new_AGEMA_signal_3418, new_AGEMA_signal_3417, new_AGEMA_signal_3416, MCOutput[43]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_11_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2962, new_AGEMA_signal_2961, new_AGEMA_signal_2960, MCInput[43]}), .c ({new_AGEMA_signal_3214, new_AGEMA_signal_3213, new_AGEMA_signal_3212, MCInst_XOR_r1_Inst_11_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_13_U3 ( .a ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, new_AGEMA_signal_3227, MCInst_XOR_r0_Inst_13_n2}), .b ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_3224, MCInst_XOR_r0_Inst_13_n1}), .c ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, new_AGEMA_signal_3425, MCOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_13_U2 ( .a ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCOutput[29]}), .b ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCOutput[13]}), .c ({new_AGEMA_signal_3226, new_AGEMA_signal_3225, new_AGEMA_signal_3224, MCInst_XOR_r0_Inst_13_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_13_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3070, new_AGEMA_signal_3069, new_AGEMA_signal_3068, MCInput[61]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, new_AGEMA_signal_3227, MCInst_XOR_r0_Inst_13_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_13_U2 ( .a ({new_AGEMA_signal_3232, new_AGEMA_signal_3231, new_AGEMA_signal_3230, MCInst_XOR_r1_Inst_13_n1}), .b ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCOutput[13]}), .c ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, MCOutput[45]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_13_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2974, new_AGEMA_signal_2973, new_AGEMA_signal_2972, MCInput[45]}), .c ({new_AGEMA_signal_3232, new_AGEMA_signal_3231, new_AGEMA_signal_3230, MCInst_XOR_r1_Inst_13_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_15_U3 ( .a ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, new_AGEMA_signal_3245, MCInst_XOR_r0_Inst_15_n2}), .b ({new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, MCInst_XOR_r0_Inst_15_n1}), .c ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, MCOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_15_U2 ( .a ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCOutput[31]}), .b ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCOutput[15]}), .c ({new_AGEMA_signal_3244, new_AGEMA_signal_3243, new_AGEMA_signal_3242, MCInst_XOR_r0_Inst_15_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_15_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3082, new_AGEMA_signal_3081, new_AGEMA_signal_3080, MCInput[63]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, new_AGEMA_signal_3245, MCInst_XOR_r0_Inst_15_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_15_U2 ( .a ({new_AGEMA_signal_3250, new_AGEMA_signal_3249, new_AGEMA_signal_3248, MCInst_XOR_r1_Inst_15_n1}), .b ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCOutput[15]}), .c ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, MCOutput[47]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_15_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2986, new_AGEMA_signal_2985, new_AGEMA_signal_2984, MCInput[47]}), .c ({new_AGEMA_signal_3250, new_AGEMA_signal_3249, new_AGEMA_signal_3248, MCInst_XOR_r1_Inst_15_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3544, new_AGEMA_signal_3543, new_AGEMA_signal_3542, AddKeyXOR1_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2617, new_AGEMA_signal_2616, new_AGEMA_signal_2615, SelectedKey[49]}), .c ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, new_AGEMA_signal_3638, AddRoundKeyOutput[49]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, new_AGEMA_signal_3353, MCOutput[49]}), .c ({new_AGEMA_signal_3544, new_AGEMA_signal_3543, new_AGEMA_signal_3542, AddKeyXOR1_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, new_AGEMA_signal_3548, AddKeyXOR1_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, new_AGEMA_signal_2633, SelectedKey[51]}), .c ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, new_AGEMA_signal_3644, AddRoundKeyOutput[51]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, new_AGEMA_signal_3365, MCOutput[51]}), .c ({new_AGEMA_signal_3550, new_AGEMA_signal_3549, new_AGEMA_signal_3548, AddKeyXOR1_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, AddKeyXOR1_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1798, new_AGEMA_signal_1797, new_AGEMA_signal_1796, SelectedKey[53]}), .c ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, new_AGEMA_signal_3650, AddRoundKeyOutput[53]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, new_AGEMA_signal_3377, MCOutput[53]}), .c ({new_AGEMA_signal_3556, new_AGEMA_signal_3555, new_AGEMA_signal_3554, AddKeyXOR1_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3562, new_AGEMA_signal_3561, new_AGEMA_signal_3560, AddKeyXOR1_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, new_AGEMA_signal_2651, SelectedKey[55]}), .c ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, new_AGEMA_signal_3656, AddRoundKeyOutput[55]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, new_AGEMA_signal_3389, MCOutput[55]}), .c ({new_AGEMA_signal_3562, new_AGEMA_signal_3561, new_AGEMA_signal_3560, AddKeyXOR1_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, new_AGEMA_signal_3566, AddKeyXOR1_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2662, new_AGEMA_signal_2661, new_AGEMA_signal_2660, SelectedKey[57]}), .c ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, AddRoundKeyOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, new_AGEMA_signal_3401, MCOutput[57]}), .c ({new_AGEMA_signal_3568, new_AGEMA_signal_3567, new_AGEMA_signal_3566, AddKeyXOR1_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, new_AGEMA_signal_3572, AddKeyXOR1_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1825, new_AGEMA_signal_1824, new_AGEMA_signal_1823, SelectedKey[59]}), .c ({new_AGEMA_signal_3670, new_AGEMA_signal_3669, new_AGEMA_signal_3668, AddRoundKeyOutput[59]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, new_AGEMA_signal_3413, MCOutput[59]}), .c ({new_AGEMA_signal_3574, new_AGEMA_signal_3573, new_AGEMA_signal_3572, AddKeyXOR1_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3580, new_AGEMA_signal_3579, new_AGEMA_signal_3578, AddKeyXOR1_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, new_AGEMA_signal_2687, SelectedKey[61]}), .c ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, new_AGEMA_signal_3674, AddRoundKeyOutput[61]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, new_AGEMA_signal_3425, MCOutput[61]}), .c ({new_AGEMA_signal_3580, new_AGEMA_signal_3579, new_AGEMA_signal_3578, AddKeyXOR1_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, new_AGEMA_signal_3584, AddKeyXOR1_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2698, new_AGEMA_signal_2697, new_AGEMA_signal_2696, SelectedKey[63]}), .c ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, new_AGEMA_signal_3680, AddRoundKeyOutput[63]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, new_AGEMA_signal_3437, MCOutput[63]}), .c ({new_AGEMA_signal_3586, new_AGEMA_signal_3585, new_AGEMA_signal_3584, AddKeyXOR1_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, AddKeyConstXOR_XORInst_0_1_n2}), .b ({new_AGEMA_signal_3088, new_AGEMA_signal_3087, new_AGEMA_signal_3086, AddKeyConstXOR_XORInst_0_1_n1}), .c ({new_AGEMA_signal_3688, new_AGEMA_signal_3687, new_AGEMA_signal_3686, AddRoundKeyOutput[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3406, new_AGEMA_signal_3405, new_AGEMA_signal_3404, MCOutput[41]}), .c ({new_AGEMA_signal_3592, new_AGEMA_signal_3591, new_AGEMA_signal_3590, AddKeyConstXOR_XORInst_0_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_3598, new_AGEMA_signal_3597, new_AGEMA_signal_3596, AddKeyConstXOR_XORInst_0_3_n2}), .b ({new_AGEMA_signal_3094, new_AGEMA_signal_3093, new_AGEMA_signal_3092, AddKeyConstXOR_XORInst_0_3_n1}), .c ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, new_AGEMA_signal_3692, AddRoundKeyOutput[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3418, new_AGEMA_signal_3417, new_AGEMA_signal_3416, MCOutput[43]}), .c ({new_AGEMA_signal_3598, new_AGEMA_signal_3597, new_AGEMA_signal_3596, AddKeyConstXOR_XORInst_0_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, AddKeyConstXOR_XORInst_1_1_n2}), .b ({new_AGEMA_signal_3100, new_AGEMA_signal_3099, new_AGEMA_signal_3098, AddKeyConstXOR_XORInst_1_1_n1}), .c ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, AddRoundKeyOutput[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3430, new_AGEMA_signal_3429, new_AGEMA_signal_3428, MCOutput[45]}), .c ({new_AGEMA_signal_3604, new_AGEMA_signal_3603, new_AGEMA_signal_3602, AddKeyConstXOR_XORInst_1_1_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, AddKeyConstXOR_XORInst_1_3_n2}), .b ({new_AGEMA_signal_3106, new_AGEMA_signal_3105, new_AGEMA_signal_3104, AddKeyConstXOR_XORInst_1_3_n1}), .c ({new_AGEMA_signal_3706, new_AGEMA_signal_3705, new_AGEMA_signal_3704, AddRoundKeyOutput[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3442, new_AGEMA_signal_3441, new_AGEMA_signal_3440, MCOutput[47]}), .c ({new_AGEMA_signal_3610, new_AGEMA_signal_3609, new_AGEMA_signal_3608, AddKeyConstXOR_XORInst_1_3_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3256, new_AGEMA_signal_3255, new_AGEMA_signal_3254, AddKeyXOR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, new_AGEMA_signal_2273, SelectedKey[1]}), .c ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, AddRoundKeyOutput[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2710, new_AGEMA_signal_2709, new_AGEMA_signal_2708, MCOutput[1]}), .c ({new_AGEMA_signal_3256, new_AGEMA_signal_3255, new_AGEMA_signal_3254, AddKeyXOR2_XORInst_0_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, new_AGEMA_signal_3260, AddKeyXOR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2284, new_AGEMA_signal_2283, new_AGEMA_signal_2282, SelectedKey[3]}), .c ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, new_AGEMA_signal_3452, AddRoundKeyOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2722, new_AGEMA_signal_2721, new_AGEMA_signal_2720, MCOutput[3]}), .c ({new_AGEMA_signal_3262, new_AGEMA_signal_3261, new_AGEMA_signal_3260, AddKeyXOR2_XORInst_0_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3268, new_AGEMA_signal_3267, new_AGEMA_signal_3266, AddKeyXOR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_2302, new_AGEMA_signal_2301, new_AGEMA_signal_2300, SelectedKey[5]}), .c ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, AddRoundKeyOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2734, new_AGEMA_signal_2733, new_AGEMA_signal_2732, MCOutput[5]}), .c ({new_AGEMA_signal_3268, new_AGEMA_signal_3267, new_AGEMA_signal_3266, AddKeyXOR2_XORInst_1_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3274, new_AGEMA_signal_3273, new_AGEMA_signal_3272, AddKeyXOR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2320, new_AGEMA_signal_2319, new_AGEMA_signal_2318, SelectedKey[7]}), .c ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, AddRoundKeyOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2746, new_AGEMA_signal_2745, new_AGEMA_signal_2744, MCOutput[7]}), .c ({new_AGEMA_signal_3274, new_AGEMA_signal_3273, new_AGEMA_signal_3272, AddKeyXOR2_XORInst_1_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3280, new_AGEMA_signal_3279, new_AGEMA_signal_3278, AddKeyXOR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_2338, new_AGEMA_signal_2337, new_AGEMA_signal_2336, SelectedKey[9]}), .c ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, new_AGEMA_signal_3470, AddRoundKeyOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2758, new_AGEMA_signal_2757, new_AGEMA_signal_2756, MCOutput[9]}), .c ({new_AGEMA_signal_3280, new_AGEMA_signal_3279, new_AGEMA_signal_3278, AddKeyXOR2_XORInst_2_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, new_AGEMA_signal_3284, AddKeyXOR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2356, new_AGEMA_signal_2355, new_AGEMA_signal_2354, SelectedKey[11]}), .c ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, new_AGEMA_signal_3476, AddRoundKeyOutput[11]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2770, new_AGEMA_signal_2769, new_AGEMA_signal_2768, MCOutput[11]}), .c ({new_AGEMA_signal_3286, new_AGEMA_signal_3285, new_AGEMA_signal_3284, AddKeyXOR2_XORInst_2_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, AddKeyXOR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_2374, new_AGEMA_signal_2373, new_AGEMA_signal_2372, SelectedKey[13]}), .c ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, AddRoundKeyOutput[13]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2782, new_AGEMA_signal_2781, new_AGEMA_signal_2780, MCOutput[13]}), .c ({new_AGEMA_signal_3292, new_AGEMA_signal_3291, new_AGEMA_signal_3290, AddKeyXOR2_XORInst_3_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, new_AGEMA_signal_3296, AddKeyXOR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2392, new_AGEMA_signal_2391, new_AGEMA_signal_2390, SelectedKey[15]}), .c ({new_AGEMA_signal_3490, new_AGEMA_signal_3489, new_AGEMA_signal_3488, AddRoundKeyOutput[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2794, new_AGEMA_signal_2793, new_AGEMA_signal_2792, MCOutput[15]}), .c ({new_AGEMA_signal_3298, new_AGEMA_signal_3297, new_AGEMA_signal_3296, AddKeyXOR2_XORInst_3_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_3304, new_AGEMA_signal_3303, new_AGEMA_signal_3302, AddKeyXOR2_XORInst_4_1_n1}), .b ({new_AGEMA_signal_2410, new_AGEMA_signal_2409, new_AGEMA_signal_2408, SelectedKey[17]}), .c ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, new_AGEMA_signal_3494, AddRoundKeyOutput[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2806, new_AGEMA_signal_2805, new_AGEMA_signal_2804, MCOutput[17]}), .c ({new_AGEMA_signal_3304, new_AGEMA_signal_3303, new_AGEMA_signal_3302, AddKeyXOR2_XORInst_4_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, new_AGEMA_signal_3308, AddKeyXOR2_XORInst_4_3_n1}), .b ({new_AGEMA_signal_2428, new_AGEMA_signal_2427, new_AGEMA_signal_2426, SelectedKey[19]}), .c ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, new_AGEMA_signal_3500, AddRoundKeyOutput[19]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2818, new_AGEMA_signal_2817, new_AGEMA_signal_2816, MCOutput[19]}), .c ({new_AGEMA_signal_3310, new_AGEMA_signal_3309, new_AGEMA_signal_3308, AddKeyXOR2_XORInst_4_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, AddKeyXOR2_XORInst_5_1_n1}), .b ({new_AGEMA_signal_2446, new_AGEMA_signal_2445, new_AGEMA_signal_2444, SelectedKey[21]}), .c ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, new_AGEMA_signal_3506, AddRoundKeyOutput[21]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2830, new_AGEMA_signal_2829, new_AGEMA_signal_2828, MCOutput[21]}), .c ({new_AGEMA_signal_3316, new_AGEMA_signal_3315, new_AGEMA_signal_3314, AddKeyXOR2_XORInst_5_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, new_AGEMA_signal_3320, AddKeyXOR2_XORInst_5_3_n1}), .b ({new_AGEMA_signal_1726, new_AGEMA_signal_1725, new_AGEMA_signal_1724, SelectedKey[23]}), .c ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_3512, AddRoundKeyOutput[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2842, new_AGEMA_signal_2841, new_AGEMA_signal_2840, MCOutput[23]}), .c ({new_AGEMA_signal_3322, new_AGEMA_signal_3321, new_AGEMA_signal_3320, AddKeyXOR2_XORInst_5_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_3328, new_AGEMA_signal_3327, new_AGEMA_signal_3326, AddKeyXOR2_XORInst_6_1_n1}), .b ({new_AGEMA_signal_1744, new_AGEMA_signal_1743, new_AGEMA_signal_1742, SelectedKey[25]}), .c ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, AddRoundKeyOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2854, new_AGEMA_signal_2853, new_AGEMA_signal_2852, MCOutput[25]}), .c ({new_AGEMA_signal_3328, new_AGEMA_signal_3327, new_AGEMA_signal_3326, AddKeyXOR2_XORInst_6_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, new_AGEMA_signal_3332, AddKeyXOR2_XORInst_6_3_n1}), .b ({new_AGEMA_signal_1762, new_AGEMA_signal_1761, new_AGEMA_signal_1760, SelectedKey[27]}), .c ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, new_AGEMA_signal_3524, AddRoundKeyOutput[27]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2866, new_AGEMA_signal_2865, new_AGEMA_signal_2864, MCOutput[27]}), .c ({new_AGEMA_signal_3334, new_AGEMA_signal_3333, new_AGEMA_signal_3332, AddKeyXOR2_XORInst_6_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_3340, new_AGEMA_signal_3339, new_AGEMA_signal_3338, AddKeyXOR2_XORInst_7_1_n1}), .b ({new_AGEMA_signal_2464, new_AGEMA_signal_2463, new_AGEMA_signal_2462, SelectedKey[29]}), .c ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, AddRoundKeyOutput[29]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2878, new_AGEMA_signal_2877, new_AGEMA_signal_2876, MCOutput[29]}), .c ({new_AGEMA_signal_3340, new_AGEMA_signal_3339, new_AGEMA_signal_3338, AddKeyXOR2_XORInst_7_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_3346, new_AGEMA_signal_3345, new_AGEMA_signal_3344, AddKeyXOR2_XORInst_7_3_n1}), .b ({new_AGEMA_signal_2482, new_AGEMA_signal_2481, new_AGEMA_signal_2480, SelectedKey[31]}), .c ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, new_AGEMA_signal_3536, AddRoundKeyOutput[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2890, new_AGEMA_signal_2889, new_AGEMA_signal_2888, MCOutput[31]}), .c ({new_AGEMA_signal_3346, new_AGEMA_signal_3345, new_AGEMA_signal_3344, AddKeyXOR2_XORInst_7_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_1_U2 ( .a ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, new_AGEMA_signal_3614, AddKeyXOR2_XORInst_8_1_n1}), .b ({new_AGEMA_signal_1771, new_AGEMA_signal_1770, new_AGEMA_signal_1769, SelectedKey[33]}), .c ({new_AGEMA_signal_3712, new_AGEMA_signal_3711, new_AGEMA_signal_3710, AddRoundKeyOutput[33]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3358, new_AGEMA_signal_3357, new_AGEMA_signal_3356, MCOutput[33]}), .c ({new_AGEMA_signal_3616, new_AGEMA_signal_3615, new_AGEMA_signal_3614, AddKeyXOR2_XORInst_8_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_3_U2 ( .a ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, new_AGEMA_signal_3620, AddKeyXOR2_XORInst_8_3_n1}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, new_AGEMA_signal_2507, SelectedKey[35]}), .c ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, new_AGEMA_signal_3716, AddRoundKeyOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3370, new_AGEMA_signal_3369, new_AGEMA_signal_3368, MCOutput[35]}), .c ({new_AGEMA_signal_3622, new_AGEMA_signal_3621, new_AGEMA_signal_3620, AddKeyXOR2_XORInst_8_3_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_1_U2 ( .a ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, AddKeyXOR2_XORInst_9_1_n1}), .b ({new_AGEMA_signal_2518, new_AGEMA_signal_2517, new_AGEMA_signal_2516, SelectedKey[37]}), .c ({new_AGEMA_signal_3724, new_AGEMA_signal_3723, new_AGEMA_signal_3722, AddRoundKeyOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3382, new_AGEMA_signal_3381, new_AGEMA_signal_3380, MCOutput[37]}), .c ({new_AGEMA_signal_3628, new_AGEMA_signal_3627, new_AGEMA_signal_3626, AddKeyXOR2_XORInst_9_1_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_3_U2 ( .a ({new_AGEMA_signal_3634, new_AGEMA_signal_3633, new_AGEMA_signal_3632, AddKeyXOR2_XORInst_9_3_n1}), .b ({new_AGEMA_signal_1789, new_AGEMA_signal_1788, new_AGEMA_signal_1787, SelectedKey[39]}), .c ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, new_AGEMA_signal_3728, AddRoundKeyOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3394, new_AGEMA_signal_3393, new_AGEMA_signal_3392, MCOutput[39]}), .c ({new_AGEMA_signal_3634, new_AGEMA_signal_3633, new_AGEMA_signal_3632, AddKeyXOR2_XORInst_9_3_n1}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U19 ( .a ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, SubCellInst_SboxInst_0_n15}), .b ({new_AGEMA_signal_1840, new_AGEMA_signal_1839, new_AGEMA_signal_1838, SubCellInst_SboxInst_0_n14}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, new_AGEMA_signal_2075, Feedback[3]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U16 ( .a ({new_AGEMA_signal_1405, new_AGEMA_signal_1404, new_AGEMA_signal_1403, SubCellInst_SboxInst_0_n11}), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, SubCellInst_SboxInst_0_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U12 ( .a ({new_AGEMA_signal_1414, new_AGEMA_signal_1413, new_AGEMA_signal_1412, SubCellInst_SboxInst_0_n6}), .b ({new_AGEMA_signal_1846, new_AGEMA_signal_1845, new_AGEMA_signal_1844, SubCellInst_SboxInst_0_n5}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, new_AGEMA_signal_2081, Feedback[1]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U7 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_1417, new_AGEMA_signal_1416, new_AGEMA_signal_1415, SubCellInst_SboxInst_0_n2}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, SubCellInst_SboxInst_0_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U19 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, new_AGEMA_signal_1424, SubCellInst_SboxInst_1_n15}), .b ({new_AGEMA_signal_1855, new_AGEMA_signal_1854, new_AGEMA_signal_1853, SubCellInst_SboxInst_1_n14}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, new_AGEMA_signal_2087, Feedback[7]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U16 ( .a ({new_AGEMA_signal_1423, new_AGEMA_signal_1422, new_AGEMA_signal_1421, SubCellInst_SboxInst_1_n11}), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_1_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U12 ( .a ({new_AGEMA_signal_1432, new_AGEMA_signal_1431, new_AGEMA_signal_1430, SubCellInst_SboxInst_1_n6}), .b ({new_AGEMA_signal_1861, new_AGEMA_signal_1860, new_AGEMA_signal_1859, SubCellInst_SboxInst_1_n5}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, new_AGEMA_signal_2093, Feedback[5]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U7 ( .a ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_1435, new_AGEMA_signal_1434, new_AGEMA_signal_1433, SubCellInst_SboxInst_1_n2}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, new_AGEMA_signal_1862, SubCellInst_SboxInst_1_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U19 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, SubCellInst_SboxInst_2_n15}), .b ({new_AGEMA_signal_1870, new_AGEMA_signal_1869, new_AGEMA_signal_1868, SubCellInst_SboxInst_2_n14}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, new_AGEMA_signal_2099, Feedback[11]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U16 ( .a ({new_AGEMA_signal_1441, new_AGEMA_signal_1440, new_AGEMA_signal_1439, SubCellInst_SboxInst_2_n11}), .b ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, SubCellInst_SboxInst_2_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U12 ( .a ({new_AGEMA_signal_1450, new_AGEMA_signal_1449, new_AGEMA_signal_1448, SubCellInst_SboxInst_2_n6}), .b ({new_AGEMA_signal_1876, new_AGEMA_signal_1875, new_AGEMA_signal_1874, SubCellInst_SboxInst_2_n5}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, new_AGEMA_signal_2105, Feedback[9]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U7 ( .a ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_1453, new_AGEMA_signal_1452, new_AGEMA_signal_1451, SubCellInst_SboxInst_2_n2}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, new_AGEMA_signal_1877, SubCellInst_SboxInst_2_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U19 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, new_AGEMA_signal_1460, SubCellInst_SboxInst_3_n15}), .b ({new_AGEMA_signal_1885, new_AGEMA_signal_1884, new_AGEMA_signal_1883, SubCellInst_SboxInst_3_n14}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, new_AGEMA_signal_2111, Feedback[15]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U16 ( .a ({new_AGEMA_signal_1459, new_AGEMA_signal_1458, new_AGEMA_signal_1457, SubCellInst_SboxInst_3_n11}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, SubCellInst_SboxInst_3_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U12 ( .a ({new_AGEMA_signal_1468, new_AGEMA_signal_1467, new_AGEMA_signal_1466, SubCellInst_SboxInst_3_n6}), .b ({new_AGEMA_signal_1891, new_AGEMA_signal_1890, new_AGEMA_signal_1889, SubCellInst_SboxInst_3_n5}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, new_AGEMA_signal_2117, Feedback[13]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U7 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_1471, new_AGEMA_signal_1470, new_AGEMA_signal_1469, SubCellInst_SboxInst_3_n2}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_3_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U19 ( .a ({new_AGEMA_signal_1480, new_AGEMA_signal_1479, new_AGEMA_signal_1478, SubCellInst_SboxInst_4_n15}), .b ({new_AGEMA_signal_1900, new_AGEMA_signal_1899, new_AGEMA_signal_1898, SubCellInst_SboxInst_4_n14}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, new_AGEMA_signal_2123, Feedback[19]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U16 ( .a ({new_AGEMA_signal_1477, new_AGEMA_signal_1476, new_AGEMA_signal_1475, SubCellInst_SboxInst_4_n11}), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, new_AGEMA_signal_1901, SubCellInst_SboxInst_4_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U12 ( .a ({new_AGEMA_signal_1486, new_AGEMA_signal_1485, new_AGEMA_signal_1484, SubCellInst_SboxInst_4_n6}), .b ({new_AGEMA_signal_1906, new_AGEMA_signal_1905, new_AGEMA_signal_1904, SubCellInst_SboxInst_4_n5}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_2131, new_AGEMA_signal_2130, new_AGEMA_signal_2129, Feedback[17]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U7 ( .a ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_1489, new_AGEMA_signal_1488, new_AGEMA_signal_1487, SubCellInst_SboxInst_4_n2}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1907, SubCellInst_SboxInst_4_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U19 ( .a ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, new_AGEMA_signal_1496, SubCellInst_SboxInst_5_n15}), .b ({new_AGEMA_signal_1915, new_AGEMA_signal_1914, new_AGEMA_signal_1913, SubCellInst_SboxInst_5_n14}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_2137, new_AGEMA_signal_2136, new_AGEMA_signal_2135, Feedback[23]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U16 ( .a ({new_AGEMA_signal_1495, new_AGEMA_signal_1494, new_AGEMA_signal_1493, SubCellInst_SboxInst_5_n11}), .b ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_5_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U12 ( .a ({new_AGEMA_signal_1504, new_AGEMA_signal_1503, new_AGEMA_signal_1502, SubCellInst_SboxInst_5_n6}), .b ({new_AGEMA_signal_1921, new_AGEMA_signal_1920, new_AGEMA_signal_1919, SubCellInst_SboxInst_5_n5}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, new_AGEMA_signal_2141, Feedback[21]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U7 ( .a ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_1507, new_AGEMA_signal_1506, new_AGEMA_signal_1505, SubCellInst_SboxInst_5_n2}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, SubCellInst_SboxInst_5_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U19 ( .a ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, SubCellInst_SboxInst_6_n15}), .b ({new_AGEMA_signal_1930, new_AGEMA_signal_1929, new_AGEMA_signal_1928, SubCellInst_SboxInst_6_n14}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, new_AGEMA_signal_2147, Feedback[27]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U16 ( .a ({new_AGEMA_signal_1513, new_AGEMA_signal_1512, new_AGEMA_signal_1511, SubCellInst_SboxInst_6_n11}), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, SubCellInst_SboxInst_6_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U12 ( .a ({new_AGEMA_signal_1522, new_AGEMA_signal_1521, new_AGEMA_signal_1520, SubCellInst_SboxInst_6_n6}), .b ({new_AGEMA_signal_1936, new_AGEMA_signal_1935, new_AGEMA_signal_1934, SubCellInst_SboxInst_6_n5}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, new_AGEMA_signal_2153, Feedback[25]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U7 ( .a ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_1525, new_AGEMA_signal_1524, new_AGEMA_signal_1523, SubCellInst_SboxInst_6_n2}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1937, SubCellInst_SboxInst_6_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U19 ( .a ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, SubCellInst_SboxInst_7_n15}), .b ({new_AGEMA_signal_1945, new_AGEMA_signal_1944, new_AGEMA_signal_1943, SubCellInst_SboxInst_7_n14}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, new_AGEMA_signal_2159, Feedback[31]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U16 ( .a ({new_AGEMA_signal_1531, new_AGEMA_signal_1530, new_AGEMA_signal_1529, SubCellInst_SboxInst_7_n11}), .b ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_7_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U12 ( .a ({new_AGEMA_signal_1540, new_AGEMA_signal_1539, new_AGEMA_signal_1538, SubCellInst_SboxInst_7_n6}), .b ({new_AGEMA_signal_1951, new_AGEMA_signal_1950, new_AGEMA_signal_1949, SubCellInst_SboxInst_7_n5}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, new_AGEMA_signal_2165, Feedback[29]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U7 ( .a ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_1543, new_AGEMA_signal_1542, new_AGEMA_signal_1541, SubCellInst_SboxInst_7_n2}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_7_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U19 ( .a ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, SubCellInst_SboxInst_8_n15}), .b ({new_AGEMA_signal_1960, new_AGEMA_signal_1959, new_AGEMA_signal_1958, SubCellInst_SboxInst_8_n14}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, new_AGEMA_signal_2171, Feedback[35]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U16 ( .a ({new_AGEMA_signal_1549, new_AGEMA_signal_1548, new_AGEMA_signal_1547, SubCellInst_SboxInst_8_n11}), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, SubCellInst_SboxInst_8_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U12 ( .a ({new_AGEMA_signal_1558, new_AGEMA_signal_1557, new_AGEMA_signal_1556, SubCellInst_SboxInst_8_n6}), .b ({new_AGEMA_signal_1966, new_AGEMA_signal_1965, new_AGEMA_signal_1964, SubCellInst_SboxInst_8_n5}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, new_AGEMA_signal_2177, Feedback[33]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U7 ( .a ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_1561, new_AGEMA_signal_1560, new_AGEMA_signal_1559, SubCellInst_SboxInst_8_n2}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, SubCellInst_SboxInst_8_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U19 ( .a ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, SubCellInst_SboxInst_9_n15}), .b ({new_AGEMA_signal_1975, new_AGEMA_signal_1974, new_AGEMA_signal_1973, SubCellInst_SboxInst_9_n14}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, new_AGEMA_signal_2183, Feedback[39]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U16 ( .a ({new_AGEMA_signal_1567, new_AGEMA_signal_1566, new_AGEMA_signal_1565, SubCellInst_SboxInst_9_n11}), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_9_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U12 ( .a ({new_AGEMA_signal_1576, new_AGEMA_signal_1575, new_AGEMA_signal_1574, SubCellInst_SboxInst_9_n6}), .b ({new_AGEMA_signal_1981, new_AGEMA_signal_1980, new_AGEMA_signal_1979, SubCellInst_SboxInst_9_n5}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, new_AGEMA_signal_2189, Feedback[37]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U7 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_1579, new_AGEMA_signal_1578, new_AGEMA_signal_1577, SubCellInst_SboxInst_9_n2}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_9_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U19 ( .a ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, SubCellInst_SboxInst_10_n15}), .b ({new_AGEMA_signal_1990, new_AGEMA_signal_1989, new_AGEMA_signal_1988, SubCellInst_SboxInst_10_n14}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, new_AGEMA_signal_2195, Feedback[43]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U16 ( .a ({new_AGEMA_signal_1585, new_AGEMA_signal_1584, new_AGEMA_signal_1583, SubCellInst_SboxInst_10_n11}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, SubCellInst_SboxInst_10_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U12 ( .a ({new_AGEMA_signal_1594, new_AGEMA_signal_1593, new_AGEMA_signal_1592, SubCellInst_SboxInst_10_n6}), .b ({new_AGEMA_signal_1996, new_AGEMA_signal_1995, new_AGEMA_signal_1994, SubCellInst_SboxInst_10_n5}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, new_AGEMA_signal_2201, Feedback[41]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U7 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_1597, new_AGEMA_signal_1596, new_AGEMA_signal_1595, SubCellInst_SboxInst_10_n2}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, SubCellInst_SboxInst_10_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U19 ( .a ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, SubCellInst_SboxInst_11_n15}), .b ({new_AGEMA_signal_2005, new_AGEMA_signal_2004, new_AGEMA_signal_2003, SubCellInst_SboxInst_11_n14}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, new_AGEMA_signal_2207, Feedback[47]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U16 ( .a ({new_AGEMA_signal_1603, new_AGEMA_signal_1602, new_AGEMA_signal_1601, SubCellInst_SboxInst_11_n11}), .b ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_11_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U12 ( .a ({new_AGEMA_signal_1612, new_AGEMA_signal_1611, new_AGEMA_signal_1610, SubCellInst_SboxInst_11_n6}), .b ({new_AGEMA_signal_2011, new_AGEMA_signal_2010, new_AGEMA_signal_2009, SubCellInst_SboxInst_11_n5}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, new_AGEMA_signal_2213, Feedback[45]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U7 ( .a ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_1615, new_AGEMA_signal_1614, new_AGEMA_signal_1613, SubCellInst_SboxInst_11_n2}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_11_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U19 ( .a ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, SubCellInst_SboxInst_12_n15}), .b ({new_AGEMA_signal_2020, new_AGEMA_signal_2019, new_AGEMA_signal_2018, SubCellInst_SboxInst_12_n14}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, new_AGEMA_signal_2219, Feedback[51]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U16 ( .a ({new_AGEMA_signal_1621, new_AGEMA_signal_1620, new_AGEMA_signal_1619, SubCellInst_SboxInst_12_n11}), .b ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, SubCellInst_SboxInst_12_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U12 ( .a ({new_AGEMA_signal_1630, new_AGEMA_signal_1629, new_AGEMA_signal_1628, SubCellInst_SboxInst_12_n6}), .b ({new_AGEMA_signal_2026, new_AGEMA_signal_2025, new_AGEMA_signal_2024, SubCellInst_SboxInst_12_n5}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, new_AGEMA_signal_2225, Feedback[49]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U7 ( .a ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_1633, new_AGEMA_signal_1632, new_AGEMA_signal_1631, SubCellInst_SboxInst_12_n2}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, SubCellInst_SboxInst_12_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U19 ( .a ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, SubCellInst_SboxInst_13_n15}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, new_AGEMA_signal_2033, SubCellInst_SboxInst_13_n14}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, new_AGEMA_signal_2231, Feedback[55]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U16 ( .a ({new_AGEMA_signal_1639, new_AGEMA_signal_1638, new_AGEMA_signal_1637, SubCellInst_SboxInst_13_n11}), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, new_AGEMA_signal_2036, SubCellInst_SboxInst_13_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U12 ( .a ({new_AGEMA_signal_1648, new_AGEMA_signal_1647, new_AGEMA_signal_1646, SubCellInst_SboxInst_13_n6}), .b ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, new_AGEMA_signal_2039, SubCellInst_SboxInst_13_n5}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, new_AGEMA_signal_2237, Feedback[53]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U7 ( .a ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_1651, new_AGEMA_signal_1650, new_AGEMA_signal_1649, SubCellInst_SboxInst_13_n2}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, SubCellInst_SboxInst_13_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U19 ( .a ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, SubCellInst_SboxInst_14_n15}), .b ({new_AGEMA_signal_2050, new_AGEMA_signal_2049, new_AGEMA_signal_2048, SubCellInst_SboxInst_14_n14}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, new_AGEMA_signal_2243, Feedback[59]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U16 ( .a ({new_AGEMA_signal_1657, new_AGEMA_signal_1656, new_AGEMA_signal_1655, SubCellInst_SboxInst_14_n11}), .b ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, SubCellInst_SboxInst_14_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U12 ( .a ({new_AGEMA_signal_1666, new_AGEMA_signal_1665, new_AGEMA_signal_1664, SubCellInst_SboxInst_14_n6}), .b ({new_AGEMA_signal_2056, new_AGEMA_signal_2055, new_AGEMA_signal_2054, SubCellInst_SboxInst_14_n5}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, new_AGEMA_signal_2249, Feedback[57]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U7 ( .a ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_1669, new_AGEMA_signal_1668, new_AGEMA_signal_1667, SubCellInst_SboxInst_14_n2}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, SubCellInst_SboxInst_14_n3}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U19 ( .a ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1676, SubCellInst_SboxInst_15_n15}), .b ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, new_AGEMA_signal_2063, SubCellInst_SboxInst_15_n14}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, new_AGEMA_signal_2255, Feedback[63]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U16 ( .a ({new_AGEMA_signal_1675, new_AGEMA_signal_1674, new_AGEMA_signal_1673, SubCellInst_SboxInst_15_n11}), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, SubCellInst_SboxInst_15_n12}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U12 ( .a ({new_AGEMA_signal_1684, new_AGEMA_signal_1683, new_AGEMA_signal_1682, SubCellInst_SboxInst_15_n6}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, new_AGEMA_signal_2069, SubCellInst_SboxInst_15_n5}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, new_AGEMA_signal_2261, Feedback[61]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U7 ( .a ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_1687, new_AGEMA_signal_1686, new_AGEMA_signal_1685, SubCellInst_SboxInst_15_n2}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, SubCellInst_SboxInst_15_n3}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, Feedback[0]}), .a ({plaintext_s3[0], plaintext_s2[0], plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, MCOutput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, Feedback[2]}), .a ({plaintext_s3[2], plaintext_s2[2], plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, MCOutput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, Feedback[4]}), .a ({plaintext_s3[4], plaintext_s2[4], plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, MCOutput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, Feedback[6]}), .a ({plaintext_s3[6], plaintext_s2[6], plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, MCOutput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, Feedback[8]}), .a ({plaintext_s3[8], plaintext_s2[8], plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, new_AGEMA_signal_2750, MCOutput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, Feedback[10]}), .a ({plaintext_s3[10], plaintext_s2[10], plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, new_AGEMA_signal_2120, Feedback[12]}), .a ({plaintext_s3[12], plaintext_s2[12], plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCOutput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, Feedback[14]}), .a ({plaintext_s3[14], plaintext_s2[14], plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, Feedback[16]}), .a ({plaintext_s3[16], plaintext_s2[16], plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, MCOutput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, Feedback[18]}), .a ({plaintext_s3[18], plaintext_s2[18], plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, MCOutput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, Feedback[20]}), .a ({plaintext_s3[20], plaintext_s2[20], plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, MCOutput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, Feedback[22]}), .a ({plaintext_s3[22], plaintext_s2[22], plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, MCOutput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, new_AGEMA_signal_2156, Feedback[24]}), .a ({plaintext_s3[24], plaintext_s2[24], plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, MCOutput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, new_AGEMA_signal_2150, Feedback[26]}), .a ({plaintext_s3[26], plaintext_s2[26], plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, Feedback[28]}), .a ({plaintext_s3[28], plaintext_s2[28], plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, Feedback[30]}), .a ({plaintext_s3[30], plaintext_s2[30], plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, new_AGEMA_signal_2180, Feedback[32]}), .a ({plaintext_s3[32], plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, MCInput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, Feedback[34]}), .a ({plaintext_s3[34], plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, MCInput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, Feedback[36]}), .a ({plaintext_s3[36], plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, MCInput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, Feedback[38]}), .a ({plaintext_s3[38], plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, MCInput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, Feedback[40]}), .a ({plaintext_s3[40], plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, new_AGEMA_signal_2942, MCInput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, Feedback[42]}), .a ({plaintext_s3[42], plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, MCInput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, new_AGEMA_signal_2216, Feedback[44]}), .a ({plaintext_s3[44], plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, new_AGEMA_signal_2966, MCInput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, Feedback[46]}), .a ({plaintext_s3[46], plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_2980, new_AGEMA_signal_2979, new_AGEMA_signal_2978, MCInput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, Feedback[48]}), .a ({plaintext_s3[48], plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, MCInput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, Feedback[50]}), .a ({plaintext_s3[50], plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_3004, new_AGEMA_signal_3003, new_AGEMA_signal_3002, MCInput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, new_AGEMA_signal_2240, Feedback[52]}), .a ({plaintext_s3[52], plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, MCInput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, Feedback[54]}), .a ({plaintext_s3[54], plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, MCInput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, Feedback[56]}), .a ({plaintext_s3[56], plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_3040, new_AGEMA_signal_3039, new_AGEMA_signal_3038, MCInput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, Feedback[58]}), .a ({plaintext_s3[58], plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, MCInput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, Feedback[60]}), .a ({plaintext_s3[60], plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, MCInput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) InputMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, Feedback[62]}), .a ({plaintext_s3[62], plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, MCInput[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_0_U3 ( .a ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, MCInst_XOR_r0_Inst_0_n2}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, MCInst_XOR_r0_Inst_0_n1}), .c ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, new_AGEMA_signal_3347, MCOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_0_U2 ( .a ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, MCOutput[16]}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, MCOutput[0]}), .c ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, new_AGEMA_signal_3107, MCInst_XOR_r0_Inst_0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2992, new_AGEMA_signal_2991, new_AGEMA_signal_2990, MCInput[48]}), .c ({new_AGEMA_signal_3112, new_AGEMA_signal_3111, new_AGEMA_signal_3110, MCInst_XOR_r0_Inst_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_0_U2 ( .a ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, new_AGEMA_signal_3113, MCInst_XOR_r1_Inst_0_n1}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, MCOutput[0]}), .c ({new_AGEMA_signal_3352, new_AGEMA_signal_3351, new_AGEMA_signal_3350, MCOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2896, new_AGEMA_signal_2895, new_AGEMA_signal_2894, MCInput[32]}), .c ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, new_AGEMA_signal_3113, MCInst_XOR_r1_Inst_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_2_U3 ( .a ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, new_AGEMA_signal_3128, MCInst_XOR_r0_Inst_2_n2}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, new_AGEMA_signal_3125, MCInst_XOR_r0_Inst_2_n1}), .c ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, new_AGEMA_signal_3359, MCOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_2_U2 ( .a ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, MCOutput[18]}), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, MCOutput[2]}), .c ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, new_AGEMA_signal_3125, MCInst_XOR_r0_Inst_2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3004, new_AGEMA_signal_3003, new_AGEMA_signal_3002, MCInput[50]}), .c ({new_AGEMA_signal_3130, new_AGEMA_signal_3129, new_AGEMA_signal_3128, MCInst_XOR_r0_Inst_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_2_U2 ( .a ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, new_AGEMA_signal_3131, MCInst_XOR_r1_Inst_2_n1}), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, MCOutput[2]}), .c ({new_AGEMA_signal_3364, new_AGEMA_signal_3363, new_AGEMA_signal_3362, MCOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2908, new_AGEMA_signal_2907, new_AGEMA_signal_2906, MCInput[34]}), .c ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, new_AGEMA_signal_3131, MCInst_XOR_r1_Inst_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_4_U3 ( .a ({new_AGEMA_signal_3148, new_AGEMA_signal_3147, new_AGEMA_signal_3146, MCInst_XOR_r0_Inst_4_n2}), .b ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, MCInst_XOR_r0_Inst_4_n1}), .c ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, new_AGEMA_signal_3371, MCOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_4_U2 ( .a ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, MCOutput[20]}), .b ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, MCOutput[4]}), .c ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, new_AGEMA_signal_3143, MCInst_XOR_r0_Inst_4_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_4_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3016, new_AGEMA_signal_3015, new_AGEMA_signal_3014, MCInput[52]}), .c ({new_AGEMA_signal_3148, new_AGEMA_signal_3147, new_AGEMA_signal_3146, MCInst_XOR_r0_Inst_4_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_4_U2 ( .a ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, new_AGEMA_signal_3149, MCInst_XOR_r1_Inst_4_n1}), .b ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, MCOutput[4]}), .c ({new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, MCOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_4_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2920, new_AGEMA_signal_2919, new_AGEMA_signal_2918, MCInput[36]}), .c ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, new_AGEMA_signal_3149, MCInst_XOR_r1_Inst_4_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_6_U3 ( .a ({new_AGEMA_signal_3166, new_AGEMA_signal_3165, new_AGEMA_signal_3164, MCInst_XOR_r0_Inst_6_n2}), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, new_AGEMA_signal_3161, MCInst_XOR_r0_Inst_6_n1}), .c ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, MCOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_6_U2 ( .a ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, MCOutput[22]}), .b ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, MCOutput[6]}), .c ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, new_AGEMA_signal_3161, MCInst_XOR_r0_Inst_6_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_6_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3028, new_AGEMA_signal_3027, new_AGEMA_signal_3026, MCInput[54]}), .c ({new_AGEMA_signal_3166, new_AGEMA_signal_3165, new_AGEMA_signal_3164, MCInst_XOR_r0_Inst_6_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_6_U2 ( .a ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, new_AGEMA_signal_3167, MCInst_XOR_r1_Inst_6_n1}), .b ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, MCOutput[6]}), .c ({new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, MCOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_6_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2932, new_AGEMA_signal_2931, new_AGEMA_signal_2930, MCInput[38]}), .c ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, new_AGEMA_signal_3167, MCInst_XOR_r1_Inst_6_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_8_U3 ( .a ({new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, MCInst_XOR_r0_Inst_8_n2}), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, new_AGEMA_signal_3179, MCInst_XOR_r0_Inst_8_n1}), .c ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, MCOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_8_U2 ( .a ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, MCOutput[24]}), .b ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, new_AGEMA_signal_2750, MCOutput[8]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, new_AGEMA_signal_3179, MCInst_XOR_r0_Inst_8_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_8_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3040, new_AGEMA_signal_3039, new_AGEMA_signal_3038, MCInput[56]}), .c ({new_AGEMA_signal_3184, new_AGEMA_signal_3183, new_AGEMA_signal_3182, MCInst_XOR_r0_Inst_8_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_8_U2 ( .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, new_AGEMA_signal_3185, MCInst_XOR_r1_Inst_8_n1}), .b ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, new_AGEMA_signal_2750, MCOutput[8]}), .c ({new_AGEMA_signal_3400, new_AGEMA_signal_3399, new_AGEMA_signal_3398, MCOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_8_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2944, new_AGEMA_signal_2943, new_AGEMA_signal_2942, MCInput[40]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, new_AGEMA_signal_3185, MCInst_XOR_r1_Inst_8_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_10_U3 ( .a ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, new_AGEMA_signal_3200, MCInst_XOR_r0_Inst_10_n2}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, new_AGEMA_signal_3197, MCInst_XOR_r0_Inst_10_n1}), .c ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, new_AGEMA_signal_3407, MCOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_10_U2 ( .a ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[26]}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[10]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, new_AGEMA_signal_3197, MCInst_XOR_r0_Inst_10_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_10_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3052, new_AGEMA_signal_3051, new_AGEMA_signal_3050, MCInput[58]}), .c ({new_AGEMA_signal_3202, new_AGEMA_signal_3201, new_AGEMA_signal_3200, MCInst_XOR_r0_Inst_10_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_10_U2 ( .a ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, new_AGEMA_signal_3203, MCInst_XOR_r1_Inst_10_n1}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[10]}), .c ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, MCOutput[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_10_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2956, new_AGEMA_signal_2955, new_AGEMA_signal_2954, MCInput[42]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, new_AGEMA_signal_3203, MCInst_XOR_r1_Inst_10_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_12_U3 ( .a ({new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_3218, MCInst_XOR_r0_Inst_12_n2}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, new_AGEMA_signal_3215, MCInst_XOR_r0_Inst_12_n1}), .c ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, MCOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_12_U2 ( .a ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[28]}), .b ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCOutput[12]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, new_AGEMA_signal_3215, MCInst_XOR_r0_Inst_12_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_12_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3064, new_AGEMA_signal_3063, new_AGEMA_signal_3062, MCInput[60]}), .c ({new_AGEMA_signal_3220, new_AGEMA_signal_3219, new_AGEMA_signal_3218, MCInst_XOR_r0_Inst_12_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_12_U2 ( .a ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, new_AGEMA_signal_3221, MCInst_XOR_r1_Inst_12_n1}), .b ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCOutput[12]}), .c ({new_AGEMA_signal_3424, new_AGEMA_signal_3423, new_AGEMA_signal_3422, MCOutput[44]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_12_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2968, new_AGEMA_signal_2967, new_AGEMA_signal_2966, MCInput[44]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, new_AGEMA_signal_3221, MCInst_XOR_r1_Inst_12_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_14_U3 ( .a ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, new_AGEMA_signal_3236, MCInst_XOR_r0_Inst_14_n2}), .b ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, new_AGEMA_signal_3233, MCInst_XOR_r0_Inst_14_n1}), .c ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, MCOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_14_U2 ( .a ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[30]}), .b ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[14]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, new_AGEMA_signal_3233, MCInst_XOR_r0_Inst_14_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r0_Inst_14_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3076, new_AGEMA_signal_3075, new_AGEMA_signal_3074, MCInput[62]}), .c ({new_AGEMA_signal_3238, new_AGEMA_signal_3237, new_AGEMA_signal_3236, MCInst_XOR_r0_Inst_14_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_14_U2 ( .a ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, new_AGEMA_signal_3239, MCInst_XOR_r1_Inst_14_n1}), .b ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[14]}), .c ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, new_AGEMA_signal_3434, MCOutput[46]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MCInst_XOR_r1_Inst_14_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2980, new_AGEMA_signal_2979, new_AGEMA_signal_2978, MCInput[46]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, new_AGEMA_signal_3239, MCInst_XOR_r1_Inst_14_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, AddKeyXOR1_XORInst_0_0_n1}), .b ({new_AGEMA_signal_2608, new_AGEMA_signal_2607, new_AGEMA_signal_2606, SelectedKey[48]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, AddRoundKeyOutput[48]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, new_AGEMA_signal_3347, MCOutput[48]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, new_AGEMA_signal_3539, AddKeyXOR1_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, AddKeyXOR1_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2626, new_AGEMA_signal_2625, new_AGEMA_signal_2624, SelectedKey[50]}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, new_AGEMA_signal_3641, AddRoundKeyOutput[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, new_AGEMA_signal_3359, MCOutput[50]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, new_AGEMA_signal_3545, AddKeyXOR1_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, new_AGEMA_signal_3551, AddKeyXOR1_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2644, new_AGEMA_signal_2643, new_AGEMA_signal_2642, SelectedKey[52]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, new_AGEMA_signal_3647, AddRoundKeyOutput[52]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, new_AGEMA_signal_3371, MCOutput[52]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, new_AGEMA_signal_3551, AddKeyXOR1_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, new_AGEMA_signal_3557, AddKeyXOR1_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1807, new_AGEMA_signal_1806, new_AGEMA_signal_1805, SelectedKey[54]}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, new_AGEMA_signal_3653, AddRoundKeyOutput[54]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, new_AGEMA_signal_3383, MCOutput[54]}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, new_AGEMA_signal_3557, AddKeyXOR1_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, AddKeyXOR1_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1816, new_AGEMA_signal_1815, new_AGEMA_signal_1814, SelectedKey[56]}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, new_AGEMA_signal_3659, AddRoundKeyOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, new_AGEMA_signal_3395, MCOutput[56]}), .c ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, new_AGEMA_signal_3563, AddKeyXOR1_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, new_AGEMA_signal_3569, AddKeyXOR1_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, new_AGEMA_signal_2669, SelectedKey[58]}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, new_AGEMA_signal_3665, AddRoundKeyOutput[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, new_AGEMA_signal_3407, MCOutput[58]}), .c ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, new_AGEMA_signal_3569, AddKeyXOR1_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3575, AddKeyXOR1_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2680, new_AGEMA_signal_2679, new_AGEMA_signal_2678, SelectedKey[60]}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, AddRoundKeyOutput[60]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, new_AGEMA_signal_3419, MCOutput[60]}), .c ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, new_AGEMA_signal_3575, AddKeyXOR1_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, new_AGEMA_signal_3581, AddKeyXOR1_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1834, new_AGEMA_signal_1833, new_AGEMA_signal_1832, SelectedKey[62]}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, new_AGEMA_signal_3677, AddRoundKeyOutput[62]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR1_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, new_AGEMA_signal_3431, MCOutput[62]}), .c ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, new_AGEMA_signal_3581, AddKeyXOR1_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, new_AGEMA_signal_3587, AddKeyConstXOR_XORInst_0_0_n2}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, new_AGEMA_signal_3083, AddKeyConstXOR_XORInst_0_0_n1}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, new_AGEMA_signal_3683, AddRoundKeyOutput[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3400, new_AGEMA_signal_3399, new_AGEMA_signal_3398, MCOutput[40]}), .c ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, new_AGEMA_signal_3587, AddKeyConstXOR_XORInst_0_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, new_AGEMA_signal_3593, AddKeyConstXOR_XORInst_0_2_n2}), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, new_AGEMA_signal_3089, AddKeyConstXOR_XORInst_0_2_n1}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, new_AGEMA_signal_3689, AddRoundKeyOutput[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3412, new_AGEMA_signal_3411, new_AGEMA_signal_3410, MCOutput[42]}), .c ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, new_AGEMA_signal_3593, AddKeyConstXOR_XORInst_0_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, AddKeyConstXOR_XORInst_1_0_n2}), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, new_AGEMA_signal_3095, AddKeyConstXOR_XORInst_1_0_n1}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, new_AGEMA_signal_3695, AddRoundKeyOutput[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3424, new_AGEMA_signal_3423, new_AGEMA_signal_3422, MCOutput[44]}), .c ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, new_AGEMA_signal_3599, AddKeyConstXOR_XORInst_1_0_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, new_AGEMA_signal_3605, AddKeyConstXOR_XORInst_1_2_n2}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, new_AGEMA_signal_3101, AddKeyConstXOR_XORInst_1_2_n1}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, new_AGEMA_signal_3701, AddRoundKeyOutput[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3436, new_AGEMA_signal_3435, new_AGEMA_signal_3434, MCOutput[46]}), .c ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, new_AGEMA_signal_3605, AddKeyConstXOR_XORInst_1_2_n2}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, AddKeyXOR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1699, new_AGEMA_signal_1698, new_AGEMA_signal_1697, SelectedKey[0]}), .c ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, AddRoundKeyOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2704, new_AGEMA_signal_2703, new_AGEMA_signal_2702, MCOutput[0]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, new_AGEMA_signal_3251, AddKeyXOR2_XORInst_0_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, new_AGEMA_signal_3257, AddKeyXOR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1708, new_AGEMA_signal_1707, new_AGEMA_signal_1706, SelectedKey[2]}), .c ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, AddRoundKeyOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2716, new_AGEMA_signal_2715, new_AGEMA_signal_2714, MCOutput[2]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, new_AGEMA_signal_3257, AddKeyXOR2_XORInst_0_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, new_AGEMA_signal_3263, AddKeyXOR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, new_AGEMA_signal_2291, SelectedKey[4]}), .c ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, AddRoundKeyOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2728, new_AGEMA_signal_2727, new_AGEMA_signal_2726, MCOutput[4]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, new_AGEMA_signal_3263, AddKeyXOR2_XORInst_1_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, new_AGEMA_signal_3269, AddKeyXOR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, new_AGEMA_signal_2309, SelectedKey[6]}), .c ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, new_AGEMA_signal_3461, AddRoundKeyOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2740, new_AGEMA_signal_2739, new_AGEMA_signal_2738, MCOutput[6]}), .c ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, new_AGEMA_signal_3269, AddKeyXOR2_XORInst_1_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, new_AGEMA_signal_3275, AddKeyXOR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, new_AGEMA_signal_2327, SelectedKey[8]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, AddRoundKeyOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2752, new_AGEMA_signal_2751, new_AGEMA_signal_2750, MCOutput[8]}), .c ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, new_AGEMA_signal_3275, AddKeyXOR2_XORInst_2_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, new_AGEMA_signal_3281, AddKeyXOR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2347, new_AGEMA_signal_2346, new_AGEMA_signal_2345, SelectedKey[10]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, AddRoundKeyOutput[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2764, new_AGEMA_signal_2763, new_AGEMA_signal_2762, MCOutput[10]}), .c ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, new_AGEMA_signal_3281, AddKeyXOR2_XORInst_2_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, AddKeyXOR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_2365, new_AGEMA_signal_2364, new_AGEMA_signal_2363, SelectedKey[12]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, new_AGEMA_signal_3479, AddRoundKeyOutput[12]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2776, new_AGEMA_signal_2775, new_AGEMA_signal_2774, MCOutput[12]}), .c ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, new_AGEMA_signal_3287, AddKeyXOR2_XORInst_3_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, new_AGEMA_signal_3293, AddKeyXOR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2383, new_AGEMA_signal_2382, new_AGEMA_signal_2381, SelectedKey[14]}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, new_AGEMA_signal_3485, AddRoundKeyOutput[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2788, new_AGEMA_signal_2787, new_AGEMA_signal_2786, MCOutput[14]}), .c ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, new_AGEMA_signal_3293, AddKeyXOR2_XORInst_3_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, new_AGEMA_signal_3299, AddKeyXOR2_XORInst_4_0_n1}), .b ({new_AGEMA_signal_2401, new_AGEMA_signal_2400, new_AGEMA_signal_2399, SelectedKey[16]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, AddRoundKeyOutput[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2800, new_AGEMA_signal_2799, new_AGEMA_signal_2798, MCOutput[16]}), .c ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, new_AGEMA_signal_3299, AddKeyXOR2_XORInst_4_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, new_AGEMA_signal_3305, AddKeyXOR2_XORInst_4_2_n1}), .b ({new_AGEMA_signal_2419, new_AGEMA_signal_2418, new_AGEMA_signal_2417, SelectedKey[18]}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, new_AGEMA_signal_3497, AddRoundKeyOutput[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2812, new_AGEMA_signal_2811, new_AGEMA_signal_2810, MCOutput[18]}), .c ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, new_AGEMA_signal_3305, AddKeyXOR2_XORInst_4_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, new_AGEMA_signal_3311, AddKeyXOR2_XORInst_5_0_n1}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, new_AGEMA_signal_2435, SelectedKey[20]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, AddRoundKeyOutput[20]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2824, new_AGEMA_signal_2823, new_AGEMA_signal_2822, MCOutput[20]}), .c ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, new_AGEMA_signal_3311, AddKeyXOR2_XORInst_5_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, new_AGEMA_signal_3317, AddKeyXOR2_XORInst_5_2_n1}), .b ({new_AGEMA_signal_1717, new_AGEMA_signal_1716, new_AGEMA_signal_1715, SelectedKey[22]}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_3509, AddRoundKeyOutput[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2836, new_AGEMA_signal_2835, new_AGEMA_signal_2834, MCOutput[22]}), .c ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, new_AGEMA_signal_3317, AddKeyXOR2_XORInst_5_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, AddKeyXOR2_XORInst_6_0_n1}), .b ({new_AGEMA_signal_1735, new_AGEMA_signal_1734, new_AGEMA_signal_1733, SelectedKey[24]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, new_AGEMA_signal_3515, AddRoundKeyOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2848, new_AGEMA_signal_2847, new_AGEMA_signal_2846, MCOutput[24]}), .c ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, new_AGEMA_signal_3323, AddKeyXOR2_XORInst_6_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, new_AGEMA_signal_3329, AddKeyXOR2_XORInst_6_2_n1}), .b ({new_AGEMA_signal_1753, new_AGEMA_signal_1752, new_AGEMA_signal_1751, SelectedKey[26]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, new_AGEMA_signal_3521, AddRoundKeyOutput[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2860, new_AGEMA_signal_2859, new_AGEMA_signal_2858, MCOutput[26]}), .c ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, new_AGEMA_signal_3329, AddKeyXOR2_XORInst_6_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, new_AGEMA_signal_3335, AddKeyXOR2_XORInst_7_0_n1}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, new_AGEMA_signal_2453, SelectedKey[28]}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, AddRoundKeyOutput[28]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2872, new_AGEMA_signal_2871, new_AGEMA_signal_2870, MCOutput[28]}), .c ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, new_AGEMA_signal_3335, AddKeyXOR2_XORInst_7_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, new_AGEMA_signal_3341, AddKeyXOR2_XORInst_7_2_n1}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, new_AGEMA_signal_2471, SelectedKey[30]}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, new_AGEMA_signal_3533, AddRoundKeyOutput[30]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2884, new_AGEMA_signal_2883, new_AGEMA_signal_2882, MCOutput[30]}), .c ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, new_AGEMA_signal_3341, AddKeyXOR2_XORInst_7_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_0_U2 ( .a ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, AddKeyXOR2_XORInst_8_0_n1}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, new_AGEMA_signal_2489, SelectedKey[32]}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, AddRoundKeyOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3352, new_AGEMA_signal_3351, new_AGEMA_signal_3350, MCOutput[32]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, new_AGEMA_signal_3611, AddKeyXOR2_XORInst_8_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_2_U2 ( .a ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3617, AddKeyXOR2_XORInst_8_2_n1}), .b ({new_AGEMA_signal_2500, new_AGEMA_signal_2499, new_AGEMA_signal_2498, SelectedKey[34]}), .c ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, new_AGEMA_signal_3713, AddRoundKeyOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_8_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3364, new_AGEMA_signal_3363, new_AGEMA_signal_3362, MCOutput[34]}), .c ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, new_AGEMA_signal_3617, AddKeyXOR2_XORInst_8_2_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_0_U2 ( .a ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, new_AGEMA_signal_3623, AddKeyXOR2_XORInst_9_0_n1}), .b ({new_AGEMA_signal_1780, new_AGEMA_signal_1779, new_AGEMA_signal_1778, SelectedKey[36]}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, new_AGEMA_signal_3719, AddRoundKeyOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3376, new_AGEMA_signal_3375, new_AGEMA_signal_3374, MCOutput[36]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, new_AGEMA_signal_3623, AddKeyXOR2_XORInst_9_0_n1}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_2_U2 ( .a ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, new_AGEMA_signal_3629, AddKeyXOR2_XORInst_9_2_n1}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, new_AGEMA_signal_2525, SelectedKey[38]}), .c ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, AddRoundKeyOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) AddKeyXOR2_XORInst_9_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3388, new_AGEMA_signal_3387, new_AGEMA_signal_3386, MCOutput[38]}), .c ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, new_AGEMA_signal_3629, AddKeyXOR2_XORInst_9_2_n1}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U17 ( .a ({new_AGEMA_signal_1408, new_AGEMA_signal_1407, new_AGEMA_signal_1406, SubCellInst_SboxInst_0_n15}), .b ({new_AGEMA_signal_1843, new_AGEMA_signal_1842, new_AGEMA_signal_1841, SubCellInst_SboxInst_0_n12}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_2080, new_AGEMA_signal_2079, new_AGEMA_signal_2078, Feedback[2]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U8 ( .a ({new_AGEMA_signal_1420, new_AGEMA_signal_1419, new_AGEMA_signal_1418, SubCellInst_SboxInst_0_n13}), .b ({new_AGEMA_signal_1849, new_AGEMA_signal_1848, new_AGEMA_signal_1847, SubCellInst_SboxInst_0_n3}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_2086, new_AGEMA_signal_2085, new_AGEMA_signal_2084, Feedback[0]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U17 ( .a ({new_AGEMA_signal_1426, new_AGEMA_signal_1425, new_AGEMA_signal_1424, SubCellInst_SboxInst_1_n15}), .b ({new_AGEMA_signal_1858, new_AGEMA_signal_1857, new_AGEMA_signal_1856, SubCellInst_SboxInst_1_n12}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_2092, new_AGEMA_signal_2091, new_AGEMA_signal_2090, Feedback[6]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U8 ( .a ({new_AGEMA_signal_1438, new_AGEMA_signal_1437, new_AGEMA_signal_1436, SubCellInst_SboxInst_1_n13}), .b ({new_AGEMA_signal_1864, new_AGEMA_signal_1863, new_AGEMA_signal_1862, SubCellInst_SboxInst_1_n3}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_2098, new_AGEMA_signal_2097, new_AGEMA_signal_2096, Feedback[4]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U17 ( .a ({new_AGEMA_signal_1444, new_AGEMA_signal_1443, new_AGEMA_signal_1442, SubCellInst_SboxInst_2_n15}), .b ({new_AGEMA_signal_1873, new_AGEMA_signal_1872, new_AGEMA_signal_1871, SubCellInst_SboxInst_2_n12}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_2104, new_AGEMA_signal_2103, new_AGEMA_signal_2102, Feedback[10]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U8 ( .a ({new_AGEMA_signal_1456, new_AGEMA_signal_1455, new_AGEMA_signal_1454, SubCellInst_SboxInst_2_n13}), .b ({new_AGEMA_signal_1879, new_AGEMA_signal_1878, new_AGEMA_signal_1877, SubCellInst_SboxInst_2_n3}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_2110, new_AGEMA_signal_2109, new_AGEMA_signal_2108, Feedback[8]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U17 ( .a ({new_AGEMA_signal_1462, new_AGEMA_signal_1461, new_AGEMA_signal_1460, SubCellInst_SboxInst_3_n15}), .b ({new_AGEMA_signal_1888, new_AGEMA_signal_1887, new_AGEMA_signal_1886, SubCellInst_SboxInst_3_n12}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_2116, new_AGEMA_signal_2115, new_AGEMA_signal_2114, Feedback[14]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U8 ( .a ({new_AGEMA_signal_1474, new_AGEMA_signal_1473, new_AGEMA_signal_1472, SubCellInst_SboxInst_3_n13}), .b ({new_AGEMA_signal_1894, new_AGEMA_signal_1893, new_AGEMA_signal_1892, SubCellInst_SboxInst_3_n3}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_2122, new_AGEMA_signal_2121, new_AGEMA_signal_2120, Feedback[12]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U17 ( .a ({new_AGEMA_signal_1480, new_AGEMA_signal_1479, new_AGEMA_signal_1478, SubCellInst_SboxInst_4_n15}), .b ({new_AGEMA_signal_1903, new_AGEMA_signal_1902, new_AGEMA_signal_1901, SubCellInst_SboxInst_4_n12}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_2128, new_AGEMA_signal_2127, new_AGEMA_signal_2126, Feedback[18]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U8 ( .a ({new_AGEMA_signal_1492, new_AGEMA_signal_1491, new_AGEMA_signal_1490, SubCellInst_SboxInst_4_n13}), .b ({new_AGEMA_signal_1909, new_AGEMA_signal_1908, new_AGEMA_signal_1907, SubCellInst_SboxInst_4_n3}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_2134, new_AGEMA_signal_2133, new_AGEMA_signal_2132, Feedback[16]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U17 ( .a ({new_AGEMA_signal_1498, new_AGEMA_signal_1497, new_AGEMA_signal_1496, SubCellInst_SboxInst_5_n15}), .b ({new_AGEMA_signal_1918, new_AGEMA_signal_1917, new_AGEMA_signal_1916, SubCellInst_SboxInst_5_n12}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_2140, new_AGEMA_signal_2139, new_AGEMA_signal_2138, Feedback[22]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U8 ( .a ({new_AGEMA_signal_1510, new_AGEMA_signal_1509, new_AGEMA_signal_1508, SubCellInst_SboxInst_5_n13}), .b ({new_AGEMA_signal_1924, new_AGEMA_signal_1923, new_AGEMA_signal_1922, SubCellInst_SboxInst_5_n3}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_2146, new_AGEMA_signal_2145, new_AGEMA_signal_2144, Feedback[20]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U17 ( .a ({new_AGEMA_signal_1516, new_AGEMA_signal_1515, new_AGEMA_signal_1514, SubCellInst_SboxInst_6_n15}), .b ({new_AGEMA_signal_1933, new_AGEMA_signal_1932, new_AGEMA_signal_1931, SubCellInst_SboxInst_6_n12}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_2152, new_AGEMA_signal_2151, new_AGEMA_signal_2150, Feedback[26]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U8 ( .a ({new_AGEMA_signal_1528, new_AGEMA_signal_1527, new_AGEMA_signal_1526, SubCellInst_SboxInst_6_n13}), .b ({new_AGEMA_signal_1939, new_AGEMA_signal_1938, new_AGEMA_signal_1937, SubCellInst_SboxInst_6_n3}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_2158, new_AGEMA_signal_2157, new_AGEMA_signal_2156, Feedback[24]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U17 ( .a ({new_AGEMA_signal_1534, new_AGEMA_signal_1533, new_AGEMA_signal_1532, SubCellInst_SboxInst_7_n15}), .b ({new_AGEMA_signal_1948, new_AGEMA_signal_1947, new_AGEMA_signal_1946, SubCellInst_SboxInst_7_n12}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_2164, new_AGEMA_signal_2163, new_AGEMA_signal_2162, Feedback[30]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U8 ( .a ({new_AGEMA_signal_1546, new_AGEMA_signal_1545, new_AGEMA_signal_1544, SubCellInst_SboxInst_7_n13}), .b ({new_AGEMA_signal_1954, new_AGEMA_signal_1953, new_AGEMA_signal_1952, SubCellInst_SboxInst_7_n3}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_2170, new_AGEMA_signal_2169, new_AGEMA_signal_2168, Feedback[28]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U17 ( .a ({new_AGEMA_signal_1552, new_AGEMA_signal_1551, new_AGEMA_signal_1550, SubCellInst_SboxInst_8_n15}), .b ({new_AGEMA_signal_1963, new_AGEMA_signal_1962, new_AGEMA_signal_1961, SubCellInst_SboxInst_8_n12}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_2176, new_AGEMA_signal_2175, new_AGEMA_signal_2174, Feedback[34]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U8 ( .a ({new_AGEMA_signal_1564, new_AGEMA_signal_1563, new_AGEMA_signal_1562, SubCellInst_SboxInst_8_n13}), .b ({new_AGEMA_signal_1969, new_AGEMA_signal_1968, new_AGEMA_signal_1967, SubCellInst_SboxInst_8_n3}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_2182, new_AGEMA_signal_2181, new_AGEMA_signal_2180, Feedback[32]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U17 ( .a ({new_AGEMA_signal_1570, new_AGEMA_signal_1569, new_AGEMA_signal_1568, SubCellInst_SboxInst_9_n15}), .b ({new_AGEMA_signal_1978, new_AGEMA_signal_1977, new_AGEMA_signal_1976, SubCellInst_SboxInst_9_n12}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_2188, new_AGEMA_signal_2187, new_AGEMA_signal_2186, Feedback[38]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U8 ( .a ({new_AGEMA_signal_1582, new_AGEMA_signal_1581, new_AGEMA_signal_1580, SubCellInst_SboxInst_9_n13}), .b ({new_AGEMA_signal_1984, new_AGEMA_signal_1983, new_AGEMA_signal_1982, SubCellInst_SboxInst_9_n3}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_2194, new_AGEMA_signal_2193, new_AGEMA_signal_2192, Feedback[36]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U17 ( .a ({new_AGEMA_signal_1588, new_AGEMA_signal_1587, new_AGEMA_signal_1586, SubCellInst_SboxInst_10_n15}), .b ({new_AGEMA_signal_1993, new_AGEMA_signal_1992, new_AGEMA_signal_1991, SubCellInst_SboxInst_10_n12}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_2200, new_AGEMA_signal_2199, new_AGEMA_signal_2198, Feedback[42]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U8 ( .a ({new_AGEMA_signal_1600, new_AGEMA_signal_1599, new_AGEMA_signal_1598, SubCellInst_SboxInst_10_n13}), .b ({new_AGEMA_signal_1999, new_AGEMA_signal_1998, new_AGEMA_signal_1997, SubCellInst_SboxInst_10_n3}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_2206, new_AGEMA_signal_2205, new_AGEMA_signal_2204, Feedback[40]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U17 ( .a ({new_AGEMA_signal_1606, new_AGEMA_signal_1605, new_AGEMA_signal_1604, SubCellInst_SboxInst_11_n15}), .b ({new_AGEMA_signal_2008, new_AGEMA_signal_2007, new_AGEMA_signal_2006, SubCellInst_SboxInst_11_n12}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_2212, new_AGEMA_signal_2211, new_AGEMA_signal_2210, Feedback[46]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U8 ( .a ({new_AGEMA_signal_1618, new_AGEMA_signal_1617, new_AGEMA_signal_1616, SubCellInst_SboxInst_11_n13}), .b ({new_AGEMA_signal_2014, new_AGEMA_signal_2013, new_AGEMA_signal_2012, SubCellInst_SboxInst_11_n3}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_2218, new_AGEMA_signal_2217, new_AGEMA_signal_2216, Feedback[44]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U17 ( .a ({new_AGEMA_signal_1624, new_AGEMA_signal_1623, new_AGEMA_signal_1622, SubCellInst_SboxInst_12_n15}), .b ({new_AGEMA_signal_2023, new_AGEMA_signal_2022, new_AGEMA_signal_2021, SubCellInst_SboxInst_12_n12}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_2224, new_AGEMA_signal_2223, new_AGEMA_signal_2222, Feedback[50]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U8 ( .a ({new_AGEMA_signal_1636, new_AGEMA_signal_1635, new_AGEMA_signal_1634, SubCellInst_SboxInst_12_n13}), .b ({new_AGEMA_signal_2029, new_AGEMA_signal_2028, new_AGEMA_signal_2027, SubCellInst_SboxInst_12_n3}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_2230, new_AGEMA_signal_2229, new_AGEMA_signal_2228, Feedback[48]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U17 ( .a ({new_AGEMA_signal_1642, new_AGEMA_signal_1641, new_AGEMA_signal_1640, SubCellInst_SboxInst_13_n15}), .b ({new_AGEMA_signal_2038, new_AGEMA_signal_2037, new_AGEMA_signal_2036, SubCellInst_SboxInst_13_n12}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_2236, new_AGEMA_signal_2235, new_AGEMA_signal_2234, Feedback[54]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U8 ( .a ({new_AGEMA_signal_1654, new_AGEMA_signal_1653, new_AGEMA_signal_1652, SubCellInst_SboxInst_13_n13}), .b ({new_AGEMA_signal_2044, new_AGEMA_signal_2043, new_AGEMA_signal_2042, SubCellInst_SboxInst_13_n3}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_2242, new_AGEMA_signal_2241, new_AGEMA_signal_2240, Feedback[52]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U17 ( .a ({new_AGEMA_signal_1660, new_AGEMA_signal_1659, new_AGEMA_signal_1658, SubCellInst_SboxInst_14_n15}), .b ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, new_AGEMA_signal_2051, SubCellInst_SboxInst_14_n12}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_2248, new_AGEMA_signal_2247, new_AGEMA_signal_2246, Feedback[58]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U8 ( .a ({new_AGEMA_signal_1672, new_AGEMA_signal_1671, new_AGEMA_signal_1670, SubCellInst_SboxInst_14_n13}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, new_AGEMA_signal_2057, SubCellInst_SboxInst_14_n3}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_2254, new_AGEMA_signal_2253, new_AGEMA_signal_2252, Feedback[56]}) ) ;
    nand_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U17 ( .a ({new_AGEMA_signal_1678, new_AGEMA_signal_1677, new_AGEMA_signal_1676, SubCellInst_SboxInst_15_n15}), .b ({new_AGEMA_signal_2068, new_AGEMA_signal_2067, new_AGEMA_signal_2066, SubCellInst_SboxInst_15_n12}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_2260, new_AGEMA_signal_2259, new_AGEMA_signal_2258, Feedback[62]}) ) ;
    nor_HPC2 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U8 ( .a ({new_AGEMA_signal_1690, new_AGEMA_signal_1689, new_AGEMA_signal_1688, SubCellInst_SboxInst_15_n13}), .b ({new_AGEMA_signal_2074, new_AGEMA_signal_2073, new_AGEMA_signal_2072, SubCellInst_SboxInst_15_n3}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_2266, new_AGEMA_signal_2265, new_AGEMA_signal_2264, Feedback[60]}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3682, new_AGEMA_signal_3681, new_AGEMA_signal_3680, AddRoundKeyOutput[63]}), .Q ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, new_AGEMA_signal_3677, AddRoundKeyOutput[62]}), .Q ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3676, new_AGEMA_signal_3675, new_AGEMA_signal_3674, AddRoundKeyOutput[61]}), .Q ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, new_AGEMA_signal_3671, AddRoundKeyOutput[60]}), .Q ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3670, new_AGEMA_signal_3669, new_AGEMA_signal_3668, AddRoundKeyOutput[59]}), .Q ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, new_AGEMA_signal_3665, AddRoundKeyOutput[58]}), .Q ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3664, new_AGEMA_signal_3663, new_AGEMA_signal_3662, AddRoundKeyOutput[57]}), .Q ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, new_AGEMA_signal_3659, AddRoundKeyOutput[56]}), .Q ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3658, new_AGEMA_signal_3657, new_AGEMA_signal_3656, AddRoundKeyOutput[55]}), .Q ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, new_AGEMA_signal_3653, AddRoundKeyOutput[54]}), .Q ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3652, new_AGEMA_signal_3651, new_AGEMA_signal_3650, AddRoundKeyOutput[53]}), .Q ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, new_AGEMA_signal_3647, AddRoundKeyOutput[52]}), .Q ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3646, new_AGEMA_signal_3645, new_AGEMA_signal_3644, AddRoundKeyOutput[51]}), .Q ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, new_AGEMA_signal_3641, AddRoundKeyOutput[50]}), .Q ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3640, new_AGEMA_signal_3639, new_AGEMA_signal_3638, AddRoundKeyOutput[49]}), .Q ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, new_AGEMA_signal_3635, AddRoundKeyOutput[48]}), .Q ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3706, new_AGEMA_signal_3705, new_AGEMA_signal_3704, AddRoundKeyOutput[47]}), .Q ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, new_AGEMA_signal_3701, AddRoundKeyOutput[46]}), .Q ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3700, new_AGEMA_signal_3699, new_AGEMA_signal_3698, AddRoundKeyOutput[45]}), .Q ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, new_AGEMA_signal_3695, AddRoundKeyOutput[44]}), .Q ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3694, new_AGEMA_signal_3693, new_AGEMA_signal_3692, AddRoundKeyOutput[43]}), .Q ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, new_AGEMA_signal_3689, AddRoundKeyOutput[42]}), .Q ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3688, new_AGEMA_signal_3687, new_AGEMA_signal_3686, AddRoundKeyOutput[41]}), .Q ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, new_AGEMA_signal_3683, AddRoundKeyOutput[40]}), .Q ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3730, new_AGEMA_signal_3729, new_AGEMA_signal_3728, AddRoundKeyOutput[39]}), .Q ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, new_AGEMA_signal_3725, AddRoundKeyOutput[38]}), .Q ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3724, new_AGEMA_signal_3723, new_AGEMA_signal_3722, AddRoundKeyOutput[37]}), .Q ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, new_AGEMA_signal_3719, AddRoundKeyOutput[36]}), .Q ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3718, new_AGEMA_signal_3717, new_AGEMA_signal_3716, AddRoundKeyOutput[35]}), .Q ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, new_AGEMA_signal_3713, AddRoundKeyOutput[34]}), .Q ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3712, new_AGEMA_signal_3711, new_AGEMA_signal_3710, AddRoundKeyOutput[33]}), .Q ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, new_AGEMA_signal_3707, AddRoundKeyOutput[32]}), .Q ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3538, new_AGEMA_signal_3537, new_AGEMA_signal_3536, AddRoundKeyOutput[31]}), .Q ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, new_AGEMA_signal_3533, AddRoundKeyOutput[30]}), .Q ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3532, new_AGEMA_signal_3531, new_AGEMA_signal_3530, AddRoundKeyOutput[29]}), .Q ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, new_AGEMA_signal_3527, AddRoundKeyOutput[28]}), .Q ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3526, new_AGEMA_signal_3525, new_AGEMA_signal_3524, AddRoundKeyOutput[27]}), .Q ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, new_AGEMA_signal_3521, AddRoundKeyOutput[26]}), .Q ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3520, new_AGEMA_signal_3519, new_AGEMA_signal_3518, AddRoundKeyOutput[25]}), .Q ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, new_AGEMA_signal_3515, AddRoundKeyOutput[24]}), .Q ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3514, new_AGEMA_signal_3513, new_AGEMA_signal_3512, AddRoundKeyOutput[23]}), .Q ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, new_AGEMA_signal_3509, AddRoundKeyOutput[22]}), .Q ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3508, new_AGEMA_signal_3507, new_AGEMA_signal_3506, AddRoundKeyOutput[21]}), .Q ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, new_AGEMA_signal_3503, AddRoundKeyOutput[20]}), .Q ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3502, new_AGEMA_signal_3501, new_AGEMA_signal_3500, AddRoundKeyOutput[19]}), .Q ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, new_AGEMA_signal_3497, AddRoundKeyOutput[18]}), .Q ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3496, new_AGEMA_signal_3495, new_AGEMA_signal_3494, AddRoundKeyOutput[17]}), .Q ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, new_AGEMA_signal_3491, AddRoundKeyOutput[16]}), .Q ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3490, new_AGEMA_signal_3489, new_AGEMA_signal_3488, AddRoundKeyOutput[15]}), .Q ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, new_AGEMA_signal_3485, AddRoundKeyOutput[14]}), .Q ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3484, new_AGEMA_signal_3483, new_AGEMA_signal_3482, AddRoundKeyOutput[13]}), .Q ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, new_AGEMA_signal_3479, AddRoundKeyOutput[12]}), .Q ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3478, new_AGEMA_signal_3477, new_AGEMA_signal_3476, AddRoundKeyOutput[11]}), .Q ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, new_AGEMA_signal_3473, AddRoundKeyOutput[10]}), .Q ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3472, new_AGEMA_signal_3471, new_AGEMA_signal_3470, AddRoundKeyOutput[9]}), .Q ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, new_AGEMA_signal_3467, AddRoundKeyOutput[8]}), .Q ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3466, new_AGEMA_signal_3465, new_AGEMA_signal_3464, AddRoundKeyOutput[7]}), .Q ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, new_AGEMA_signal_3461, AddRoundKeyOutput[6]}), .Q ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3460, new_AGEMA_signal_3459, new_AGEMA_signal_3458, AddRoundKeyOutput[5]}), .Q ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, new_AGEMA_signal_3455, AddRoundKeyOutput[4]}), .Q ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3454, new_AGEMA_signal_3453, new_AGEMA_signal_3452, AddRoundKeyOutput[3]}), .Q ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, new_AGEMA_signal_3449, AddRoundKeyOutput[2]}), .Q ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3448, new_AGEMA_signal_3447, new_AGEMA_signal_3446, AddRoundKeyOutput[1]}), .Q ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, new_AGEMA_signal_3443, AddRoundKeyOutput[0]}), .Q ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_6__FF_FF ( .CK (clk_gated), .D (FSMUpdate[6]), .Q (FSMReg[6]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (FSMUpdate[5]), .Q (FSMReg[5]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (FSMUpdate[4]), .Q (FSMReg[4]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (FSMUpdate[3]), .Q (FSMReg[3]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (FSMUpdate[2]), .Q (FSMReg[2]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (FSMUpdate[1]), .Q (FSMReg[1]), .QN () ) ;
    DFF_X1 FSMRegInst_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (FSMUpdate[0]), .Q (FSMReg[0]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (selectsNext[1]), .Q (selectsReg[1]), .QN () ) ;
    DFF_X1 selectsRegInst_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (selectsNext[0]), .Q (selectsReg[0]), .QN () ) ;
    DFF_X1 done_reg_FF_FF ( .CK (clk_gated), .D (done_internal), .Q (done), .QN () ) ;
endmodule
