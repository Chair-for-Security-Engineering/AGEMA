/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module LED_HPC2_Pipeline_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    wire n15 ;
    wire n14 ;
    wire n16 ;
    wire n17 ;
    wire n18 ;
    wire n19 ;
    wire n20 ;
    wire LED_128_Instance_n34 ;
    wire LED_128_Instance_n33 ;
    wire LED_128_Instance_n32 ;
    wire LED_128_Instance_n23 ;
    wire LED_128_Instance_n21 ;
    wire LED_128_Instance_n20 ;
    wire LED_128_Instance_n19 ;
    wire LED_128_Instance_n18 ;
    wire LED_128_Instance_n17 ;
    wire LED_128_Instance_n16 ;
    wire LED_128_Instance_n15 ;
    wire LED_128_Instance_n14 ;
    wire LED_128_Instance_n13 ;
    wire LED_128_Instance_n12 ;
    wire LED_128_Instance_n11 ;
    wire LED_128_Instance_n10 ;
    wire LED_128_Instance_n2 ;
    wire LED_128_Instance_n1 ;
    wire LED_128_Instance_n27 ;
    wire LED_128_Instance_N9 ;
    wire LED_128_Instance_n28 ;
    wire LED_128_Instance_N8 ;
    wire LED_128_Instance_n30 ;
    wire LED_128_Instance_N7 ;
    wire LED_128_Instance_n5 ;
    wire LED_128_Instance_N6 ;
    wire LED_128_Instance_n29 ;
    wire LED_128_Instance_N5 ;
    wire LED_128_Instance_n6 ;
    wire LED_128_Instance_N4 ;
    wire LED_128_Instance_n24 ;
    wire LED_128_Instance_N13 ;
    wire LED_128_Instance_n25 ;
    wire LED_128_Instance_N12 ;
    wire LED_128_Instance_n8 ;
    wire LED_128_Instance_n26 ;
    wire LED_128_Instance_N11 ;
    wire LED_128_Instance_n4 ;
    wire LED_128_Instance_N10 ;
    wire LED_128_Instance_n31 ;
    wire LED_128_Instance_addroundkey_out_0_ ;
    wire LED_128_Instance_addroundkey_out_1_ ;
    wire LED_128_Instance_addroundkey_out_2_ ;
    wire LED_128_Instance_addroundkey_out_3_ ;
    wire LED_128_Instance_addroundkey_out_4_ ;
    wire LED_128_Instance_addroundkey_out_5_ ;
    wire LED_128_Instance_addroundkey_out_6_ ;
    wire LED_128_Instance_addroundkey_out_16_ ;
    wire LED_128_Instance_addroundkey_out_17_ ;
    wire LED_128_Instance_addroundkey_out_18_ ;
    wire LED_128_Instance_addroundkey_out_19_ ;
    wire LED_128_Instance_addroundkey_out_20_ ;
    wire LED_128_Instance_addroundkey_out_21_ ;
    wire LED_128_Instance_addroundkey_out_22_ ;
    wire LED_128_Instance_addroundkey_out_32_ ;
    wire LED_128_Instance_addroundkey_out_33_ ;
    wire LED_128_Instance_addroundkey_out_34_ ;
    wire LED_128_Instance_addroundkey_out_35_ ;
    wire LED_128_Instance_addroundkey_out_36_ ;
    wire LED_128_Instance_addroundkey_out_37_ ;
    wire LED_128_Instance_addroundkey_out_38_ ;
    wire LED_128_Instance_addroundkey_out_48_ ;
    wire LED_128_Instance_addroundkey_out_49_ ;
    wire LED_128_Instance_addroundkey_out_50_ ;
    wire LED_128_Instance_addroundkey_out_51_ ;
    wire LED_128_Instance_addroundkey_out_52_ ;
    wire LED_128_Instance_addroundkey_out_53_ ;
    wire LED_128_Instance_addroundkey_out_54_ ;
    wire LED_128_Instance_n22 ;
    wire LED_128_Instance_MUX_state0_n11 ;
    wire LED_128_Instance_MUX_state0_n10 ;
    wire LED_128_Instance_MUX_state0_n9 ;
    wire LED_128_Instance_MUX_state0_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n10 ;
    wire LED_128_Instance_MUX_current_roundkey_n9 ;
    wire LED_128_Instance_MUX_current_roundkey_n8 ;
    wire LED_128_Instance_MUX_current_roundkey_n7 ;
    wire LED_128_Instance_MUX_addroundkey_out_n9 ;
    wire LED_128_Instance_MUX_addroundkey_out_n8 ;
    wire LED_128_Instance_MUX_addroundkey_out_n7 ;
    wire LED_128_Instance_SBox_Instance_0_n3 ;
    wire LED_128_Instance_SBox_Instance_0_n2 ;
    wire LED_128_Instance_SBox_Instance_0_n1 ;
    wire LED_128_Instance_SBox_Instance_0_L8 ;
    wire LED_128_Instance_SBox_Instance_0_L7 ;
    wire LED_128_Instance_SBox_Instance_0_T3 ;
    wire LED_128_Instance_SBox_Instance_0_T1 ;
    wire LED_128_Instance_SBox_Instance_0_Q7 ;
    wire LED_128_Instance_SBox_Instance_0_Q6 ;
    wire LED_128_Instance_SBox_Instance_0_L5 ;
    wire LED_128_Instance_SBox_Instance_0_T2 ;
    wire LED_128_Instance_SBox_Instance_0_L4 ;
    wire LED_128_Instance_SBox_Instance_0_Q3 ;
    wire LED_128_Instance_SBox_Instance_0_L3 ;
    wire LED_128_Instance_SBox_Instance_0_Q2 ;
    wire LED_128_Instance_SBox_Instance_0_T0 ;
    wire LED_128_Instance_SBox_Instance_0_L2 ;
    wire LED_128_Instance_SBox_Instance_0_L1 ;
    wire LED_128_Instance_SBox_Instance_0_L0 ;
    wire LED_128_Instance_SBox_Instance_1_n3 ;
    wire LED_128_Instance_SBox_Instance_1_n2 ;
    wire LED_128_Instance_SBox_Instance_1_n1 ;
    wire LED_128_Instance_SBox_Instance_1_L8 ;
    wire LED_128_Instance_SBox_Instance_1_L7 ;
    wire LED_128_Instance_SBox_Instance_1_T3 ;
    wire LED_128_Instance_SBox_Instance_1_T1 ;
    wire LED_128_Instance_SBox_Instance_1_Q7 ;
    wire LED_128_Instance_SBox_Instance_1_Q6 ;
    wire LED_128_Instance_SBox_Instance_1_L5 ;
    wire LED_128_Instance_SBox_Instance_1_T2 ;
    wire LED_128_Instance_SBox_Instance_1_L4 ;
    wire LED_128_Instance_SBox_Instance_1_Q3 ;
    wire LED_128_Instance_SBox_Instance_1_L3 ;
    wire LED_128_Instance_SBox_Instance_1_Q2 ;
    wire LED_128_Instance_SBox_Instance_1_T0 ;
    wire LED_128_Instance_SBox_Instance_1_L2 ;
    wire LED_128_Instance_SBox_Instance_1_L1 ;
    wire LED_128_Instance_SBox_Instance_1_L0 ;
    wire LED_128_Instance_SBox_Instance_2_n3 ;
    wire LED_128_Instance_SBox_Instance_2_n2 ;
    wire LED_128_Instance_SBox_Instance_2_n1 ;
    wire LED_128_Instance_SBox_Instance_2_L8 ;
    wire LED_128_Instance_SBox_Instance_2_L7 ;
    wire LED_128_Instance_SBox_Instance_2_T3 ;
    wire LED_128_Instance_SBox_Instance_2_T1 ;
    wire LED_128_Instance_SBox_Instance_2_Q7 ;
    wire LED_128_Instance_SBox_Instance_2_Q6 ;
    wire LED_128_Instance_SBox_Instance_2_L5 ;
    wire LED_128_Instance_SBox_Instance_2_T2 ;
    wire LED_128_Instance_SBox_Instance_2_L4 ;
    wire LED_128_Instance_SBox_Instance_2_Q3 ;
    wire LED_128_Instance_SBox_Instance_2_L3 ;
    wire LED_128_Instance_SBox_Instance_2_Q2 ;
    wire LED_128_Instance_SBox_Instance_2_T0 ;
    wire LED_128_Instance_SBox_Instance_2_L2 ;
    wire LED_128_Instance_SBox_Instance_2_L1 ;
    wire LED_128_Instance_SBox_Instance_2_L0 ;
    wire LED_128_Instance_SBox_Instance_3_n3 ;
    wire LED_128_Instance_SBox_Instance_3_n2 ;
    wire LED_128_Instance_SBox_Instance_3_n1 ;
    wire LED_128_Instance_SBox_Instance_3_L8 ;
    wire LED_128_Instance_SBox_Instance_3_L7 ;
    wire LED_128_Instance_SBox_Instance_3_T3 ;
    wire LED_128_Instance_SBox_Instance_3_T1 ;
    wire LED_128_Instance_SBox_Instance_3_Q7 ;
    wire LED_128_Instance_SBox_Instance_3_Q6 ;
    wire LED_128_Instance_SBox_Instance_3_L5 ;
    wire LED_128_Instance_SBox_Instance_3_T2 ;
    wire LED_128_Instance_SBox_Instance_3_L4 ;
    wire LED_128_Instance_SBox_Instance_3_Q3 ;
    wire LED_128_Instance_SBox_Instance_3_L3 ;
    wire LED_128_Instance_SBox_Instance_3_Q2 ;
    wire LED_128_Instance_SBox_Instance_3_T0 ;
    wire LED_128_Instance_SBox_Instance_3_L2 ;
    wire LED_128_Instance_SBox_Instance_3_L1 ;
    wire LED_128_Instance_SBox_Instance_3_L0 ;
    wire LED_128_Instance_SBox_Instance_4_n3 ;
    wire LED_128_Instance_SBox_Instance_4_n2 ;
    wire LED_128_Instance_SBox_Instance_4_n1 ;
    wire LED_128_Instance_SBox_Instance_4_L8 ;
    wire LED_128_Instance_SBox_Instance_4_L7 ;
    wire LED_128_Instance_SBox_Instance_4_T3 ;
    wire LED_128_Instance_SBox_Instance_4_T1 ;
    wire LED_128_Instance_SBox_Instance_4_Q7 ;
    wire LED_128_Instance_SBox_Instance_4_Q6 ;
    wire LED_128_Instance_SBox_Instance_4_L5 ;
    wire LED_128_Instance_SBox_Instance_4_T2 ;
    wire LED_128_Instance_SBox_Instance_4_L4 ;
    wire LED_128_Instance_SBox_Instance_4_Q3 ;
    wire LED_128_Instance_SBox_Instance_4_L3 ;
    wire LED_128_Instance_SBox_Instance_4_Q2 ;
    wire LED_128_Instance_SBox_Instance_4_T0 ;
    wire LED_128_Instance_SBox_Instance_4_L2 ;
    wire LED_128_Instance_SBox_Instance_4_L1 ;
    wire LED_128_Instance_SBox_Instance_4_L0 ;
    wire LED_128_Instance_SBox_Instance_5_n3 ;
    wire LED_128_Instance_SBox_Instance_5_n2 ;
    wire LED_128_Instance_SBox_Instance_5_n1 ;
    wire LED_128_Instance_SBox_Instance_5_L8 ;
    wire LED_128_Instance_SBox_Instance_5_L7 ;
    wire LED_128_Instance_SBox_Instance_5_T3 ;
    wire LED_128_Instance_SBox_Instance_5_T1 ;
    wire LED_128_Instance_SBox_Instance_5_Q7 ;
    wire LED_128_Instance_SBox_Instance_5_Q6 ;
    wire LED_128_Instance_SBox_Instance_5_L5 ;
    wire LED_128_Instance_SBox_Instance_5_T2 ;
    wire LED_128_Instance_SBox_Instance_5_L4 ;
    wire LED_128_Instance_SBox_Instance_5_Q3 ;
    wire LED_128_Instance_SBox_Instance_5_L3 ;
    wire LED_128_Instance_SBox_Instance_5_Q2 ;
    wire LED_128_Instance_SBox_Instance_5_T0 ;
    wire LED_128_Instance_SBox_Instance_5_L2 ;
    wire LED_128_Instance_SBox_Instance_5_L1 ;
    wire LED_128_Instance_SBox_Instance_5_L0 ;
    wire LED_128_Instance_SBox_Instance_6_n3 ;
    wire LED_128_Instance_SBox_Instance_6_n2 ;
    wire LED_128_Instance_SBox_Instance_6_n1 ;
    wire LED_128_Instance_SBox_Instance_6_L8 ;
    wire LED_128_Instance_SBox_Instance_6_L7 ;
    wire LED_128_Instance_SBox_Instance_6_T3 ;
    wire LED_128_Instance_SBox_Instance_6_T1 ;
    wire LED_128_Instance_SBox_Instance_6_Q7 ;
    wire LED_128_Instance_SBox_Instance_6_Q6 ;
    wire LED_128_Instance_SBox_Instance_6_L5 ;
    wire LED_128_Instance_SBox_Instance_6_T2 ;
    wire LED_128_Instance_SBox_Instance_6_L4 ;
    wire LED_128_Instance_SBox_Instance_6_Q3 ;
    wire LED_128_Instance_SBox_Instance_6_L3 ;
    wire LED_128_Instance_SBox_Instance_6_Q2 ;
    wire LED_128_Instance_SBox_Instance_6_T0 ;
    wire LED_128_Instance_SBox_Instance_6_L2 ;
    wire LED_128_Instance_SBox_Instance_6_L1 ;
    wire LED_128_Instance_SBox_Instance_6_L0 ;
    wire LED_128_Instance_SBox_Instance_7_n3 ;
    wire LED_128_Instance_SBox_Instance_7_n2 ;
    wire LED_128_Instance_SBox_Instance_7_n1 ;
    wire LED_128_Instance_SBox_Instance_7_L8 ;
    wire LED_128_Instance_SBox_Instance_7_L7 ;
    wire LED_128_Instance_SBox_Instance_7_T3 ;
    wire LED_128_Instance_SBox_Instance_7_T1 ;
    wire LED_128_Instance_SBox_Instance_7_Q7 ;
    wire LED_128_Instance_SBox_Instance_7_Q6 ;
    wire LED_128_Instance_SBox_Instance_7_L5 ;
    wire LED_128_Instance_SBox_Instance_7_T2 ;
    wire LED_128_Instance_SBox_Instance_7_L4 ;
    wire LED_128_Instance_SBox_Instance_7_Q3 ;
    wire LED_128_Instance_SBox_Instance_7_L3 ;
    wire LED_128_Instance_SBox_Instance_7_Q2 ;
    wire LED_128_Instance_SBox_Instance_7_T0 ;
    wire LED_128_Instance_SBox_Instance_7_L2 ;
    wire LED_128_Instance_SBox_Instance_7_L1 ;
    wire LED_128_Instance_SBox_Instance_7_L0 ;
    wire LED_128_Instance_SBox_Instance_8_n3 ;
    wire LED_128_Instance_SBox_Instance_8_n2 ;
    wire LED_128_Instance_SBox_Instance_8_n1 ;
    wire LED_128_Instance_SBox_Instance_8_L8 ;
    wire LED_128_Instance_SBox_Instance_8_L7 ;
    wire LED_128_Instance_SBox_Instance_8_T3 ;
    wire LED_128_Instance_SBox_Instance_8_T1 ;
    wire LED_128_Instance_SBox_Instance_8_Q7 ;
    wire LED_128_Instance_SBox_Instance_8_Q6 ;
    wire LED_128_Instance_SBox_Instance_8_L5 ;
    wire LED_128_Instance_SBox_Instance_8_T2 ;
    wire LED_128_Instance_SBox_Instance_8_L4 ;
    wire LED_128_Instance_SBox_Instance_8_Q3 ;
    wire LED_128_Instance_SBox_Instance_8_L3 ;
    wire LED_128_Instance_SBox_Instance_8_Q2 ;
    wire LED_128_Instance_SBox_Instance_8_T0 ;
    wire LED_128_Instance_SBox_Instance_8_L2 ;
    wire LED_128_Instance_SBox_Instance_8_L1 ;
    wire LED_128_Instance_SBox_Instance_8_L0 ;
    wire LED_128_Instance_SBox_Instance_9_n3 ;
    wire LED_128_Instance_SBox_Instance_9_n2 ;
    wire LED_128_Instance_SBox_Instance_9_n1 ;
    wire LED_128_Instance_SBox_Instance_9_L8 ;
    wire LED_128_Instance_SBox_Instance_9_L7 ;
    wire LED_128_Instance_SBox_Instance_9_T3 ;
    wire LED_128_Instance_SBox_Instance_9_T1 ;
    wire LED_128_Instance_SBox_Instance_9_Q7 ;
    wire LED_128_Instance_SBox_Instance_9_Q6 ;
    wire LED_128_Instance_SBox_Instance_9_L5 ;
    wire LED_128_Instance_SBox_Instance_9_T2 ;
    wire LED_128_Instance_SBox_Instance_9_L4 ;
    wire LED_128_Instance_SBox_Instance_9_Q3 ;
    wire LED_128_Instance_SBox_Instance_9_L3 ;
    wire LED_128_Instance_SBox_Instance_9_Q2 ;
    wire LED_128_Instance_SBox_Instance_9_T0 ;
    wire LED_128_Instance_SBox_Instance_9_L2 ;
    wire LED_128_Instance_SBox_Instance_9_L1 ;
    wire LED_128_Instance_SBox_Instance_9_L0 ;
    wire LED_128_Instance_SBox_Instance_10_n3 ;
    wire LED_128_Instance_SBox_Instance_10_n2 ;
    wire LED_128_Instance_SBox_Instance_10_n1 ;
    wire LED_128_Instance_SBox_Instance_10_L8 ;
    wire LED_128_Instance_SBox_Instance_10_L7 ;
    wire LED_128_Instance_SBox_Instance_10_T3 ;
    wire LED_128_Instance_SBox_Instance_10_T1 ;
    wire LED_128_Instance_SBox_Instance_10_Q7 ;
    wire LED_128_Instance_SBox_Instance_10_Q6 ;
    wire LED_128_Instance_SBox_Instance_10_L5 ;
    wire LED_128_Instance_SBox_Instance_10_T2 ;
    wire LED_128_Instance_SBox_Instance_10_L4 ;
    wire LED_128_Instance_SBox_Instance_10_Q3 ;
    wire LED_128_Instance_SBox_Instance_10_L3 ;
    wire LED_128_Instance_SBox_Instance_10_Q2 ;
    wire LED_128_Instance_SBox_Instance_10_T0 ;
    wire LED_128_Instance_SBox_Instance_10_L2 ;
    wire LED_128_Instance_SBox_Instance_10_L1 ;
    wire LED_128_Instance_SBox_Instance_10_L0 ;
    wire LED_128_Instance_SBox_Instance_11_n3 ;
    wire LED_128_Instance_SBox_Instance_11_n2 ;
    wire LED_128_Instance_SBox_Instance_11_n1 ;
    wire LED_128_Instance_SBox_Instance_11_L8 ;
    wire LED_128_Instance_SBox_Instance_11_L7 ;
    wire LED_128_Instance_SBox_Instance_11_T3 ;
    wire LED_128_Instance_SBox_Instance_11_T1 ;
    wire LED_128_Instance_SBox_Instance_11_Q7 ;
    wire LED_128_Instance_SBox_Instance_11_Q6 ;
    wire LED_128_Instance_SBox_Instance_11_L5 ;
    wire LED_128_Instance_SBox_Instance_11_T2 ;
    wire LED_128_Instance_SBox_Instance_11_L4 ;
    wire LED_128_Instance_SBox_Instance_11_Q3 ;
    wire LED_128_Instance_SBox_Instance_11_L3 ;
    wire LED_128_Instance_SBox_Instance_11_Q2 ;
    wire LED_128_Instance_SBox_Instance_11_T0 ;
    wire LED_128_Instance_SBox_Instance_11_L2 ;
    wire LED_128_Instance_SBox_Instance_11_L1 ;
    wire LED_128_Instance_SBox_Instance_11_L0 ;
    wire LED_128_Instance_SBox_Instance_12_n3 ;
    wire LED_128_Instance_SBox_Instance_12_n2 ;
    wire LED_128_Instance_SBox_Instance_12_n1 ;
    wire LED_128_Instance_SBox_Instance_12_L8 ;
    wire LED_128_Instance_SBox_Instance_12_L7 ;
    wire LED_128_Instance_SBox_Instance_12_T3 ;
    wire LED_128_Instance_SBox_Instance_12_T1 ;
    wire LED_128_Instance_SBox_Instance_12_Q7 ;
    wire LED_128_Instance_SBox_Instance_12_Q6 ;
    wire LED_128_Instance_SBox_Instance_12_L5 ;
    wire LED_128_Instance_SBox_Instance_12_T2 ;
    wire LED_128_Instance_SBox_Instance_12_L4 ;
    wire LED_128_Instance_SBox_Instance_12_Q3 ;
    wire LED_128_Instance_SBox_Instance_12_L3 ;
    wire LED_128_Instance_SBox_Instance_12_Q2 ;
    wire LED_128_Instance_SBox_Instance_12_T0 ;
    wire LED_128_Instance_SBox_Instance_12_L2 ;
    wire LED_128_Instance_SBox_Instance_12_L1 ;
    wire LED_128_Instance_SBox_Instance_12_L0 ;
    wire LED_128_Instance_SBox_Instance_13_n3 ;
    wire LED_128_Instance_SBox_Instance_13_n2 ;
    wire LED_128_Instance_SBox_Instance_13_n1 ;
    wire LED_128_Instance_SBox_Instance_13_L8 ;
    wire LED_128_Instance_SBox_Instance_13_L7 ;
    wire LED_128_Instance_SBox_Instance_13_T3 ;
    wire LED_128_Instance_SBox_Instance_13_T1 ;
    wire LED_128_Instance_SBox_Instance_13_Q7 ;
    wire LED_128_Instance_SBox_Instance_13_Q6 ;
    wire LED_128_Instance_SBox_Instance_13_L5 ;
    wire LED_128_Instance_SBox_Instance_13_T2 ;
    wire LED_128_Instance_SBox_Instance_13_L4 ;
    wire LED_128_Instance_SBox_Instance_13_Q3 ;
    wire LED_128_Instance_SBox_Instance_13_L3 ;
    wire LED_128_Instance_SBox_Instance_13_Q2 ;
    wire LED_128_Instance_SBox_Instance_13_T0 ;
    wire LED_128_Instance_SBox_Instance_13_L2 ;
    wire LED_128_Instance_SBox_Instance_13_L1 ;
    wire LED_128_Instance_SBox_Instance_13_L0 ;
    wire LED_128_Instance_SBox_Instance_14_n3 ;
    wire LED_128_Instance_SBox_Instance_14_n2 ;
    wire LED_128_Instance_SBox_Instance_14_n1 ;
    wire LED_128_Instance_SBox_Instance_14_L8 ;
    wire LED_128_Instance_SBox_Instance_14_L7 ;
    wire LED_128_Instance_SBox_Instance_14_T3 ;
    wire LED_128_Instance_SBox_Instance_14_T1 ;
    wire LED_128_Instance_SBox_Instance_14_Q7 ;
    wire LED_128_Instance_SBox_Instance_14_Q6 ;
    wire LED_128_Instance_SBox_Instance_14_L5 ;
    wire LED_128_Instance_SBox_Instance_14_T2 ;
    wire LED_128_Instance_SBox_Instance_14_L4 ;
    wire LED_128_Instance_SBox_Instance_14_Q3 ;
    wire LED_128_Instance_SBox_Instance_14_L3 ;
    wire LED_128_Instance_SBox_Instance_14_Q2 ;
    wire LED_128_Instance_SBox_Instance_14_T0 ;
    wire LED_128_Instance_SBox_Instance_14_L2 ;
    wire LED_128_Instance_SBox_Instance_14_L1 ;
    wire LED_128_Instance_SBox_Instance_14_L0 ;
    wire LED_128_Instance_SBox_Instance_15_n3 ;
    wire LED_128_Instance_SBox_Instance_15_n2 ;
    wire LED_128_Instance_SBox_Instance_15_n1 ;
    wire LED_128_Instance_SBox_Instance_15_L8 ;
    wire LED_128_Instance_SBox_Instance_15_L7 ;
    wire LED_128_Instance_SBox_Instance_15_T3 ;
    wire LED_128_Instance_SBox_Instance_15_T1 ;
    wire LED_128_Instance_SBox_Instance_15_Q7 ;
    wire LED_128_Instance_SBox_Instance_15_Q6 ;
    wire LED_128_Instance_SBox_Instance_15_L5 ;
    wire LED_128_Instance_SBox_Instance_15_T2 ;
    wire LED_128_Instance_SBox_Instance_15_L4 ;
    wire LED_128_Instance_SBox_Instance_15_Q3 ;
    wire LED_128_Instance_SBox_Instance_15_L3 ;
    wire LED_128_Instance_SBox_Instance_15_Q2 ;
    wire LED_128_Instance_SBox_Instance_15_T0 ;
    wire LED_128_Instance_SBox_Instance_15_L2 ;
    wire LED_128_Instance_SBox_Instance_15_L1 ;
    wire LED_128_Instance_SBox_Instance_15_L0 ;
    wire LED_128_Instance_MCS_Instance_0_n38 ;
    wire LED_128_Instance_MCS_Instance_0_n37 ;
    wire LED_128_Instance_MCS_Instance_0_n36 ;
    wire LED_128_Instance_MCS_Instance_0_n35 ;
    wire LED_128_Instance_MCS_Instance_0_n34 ;
    wire LED_128_Instance_MCS_Instance_0_n33 ;
    wire LED_128_Instance_MCS_Instance_0_n32 ;
    wire LED_128_Instance_MCS_Instance_0_n31 ;
    wire LED_128_Instance_MCS_Instance_0_n30 ;
    wire LED_128_Instance_MCS_Instance_0_n29 ;
    wire LED_128_Instance_MCS_Instance_0_n28 ;
    wire LED_128_Instance_MCS_Instance_0_n27 ;
    wire LED_128_Instance_MCS_Instance_0_n26 ;
    wire LED_128_Instance_MCS_Instance_0_n25 ;
    wire LED_128_Instance_MCS_Instance_0_n24 ;
    wire LED_128_Instance_MCS_Instance_0_n23 ;
    wire LED_128_Instance_MCS_Instance_0_n22 ;
    wire LED_128_Instance_MCS_Instance_0_n21 ;
    wire LED_128_Instance_MCS_Instance_0_n20 ;
    wire LED_128_Instance_MCS_Instance_0_n19 ;
    wire LED_128_Instance_MCS_Instance_0_n18 ;
    wire LED_128_Instance_MCS_Instance_0_n17 ;
    wire LED_128_Instance_MCS_Instance_0_n16 ;
    wire LED_128_Instance_MCS_Instance_0_n15 ;
    wire LED_128_Instance_MCS_Instance_0_n14 ;
    wire LED_128_Instance_MCS_Instance_0_n13 ;
    wire LED_128_Instance_MCS_Instance_0_n12 ;
    wire LED_128_Instance_MCS_Instance_0_n11 ;
    wire LED_128_Instance_MCS_Instance_0_n10 ;
    wire LED_128_Instance_MCS_Instance_0_n9 ;
    wire LED_128_Instance_MCS_Instance_0_n8 ;
    wire LED_128_Instance_MCS_Instance_0_n7 ;
    wire LED_128_Instance_MCS_Instance_0_n6 ;
    wire LED_128_Instance_MCS_Instance_0_n5 ;
    wire LED_128_Instance_MCS_Instance_0_n4 ;
    wire LED_128_Instance_MCS_Instance_0_n3 ;
    wire LED_128_Instance_MCS_Instance_0_n2 ;
    wire LED_128_Instance_MCS_Instance_0_n1 ;
    wire LED_128_Instance_MCS_Instance_1_n38 ;
    wire LED_128_Instance_MCS_Instance_1_n37 ;
    wire LED_128_Instance_MCS_Instance_1_n36 ;
    wire LED_128_Instance_MCS_Instance_1_n35 ;
    wire LED_128_Instance_MCS_Instance_1_n34 ;
    wire LED_128_Instance_MCS_Instance_1_n33 ;
    wire LED_128_Instance_MCS_Instance_1_n32 ;
    wire LED_128_Instance_MCS_Instance_1_n31 ;
    wire LED_128_Instance_MCS_Instance_1_n30 ;
    wire LED_128_Instance_MCS_Instance_1_n29 ;
    wire LED_128_Instance_MCS_Instance_1_n28 ;
    wire LED_128_Instance_MCS_Instance_1_n27 ;
    wire LED_128_Instance_MCS_Instance_1_n26 ;
    wire LED_128_Instance_MCS_Instance_1_n25 ;
    wire LED_128_Instance_MCS_Instance_1_n24 ;
    wire LED_128_Instance_MCS_Instance_1_n23 ;
    wire LED_128_Instance_MCS_Instance_1_n22 ;
    wire LED_128_Instance_MCS_Instance_1_n21 ;
    wire LED_128_Instance_MCS_Instance_1_n20 ;
    wire LED_128_Instance_MCS_Instance_1_n19 ;
    wire LED_128_Instance_MCS_Instance_1_n18 ;
    wire LED_128_Instance_MCS_Instance_1_n17 ;
    wire LED_128_Instance_MCS_Instance_1_n16 ;
    wire LED_128_Instance_MCS_Instance_1_n15 ;
    wire LED_128_Instance_MCS_Instance_1_n14 ;
    wire LED_128_Instance_MCS_Instance_1_n13 ;
    wire LED_128_Instance_MCS_Instance_1_n12 ;
    wire LED_128_Instance_MCS_Instance_1_n11 ;
    wire LED_128_Instance_MCS_Instance_1_n10 ;
    wire LED_128_Instance_MCS_Instance_1_n9 ;
    wire LED_128_Instance_MCS_Instance_1_n8 ;
    wire LED_128_Instance_MCS_Instance_1_n7 ;
    wire LED_128_Instance_MCS_Instance_1_n6 ;
    wire LED_128_Instance_MCS_Instance_1_n5 ;
    wire LED_128_Instance_MCS_Instance_1_n4 ;
    wire LED_128_Instance_MCS_Instance_1_n3 ;
    wire LED_128_Instance_MCS_Instance_1_n2 ;
    wire LED_128_Instance_MCS_Instance_1_n1 ;
    wire LED_128_Instance_MCS_Instance_2_n38 ;
    wire LED_128_Instance_MCS_Instance_2_n37 ;
    wire LED_128_Instance_MCS_Instance_2_n36 ;
    wire LED_128_Instance_MCS_Instance_2_n35 ;
    wire LED_128_Instance_MCS_Instance_2_n34 ;
    wire LED_128_Instance_MCS_Instance_2_n33 ;
    wire LED_128_Instance_MCS_Instance_2_n32 ;
    wire LED_128_Instance_MCS_Instance_2_n31 ;
    wire LED_128_Instance_MCS_Instance_2_n30 ;
    wire LED_128_Instance_MCS_Instance_2_n29 ;
    wire LED_128_Instance_MCS_Instance_2_n28 ;
    wire LED_128_Instance_MCS_Instance_2_n27 ;
    wire LED_128_Instance_MCS_Instance_2_n26 ;
    wire LED_128_Instance_MCS_Instance_2_n25 ;
    wire LED_128_Instance_MCS_Instance_2_n24 ;
    wire LED_128_Instance_MCS_Instance_2_n23 ;
    wire LED_128_Instance_MCS_Instance_2_n22 ;
    wire LED_128_Instance_MCS_Instance_2_n21 ;
    wire LED_128_Instance_MCS_Instance_2_n20 ;
    wire LED_128_Instance_MCS_Instance_2_n19 ;
    wire LED_128_Instance_MCS_Instance_2_n18 ;
    wire LED_128_Instance_MCS_Instance_2_n17 ;
    wire LED_128_Instance_MCS_Instance_2_n16 ;
    wire LED_128_Instance_MCS_Instance_2_n15 ;
    wire LED_128_Instance_MCS_Instance_2_n14 ;
    wire LED_128_Instance_MCS_Instance_2_n13 ;
    wire LED_128_Instance_MCS_Instance_2_n12 ;
    wire LED_128_Instance_MCS_Instance_2_n11 ;
    wire LED_128_Instance_MCS_Instance_2_n10 ;
    wire LED_128_Instance_MCS_Instance_2_n9 ;
    wire LED_128_Instance_MCS_Instance_2_n8 ;
    wire LED_128_Instance_MCS_Instance_2_n7 ;
    wire LED_128_Instance_MCS_Instance_2_n6 ;
    wire LED_128_Instance_MCS_Instance_2_n5 ;
    wire LED_128_Instance_MCS_Instance_2_n4 ;
    wire LED_128_Instance_MCS_Instance_2_n3 ;
    wire LED_128_Instance_MCS_Instance_2_n2 ;
    wire LED_128_Instance_MCS_Instance_2_n1 ;
    wire LED_128_Instance_MCS_Instance_3_n38 ;
    wire LED_128_Instance_MCS_Instance_3_n37 ;
    wire LED_128_Instance_MCS_Instance_3_n36 ;
    wire LED_128_Instance_MCS_Instance_3_n35 ;
    wire LED_128_Instance_MCS_Instance_3_n34 ;
    wire LED_128_Instance_MCS_Instance_3_n33 ;
    wire LED_128_Instance_MCS_Instance_3_n32 ;
    wire LED_128_Instance_MCS_Instance_3_n31 ;
    wire LED_128_Instance_MCS_Instance_3_n30 ;
    wire LED_128_Instance_MCS_Instance_3_n29 ;
    wire LED_128_Instance_MCS_Instance_3_n28 ;
    wire LED_128_Instance_MCS_Instance_3_n27 ;
    wire LED_128_Instance_MCS_Instance_3_n26 ;
    wire LED_128_Instance_MCS_Instance_3_n25 ;
    wire LED_128_Instance_MCS_Instance_3_n24 ;
    wire LED_128_Instance_MCS_Instance_3_n23 ;
    wire LED_128_Instance_MCS_Instance_3_n22 ;
    wire LED_128_Instance_MCS_Instance_3_n21 ;
    wire LED_128_Instance_MCS_Instance_3_n20 ;
    wire LED_128_Instance_MCS_Instance_3_n19 ;
    wire LED_128_Instance_MCS_Instance_3_n18 ;
    wire LED_128_Instance_MCS_Instance_3_n17 ;
    wire LED_128_Instance_MCS_Instance_3_n16 ;
    wire LED_128_Instance_MCS_Instance_3_n15 ;
    wire LED_128_Instance_MCS_Instance_3_n14 ;
    wire LED_128_Instance_MCS_Instance_3_n13 ;
    wire LED_128_Instance_MCS_Instance_3_n12 ;
    wire LED_128_Instance_MCS_Instance_3_n11 ;
    wire LED_128_Instance_MCS_Instance_3_n10 ;
    wire LED_128_Instance_MCS_Instance_3_n9 ;
    wire LED_128_Instance_MCS_Instance_3_n8 ;
    wire LED_128_Instance_MCS_Instance_3_n7 ;
    wire LED_128_Instance_MCS_Instance_3_n6 ;
    wire LED_128_Instance_MCS_Instance_3_n5 ;
    wire LED_128_Instance_MCS_Instance_3_n4 ;
    wire LED_128_Instance_MCS_Instance_3_n3 ;
    wire LED_128_Instance_MCS_Instance_3_n2 ;
    wire LED_128_Instance_MCS_Instance_3_n1 ;
    wire LED_128_Instance_ks_reg_0__Q ;
    wire [5:0] roundconstant ;
    wire [63:0] LED_128_Instance_subcells_out ;
    wire [63:0] LED_128_Instance_addconst_out ;
    wire [63:0] LED_128_Instance_addroundkey_tmp ;
    wire [63:0] LED_128_Instance_current_roundkey ;
    wire [63:0] LED_128_Instance_state1 ;
    wire [63:0] LED_128_Instance_state0 ;
    wire [63:0] LED_128_Instance_mixcolumns_out ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;

    /* cells in depth 0 */
    NOR2_X1 U16 ( .A1 (roundconstant[4]), .A2 (roundconstant[1]), .ZN (n14) ) ;
    NAND2_X1 U17 ( .A1 (roundconstant[0]), .A2 (n14), .ZN (n16) ) ;
    NOR2_X1 U18 ( .A1 (roundconstant[5]), .A2 (n16), .ZN (n17) ) ;
    NAND2_X1 U19 ( .A1 (roundconstant[3]), .A2 (n17), .ZN (n18) ) ;
    NOR2_X1 U20 ( .A1 (roundconstant[2]), .A2 (n18), .ZN (n19) ) ;
    NOR2_X1 U21 ( .A1 (OUT_done), .A2 (n19), .ZN (n20) ) ;
    NOR2_X1 U22 ( .A1 (IN_reset), .A2 (n20), .ZN (n15) ) ;
    NAND2_X1 LED_128_Instance_U30 ( .A1 (LED_128_Instance_n33), .A2 (LED_128_Instance_n32), .ZN (LED_128_Instance_n34) ) ;
    XNOR2_X1 LED_128_Instance_U29 ( .A (LED_128_Instance_n25), .B (LED_128_Instance_n23), .ZN (LED_128_Instance_n32) ) ;
    XOR2_X1 LED_128_Instance_U28 ( .A (LED_128_Instance_n4), .B (LED_128_Instance_n26), .Z (LED_128_Instance_n23) ) ;
    NAND2_X1 LED_128_Instance_U27 ( .A1 (LED_128_Instance_n21), .A2 (LED_128_Instance_n20), .ZN (LED_128_Instance_n33) ) ;
    NAND2_X1 LED_128_Instance_U26 ( .A1 (LED_128_Instance_n19), .A2 (LED_128_Instance_n18), .ZN (LED_128_Instance_n20) ) ;
    NOR2_X1 LED_128_Instance_U25 ( .A1 (LED_128_Instance_n24), .A2 (LED_128_Instance_n1), .ZN (LED_128_Instance_n18) ) ;
    NOR2_X1 LED_128_Instance_U24 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n19) ) ;
    NAND2_X1 LED_128_Instance_U23 ( .A1 (LED_128_Instance_n1), .A2 (LED_128_Instance_n17), .ZN (LED_128_Instance_n21) ) ;
    AND2_X1 LED_128_Instance_U22 ( .A1 (LED_128_Instance_n8), .A2 (LED_128_Instance_n4), .ZN (LED_128_Instance_n17) ) ;
    NAND2_X1 LED_128_Instance_U21 ( .A1 (LED_128_Instance_n29), .A2 (LED_128_Instance_n14), .ZN (LED_128_Instance_n15) ) ;
    NOR2_X1 LED_128_Instance_U20 ( .A1 (LED_128_Instance_n6), .A2 (LED_128_Instance_n13), .ZN (LED_128_Instance_n14) ) ;
    NAND2_X1 LED_128_Instance_U19 ( .A1 (LED_128_Instance_n5), .A2 (roundconstant[3]), .ZN (LED_128_Instance_n13) ) ;
    NAND2_X1 LED_128_Instance_U18 ( .A1 (LED_128_Instance_n28), .A2 (LED_128_Instance_n27), .ZN (LED_128_Instance_n16) ) ;
    NOR2_X1 LED_128_Instance_U17 ( .A1 (LED_128_Instance_n28), .A2 (IN_reset), .ZN (LED_128_Instance_N9) ) ;
    NOR2_X1 LED_128_Instance_U16 ( .A1 (IN_reset), .A2 (LED_128_Instance_n30), .ZN (LED_128_Instance_N8) ) ;
    NOR2_X1 LED_128_Instance_U15 ( .A1 (IN_reset), .A2 (LED_128_Instance_n5), .ZN (LED_128_Instance_N7) ) ;
    NOR2_X1 LED_128_Instance_U14 ( .A1 (IN_reset), .A2 (LED_128_Instance_n29), .ZN (LED_128_Instance_N6) ) ;
    NOR2_X1 LED_128_Instance_U13 ( .A1 (IN_reset), .A2 (LED_128_Instance_n6), .ZN (LED_128_Instance_N5) ) ;
    NOR2_X1 LED_128_Instance_U12 ( .A1 (LED_128_Instance_n1), .A2 (IN_reset), .ZN (LED_128_Instance_N13) ) ;
    NOR2_X1 LED_128_Instance_U11 ( .A1 (LED_128_Instance_n8), .A2 (IN_reset), .ZN (LED_128_Instance_N12) ) ;
    NOR2_X1 LED_128_Instance_U10 ( .A1 (LED_128_Instance_n4), .A2 (IN_reset), .ZN (LED_128_Instance_N11) ) ;
    NOR2_X1 LED_128_Instance_U9 ( .A1 (LED_128_Instance_n2), .A2 (IN_reset), .ZN (LED_128_Instance_N10) ) ;
    OR2_X1 LED_128_Instance_U8 ( .A1 (LED_128_Instance_n2), .A2 (LED_128_Instance_n21), .ZN (LED_128_Instance_n11) ) ;
    NAND2_X1 LED_128_Instance_U7 ( .A1 (LED_128_Instance_n34), .A2 (LED_128_Instance_n11), .ZN (LED_128_Instance_n31) ) ;
    NOR2_X1 LED_128_Instance_U6 ( .A1 (LED_128_Instance_n16), .A2 (LED_128_Instance_n15), .ZN (LED_128_Instance_n22) ) ;
    INV_X1 LED_128_Instance_U5 ( .A (LED_128_Instance_n11), .ZN (LED_128_Instance_n12) ) ;
    OR2_X1 LED_128_Instance_U4 ( .A1 (IN_reset), .A2 (LED_128_Instance_n10), .ZN (LED_128_Instance_N4) ) ;
    XNOR2_X1 LED_128_Instance_U3 ( .A (LED_128_Instance_n28), .B (LED_128_Instance_n27), .ZN (LED_128_Instance_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U4 ( .A (LED_128_Instance_n22), .ZN (LED_128_Instance_MUX_state0_n11) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U3 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n8) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U2 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n10) ) ;
    INV_X1 LED_128_Instance_MUX_state0_U1 ( .A (LED_128_Instance_MUX_state0_n11), .ZN (LED_128_Instance_MUX_state0_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U4 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n9) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U3 ( .A (LED_128_Instance_n12), .ZN (LED_128_Instance_MUX_current_roundkey_n10) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U2 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n7) ) ;
    INV_X1 LED_128_Instance_MUX_current_roundkey_U1 ( .A (LED_128_Instance_MUX_current_roundkey_n10), .ZN (LED_128_Instance_MUX_current_roundkey_n8) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_0_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({new_AGEMA_signal_1330, LED_128_Instance_current_roundkey[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_1_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({new_AGEMA_signal_1395, LED_128_Instance_current_roundkey[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_2_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_3_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({new_AGEMA_signal_1333, LED_128_Instance_current_roundkey[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({new_AGEMA_signal_1401, LED_128_Instance_current_roundkey[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({new_AGEMA_signal_1407, LED_128_Instance_current_roundkey[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({new_AGEMA_signal_1410, LED_128_Instance_current_roundkey[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({new_AGEMA_signal_1413, LED_128_Instance_current_roundkey[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({new_AGEMA_signal_1416, LED_128_Instance_current_roundkey[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({new_AGEMA_signal_1419, LED_128_Instance_current_roundkey[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({new_AGEMA_signal_1422, LED_128_Instance_current_roundkey[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({new_AGEMA_signal_1425, LED_128_Instance_current_roundkey[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({new_AGEMA_signal_1428, LED_128_Instance_current_roundkey[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({new_AGEMA_signal_1431, LED_128_Instance_current_roundkey[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({new_AGEMA_signal_1434, LED_128_Instance_current_roundkey[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_16_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({new_AGEMA_signal_1336, LED_128_Instance_current_roundkey[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_17_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({new_AGEMA_signal_1437, LED_128_Instance_current_roundkey[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_18_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({new_AGEMA_signal_1440, LED_128_Instance_current_roundkey[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_19_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({new_AGEMA_signal_1339, LED_128_Instance_current_roundkey[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n9), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({new_AGEMA_signal_1443, LED_128_Instance_current_roundkey[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_21_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({new_AGEMA_signal_1446, LED_128_Instance_current_roundkey[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_22_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({new_AGEMA_signal_1342, LED_128_Instance_current_roundkey[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_23_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({new_AGEMA_signal_1449, LED_128_Instance_current_roundkey[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_24_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({new_AGEMA_signal_1345, LED_128_Instance_current_roundkey[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_25_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({new_AGEMA_signal_1452, LED_128_Instance_current_roundkey[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_26_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({new_AGEMA_signal_1348, LED_128_Instance_current_roundkey[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_27_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({new_AGEMA_signal_1455, LED_128_Instance_current_roundkey[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_28_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({new_AGEMA_signal_1351, LED_128_Instance_current_roundkey[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({new_AGEMA_signal_1458, LED_128_Instance_current_roundkey[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({new_AGEMA_signal_1461, LED_128_Instance_current_roundkey[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({new_AGEMA_signal_1464, LED_128_Instance_current_roundkey[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_32_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({new_AGEMA_signal_1354, LED_128_Instance_current_roundkey[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({new_AGEMA_signal_1467, LED_128_Instance_current_roundkey[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_34_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({new_AGEMA_signal_1357, LED_128_Instance_current_roundkey[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_35_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({new_AGEMA_signal_1360, LED_128_Instance_current_roundkey[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_36_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({new_AGEMA_signal_1363, LED_128_Instance_current_roundkey[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_37_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({new_AGEMA_signal_1470, LED_128_Instance_current_roundkey[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({new_AGEMA_signal_1473, LED_128_Instance_current_roundkey[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_39_U1 ( .s (LED_128_Instance_n12), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({new_AGEMA_signal_1366, LED_128_Instance_current_roundkey[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({new_AGEMA_signal_1476, LED_128_Instance_current_roundkey[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({new_AGEMA_signal_1479, LED_128_Instance_current_roundkey[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({new_AGEMA_signal_1482, LED_128_Instance_current_roundkey[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_43_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({new_AGEMA_signal_1485, LED_128_Instance_current_roundkey[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({new_AGEMA_signal_1488, LED_128_Instance_current_roundkey[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({new_AGEMA_signal_1491, LED_128_Instance_current_roundkey[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({new_AGEMA_signal_1494, LED_128_Instance_current_roundkey[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_47_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({new_AGEMA_signal_1497, LED_128_Instance_current_roundkey[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_48_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({new_AGEMA_signal_1500, LED_128_Instance_current_roundkey[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_49_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({new_AGEMA_signal_1503, LED_128_Instance_current_roundkey[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_50_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({new_AGEMA_signal_1506, LED_128_Instance_current_roundkey[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_51_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n8), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({new_AGEMA_signal_1509, LED_128_Instance_current_roundkey[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_52_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({new_AGEMA_signal_1512, LED_128_Instance_current_roundkey[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_53_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({new_AGEMA_signal_1515, LED_128_Instance_current_roundkey[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({new_AGEMA_signal_1518, LED_128_Instance_current_roundkey[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({new_AGEMA_signal_1521, LED_128_Instance_current_roundkey[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({new_AGEMA_signal_1524, LED_128_Instance_current_roundkey[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({new_AGEMA_signal_1527, LED_128_Instance_current_roundkey[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({new_AGEMA_signal_1530, LED_128_Instance_current_roundkey[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({new_AGEMA_signal_1533, LED_128_Instance_current_roundkey[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({new_AGEMA_signal_1536, LED_128_Instance_current_roundkey[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({new_AGEMA_signal_1539, LED_128_Instance_current_roundkey[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({new_AGEMA_signal_1542, LED_128_Instance_current_roundkey[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_current_roundkey_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_current_roundkey_n7), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({new_AGEMA_signal_1545, LED_128_Instance_current_roundkey[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U64 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({new_AGEMA_signal_1416, LED_128_Instance_current_roundkey[9]}), .c ({new_AGEMA_signal_1554, LED_128_Instance_addroundkey_tmp[9]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U63 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({new_AGEMA_signal_1413, LED_128_Instance_current_roundkey[8]}), .c ({new_AGEMA_signal_1556, LED_128_Instance_addroundkey_tmp[8]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U62 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({new_AGEMA_signal_1410, LED_128_Instance_current_roundkey[7]}), .c ({new_AGEMA_signal_1558, LED_128_Instance_addroundkey_tmp[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U61 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({new_AGEMA_signal_1407, LED_128_Instance_current_roundkey[6]}), .c ({new_AGEMA_signal_1560, LED_128_Instance_addroundkey_tmp[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U60 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({new_AGEMA_signal_1545, LED_128_Instance_current_roundkey[63]}), .c ({new_AGEMA_signal_1562, LED_128_Instance_addroundkey_tmp[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U59 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({new_AGEMA_signal_1542, LED_128_Instance_current_roundkey[62]}), .c ({new_AGEMA_signal_1564, LED_128_Instance_addroundkey_tmp[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U58 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({new_AGEMA_signal_1539, LED_128_Instance_current_roundkey[61]}), .c ({new_AGEMA_signal_1566, LED_128_Instance_addroundkey_tmp[61]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U57 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({new_AGEMA_signal_1536, LED_128_Instance_current_roundkey[60]}), .c ({new_AGEMA_signal_1568, LED_128_Instance_addroundkey_tmp[60]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U56 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({new_AGEMA_signal_1404, LED_128_Instance_current_roundkey[5]}), .c ({new_AGEMA_signal_1570, LED_128_Instance_addroundkey_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U55 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({new_AGEMA_signal_1533, LED_128_Instance_current_roundkey[59]}), .c ({new_AGEMA_signal_1572, LED_128_Instance_addroundkey_tmp[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U54 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({new_AGEMA_signal_1530, LED_128_Instance_current_roundkey[58]}), .c ({new_AGEMA_signal_1574, LED_128_Instance_addroundkey_tmp[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U53 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({new_AGEMA_signal_1527, LED_128_Instance_current_roundkey[57]}), .c ({new_AGEMA_signal_1576, LED_128_Instance_addroundkey_tmp[57]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U52 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({new_AGEMA_signal_1524, LED_128_Instance_current_roundkey[56]}), .c ({new_AGEMA_signal_1578, LED_128_Instance_addroundkey_tmp[56]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U51 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({new_AGEMA_signal_1521, LED_128_Instance_current_roundkey[55]}), .c ({new_AGEMA_signal_1580, LED_128_Instance_addroundkey_tmp[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U50 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({new_AGEMA_signal_1518, LED_128_Instance_current_roundkey[54]}), .c ({new_AGEMA_signal_1582, LED_128_Instance_addroundkey_tmp[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U49 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({new_AGEMA_signal_1515, LED_128_Instance_current_roundkey[53]}), .c ({new_AGEMA_signal_1584, LED_128_Instance_addroundkey_tmp[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U48 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({new_AGEMA_signal_1512, LED_128_Instance_current_roundkey[52]}), .c ({new_AGEMA_signal_1586, LED_128_Instance_addroundkey_tmp[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U47 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({new_AGEMA_signal_1509, LED_128_Instance_current_roundkey[51]}), .c ({new_AGEMA_signal_1588, LED_128_Instance_addroundkey_tmp[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U46 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({new_AGEMA_signal_1506, LED_128_Instance_current_roundkey[50]}), .c ({new_AGEMA_signal_1590, LED_128_Instance_addroundkey_tmp[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U45 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({new_AGEMA_signal_1401, LED_128_Instance_current_roundkey[4]}), .c ({new_AGEMA_signal_1592, LED_128_Instance_addroundkey_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U44 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({new_AGEMA_signal_1503, LED_128_Instance_current_roundkey[49]}), .c ({new_AGEMA_signal_1594, LED_128_Instance_addroundkey_tmp[49]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U43 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({new_AGEMA_signal_1500, LED_128_Instance_current_roundkey[48]}), .c ({new_AGEMA_signal_1596, LED_128_Instance_addroundkey_tmp[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U42 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({new_AGEMA_signal_1497, LED_128_Instance_current_roundkey[47]}), .c ({new_AGEMA_signal_1598, LED_128_Instance_addroundkey_tmp[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U41 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({new_AGEMA_signal_1494, LED_128_Instance_current_roundkey[46]}), .c ({new_AGEMA_signal_1600, LED_128_Instance_addroundkey_tmp[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U40 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({new_AGEMA_signal_1491, LED_128_Instance_current_roundkey[45]}), .c ({new_AGEMA_signal_1602, LED_128_Instance_addroundkey_tmp[45]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U39 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({new_AGEMA_signal_1488, LED_128_Instance_current_roundkey[44]}), .c ({new_AGEMA_signal_1604, LED_128_Instance_addroundkey_tmp[44]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U38 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({new_AGEMA_signal_1485, LED_128_Instance_current_roundkey[43]}), .c ({new_AGEMA_signal_1606, LED_128_Instance_addroundkey_tmp[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U37 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({new_AGEMA_signal_1482, LED_128_Instance_current_roundkey[42]}), .c ({new_AGEMA_signal_1608, LED_128_Instance_addroundkey_tmp[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U36 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({new_AGEMA_signal_1479, LED_128_Instance_current_roundkey[41]}), .c ({new_AGEMA_signal_1610, LED_128_Instance_addroundkey_tmp[41]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U35 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({new_AGEMA_signal_1476, LED_128_Instance_current_roundkey[40]}), .c ({new_AGEMA_signal_1612, LED_128_Instance_addroundkey_tmp[40]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U34 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({new_AGEMA_signal_1333, LED_128_Instance_current_roundkey[3]}), .c ({new_AGEMA_signal_1368, LED_128_Instance_addroundkey_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U33 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({new_AGEMA_signal_1366, LED_128_Instance_current_roundkey[39]}), .c ({new_AGEMA_signal_1370, LED_128_Instance_addroundkey_tmp[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U32 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({new_AGEMA_signal_1473, LED_128_Instance_current_roundkey[38]}), .c ({new_AGEMA_signal_1614, LED_128_Instance_addroundkey_tmp[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U31 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({new_AGEMA_signal_1470, LED_128_Instance_current_roundkey[37]}), .c ({new_AGEMA_signal_1616, LED_128_Instance_addroundkey_tmp[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U30 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({new_AGEMA_signal_1363, LED_128_Instance_current_roundkey[36]}), .c ({new_AGEMA_signal_1372, LED_128_Instance_addroundkey_tmp[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U29 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({new_AGEMA_signal_1360, LED_128_Instance_current_roundkey[35]}), .c ({new_AGEMA_signal_1374, LED_128_Instance_addroundkey_tmp[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U28 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({new_AGEMA_signal_1357, LED_128_Instance_current_roundkey[34]}), .c ({new_AGEMA_signal_1376, LED_128_Instance_addroundkey_tmp[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U27 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({new_AGEMA_signal_1467, LED_128_Instance_current_roundkey[33]}), .c ({new_AGEMA_signal_1618, LED_128_Instance_addroundkey_tmp[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U26 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({new_AGEMA_signal_1354, LED_128_Instance_current_roundkey[32]}), .c ({new_AGEMA_signal_1378, LED_128_Instance_addroundkey_tmp[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U25 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({new_AGEMA_signal_1464, LED_128_Instance_current_roundkey[31]}), .c ({new_AGEMA_signal_1620, LED_128_Instance_addroundkey_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U24 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({new_AGEMA_signal_1461, LED_128_Instance_current_roundkey[30]}), .c ({new_AGEMA_signal_1622, LED_128_Instance_addroundkey_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U23 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({new_AGEMA_signal_1398, LED_128_Instance_current_roundkey[2]}), .c ({new_AGEMA_signal_1624, LED_128_Instance_addroundkey_tmp[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U22 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({new_AGEMA_signal_1458, LED_128_Instance_current_roundkey[29]}), .c ({new_AGEMA_signal_1626, LED_128_Instance_addroundkey_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U21 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({new_AGEMA_signal_1351, LED_128_Instance_current_roundkey[28]}), .c ({new_AGEMA_signal_1380, LED_128_Instance_addroundkey_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U20 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({new_AGEMA_signal_1455, LED_128_Instance_current_roundkey[27]}), .c ({new_AGEMA_signal_1628, LED_128_Instance_addroundkey_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U19 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({new_AGEMA_signal_1348, LED_128_Instance_current_roundkey[26]}), .c ({new_AGEMA_signal_1382, LED_128_Instance_addroundkey_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U18 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({new_AGEMA_signal_1452, LED_128_Instance_current_roundkey[25]}), .c ({new_AGEMA_signal_1630, LED_128_Instance_addroundkey_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U17 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({new_AGEMA_signal_1345, LED_128_Instance_current_roundkey[24]}), .c ({new_AGEMA_signal_1384, LED_128_Instance_addroundkey_tmp[24]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U16 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({new_AGEMA_signal_1449, LED_128_Instance_current_roundkey[23]}), .c ({new_AGEMA_signal_1632, LED_128_Instance_addroundkey_tmp[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U15 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({new_AGEMA_signal_1342, LED_128_Instance_current_roundkey[22]}), .c ({new_AGEMA_signal_1386, LED_128_Instance_addroundkey_tmp[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U14 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({new_AGEMA_signal_1446, LED_128_Instance_current_roundkey[21]}), .c ({new_AGEMA_signal_1634, LED_128_Instance_addroundkey_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U13 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({new_AGEMA_signal_1443, LED_128_Instance_current_roundkey[20]}), .c ({new_AGEMA_signal_1636, LED_128_Instance_addroundkey_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U12 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({new_AGEMA_signal_1395, LED_128_Instance_current_roundkey[1]}), .c ({new_AGEMA_signal_1638, LED_128_Instance_addroundkey_tmp[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U11 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({new_AGEMA_signal_1339, LED_128_Instance_current_roundkey[19]}), .c ({new_AGEMA_signal_1388, LED_128_Instance_addroundkey_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U10 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({new_AGEMA_signal_1440, LED_128_Instance_current_roundkey[18]}), .c ({new_AGEMA_signal_1640, LED_128_Instance_addroundkey_tmp[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U9 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({new_AGEMA_signal_1437, LED_128_Instance_current_roundkey[17]}), .c ({new_AGEMA_signal_1642, LED_128_Instance_addroundkey_tmp[17]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U8 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({new_AGEMA_signal_1336, LED_128_Instance_current_roundkey[16]}), .c ({new_AGEMA_signal_1390, LED_128_Instance_addroundkey_tmp[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U7 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({new_AGEMA_signal_1434, LED_128_Instance_current_roundkey[15]}), .c ({new_AGEMA_signal_1644, LED_128_Instance_addroundkey_tmp[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U6 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({new_AGEMA_signal_1431, LED_128_Instance_current_roundkey[14]}), .c ({new_AGEMA_signal_1646, LED_128_Instance_addroundkey_tmp[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U5 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({new_AGEMA_signal_1428, LED_128_Instance_current_roundkey[13]}), .c ({new_AGEMA_signal_1648, LED_128_Instance_addroundkey_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U4 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({new_AGEMA_signal_1425, LED_128_Instance_current_roundkey[12]}), .c ({new_AGEMA_signal_1650, LED_128_Instance_addroundkey_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U3 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({new_AGEMA_signal_1422, LED_128_Instance_current_roundkey[11]}), .c ({new_AGEMA_signal_1652, LED_128_Instance_addroundkey_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U2 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({new_AGEMA_signal_1419, LED_128_Instance_current_roundkey[10]}), .c ({new_AGEMA_signal_1654, LED_128_Instance_addroundkey_tmp[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_addRoundKey_instance_U1 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({new_AGEMA_signal_1330, LED_128_Instance_current_roundkey[0]}), .c ({new_AGEMA_signal_1392, LED_128_Instance_addroundkey_tmp[0]}) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U3 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n7) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U2 ( .A (LED_128_Instance_n31), .ZN (LED_128_Instance_MUX_addroundkey_out_n9) ) ;
    INV_X1 LED_128_Instance_MUX_addroundkey_out_U1 ( .A (LED_128_Instance_MUX_addroundkey_out_n9), .ZN (LED_128_Instance_MUX_addroundkey_out_n8) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_0_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({new_AGEMA_signal_1392, LED_128_Instance_addroundkey_tmp[0]}), .c ({new_AGEMA_signal_1546, LED_128_Instance_addroundkey_out_0_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_1_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({new_AGEMA_signal_1638, LED_128_Instance_addroundkey_tmp[1]}), .c ({new_AGEMA_signal_1666, LED_128_Instance_addroundkey_out_1_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_2_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({new_AGEMA_signal_1624, LED_128_Instance_addroundkey_tmp[2]}), .c ({new_AGEMA_signal_1667, LED_128_Instance_addroundkey_out_2_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_3_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({new_AGEMA_signal_1368, LED_128_Instance_addroundkey_tmp[3]}), .c ({new_AGEMA_signal_1547, LED_128_Instance_addroundkey_out_3_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_4_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({new_AGEMA_signal_1592, LED_128_Instance_addroundkey_tmp[4]}), .c ({new_AGEMA_signal_1668, LED_128_Instance_addroundkey_out_4_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_5_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({new_AGEMA_signal_1570, LED_128_Instance_addroundkey_tmp[5]}), .c ({new_AGEMA_signal_1669, LED_128_Instance_addroundkey_out_5_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_6_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({new_AGEMA_signal_1560, LED_128_Instance_addroundkey_tmp[6]}), .c ({new_AGEMA_signal_1670, LED_128_Instance_addroundkey_out_6_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_7_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({new_AGEMA_signal_1558, LED_128_Instance_addroundkey_tmp[7]}), .c ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_8_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({new_AGEMA_signal_1556, LED_128_Instance_addroundkey_tmp[8]}), .c ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_9_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({new_AGEMA_signal_1554, LED_128_Instance_addroundkey_tmp[9]}), .c ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_10_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({new_AGEMA_signal_1654, LED_128_Instance_addroundkey_tmp[10]}), .c ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_11_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({new_AGEMA_signal_1652, LED_128_Instance_addroundkey_tmp[11]}), .c ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_12_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({new_AGEMA_signal_1650, LED_128_Instance_addroundkey_tmp[12]}), .c ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_13_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({new_AGEMA_signal_1648, LED_128_Instance_addroundkey_tmp[13]}), .c ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_14_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({new_AGEMA_signal_1646, LED_128_Instance_addroundkey_tmp[14]}), .c ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_15_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({new_AGEMA_signal_1644, LED_128_Instance_addroundkey_tmp[15]}), .c ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_16_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({new_AGEMA_signal_1390, LED_128_Instance_addroundkey_tmp[16]}), .c ({new_AGEMA_signal_1548, LED_128_Instance_addroundkey_out_16_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_17_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({new_AGEMA_signal_1642, LED_128_Instance_addroundkey_tmp[17]}), .c ({new_AGEMA_signal_1680, LED_128_Instance_addroundkey_out_17_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_18_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({new_AGEMA_signal_1640, LED_128_Instance_addroundkey_tmp[18]}), .c ({new_AGEMA_signal_1681, LED_128_Instance_addroundkey_out_18_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_19_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({new_AGEMA_signal_1388, LED_128_Instance_addroundkey_tmp[19]}), .c ({new_AGEMA_signal_1549, LED_128_Instance_addroundkey_out_19_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_20_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n8), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({new_AGEMA_signal_1636, LED_128_Instance_addroundkey_tmp[20]}), .c ({new_AGEMA_signal_1682, LED_128_Instance_addroundkey_out_20_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_21_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({new_AGEMA_signal_1634, LED_128_Instance_addroundkey_tmp[21]}), .c ({new_AGEMA_signal_1683, LED_128_Instance_addroundkey_out_21_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_22_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({new_AGEMA_signal_1386, LED_128_Instance_addroundkey_tmp[22]}), .c ({new_AGEMA_signal_1550, LED_128_Instance_addroundkey_out_22_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_23_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({new_AGEMA_signal_1632, LED_128_Instance_addroundkey_tmp[23]}), .c ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_24_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({new_AGEMA_signal_1384, LED_128_Instance_addroundkey_tmp[24]}), .c ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_25_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({new_AGEMA_signal_1630, LED_128_Instance_addroundkey_tmp[25]}), .c ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_26_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({new_AGEMA_signal_1382, LED_128_Instance_addroundkey_tmp[26]}), .c ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_27_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({new_AGEMA_signal_1628, LED_128_Instance_addroundkey_tmp[27]}), .c ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_28_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({new_AGEMA_signal_1380, LED_128_Instance_addroundkey_tmp[28]}), .c ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_29_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({new_AGEMA_signal_1626, LED_128_Instance_addroundkey_tmp[29]}), .c ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_30_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({new_AGEMA_signal_1622, LED_128_Instance_addroundkey_tmp[30]}), .c ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_31_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({new_AGEMA_signal_1620, LED_128_Instance_addroundkey_tmp[31]}), .c ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_32_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({new_AGEMA_signal_1378, LED_128_Instance_addroundkey_tmp[32]}), .c ({new_AGEMA_signal_1656, LED_128_Instance_addroundkey_out_32_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_33_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({new_AGEMA_signal_1618, LED_128_Instance_addroundkey_tmp[33]}), .c ({new_AGEMA_signal_1690, LED_128_Instance_addroundkey_out_33_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_34_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({new_AGEMA_signal_1376, LED_128_Instance_addroundkey_tmp[34]}), .c ({new_AGEMA_signal_1657, LED_128_Instance_addroundkey_out_34_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_35_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({new_AGEMA_signal_1374, LED_128_Instance_addroundkey_tmp[35]}), .c ({new_AGEMA_signal_1658, LED_128_Instance_addroundkey_out_35_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_36_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({new_AGEMA_signal_1372, LED_128_Instance_addroundkey_tmp[36]}), .c ({new_AGEMA_signal_1659, LED_128_Instance_addroundkey_out_36_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_37_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({new_AGEMA_signal_1616, LED_128_Instance_addroundkey_tmp[37]}), .c ({new_AGEMA_signal_1691, LED_128_Instance_addroundkey_out_37_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_38_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({new_AGEMA_signal_1614, LED_128_Instance_addroundkey_tmp[38]}), .c ({new_AGEMA_signal_1692, LED_128_Instance_addroundkey_out_38_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_39_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({new_AGEMA_signal_1370, LED_128_Instance_addroundkey_tmp[39]}), .c ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_40_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({new_AGEMA_signal_1612, LED_128_Instance_addroundkey_tmp[40]}), .c ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_41_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({new_AGEMA_signal_1610, LED_128_Instance_addroundkey_tmp[41]}), .c ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_42_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({new_AGEMA_signal_1608, LED_128_Instance_addroundkey_tmp[42]}), .c ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_43_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({new_AGEMA_signal_1606, LED_128_Instance_addroundkey_tmp[43]}), .c ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_44_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({new_AGEMA_signal_1604, LED_128_Instance_addroundkey_tmp[44]}), .c ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_45_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({new_AGEMA_signal_1602, LED_128_Instance_addroundkey_tmp[45]}), .c ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_46_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({new_AGEMA_signal_1600, LED_128_Instance_addroundkey_tmp[46]}), .c ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_47_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({new_AGEMA_signal_1598, LED_128_Instance_addroundkey_tmp[47]}), .c ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_48_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({new_AGEMA_signal_1596, LED_128_Instance_addroundkey_tmp[48]}), .c ({new_AGEMA_signal_1701, LED_128_Instance_addroundkey_out_48_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_49_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({new_AGEMA_signal_1594, LED_128_Instance_addroundkey_tmp[49]}), .c ({new_AGEMA_signal_1702, LED_128_Instance_addroundkey_out_49_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_50_U1 ( .s (LED_128_Instance_n31), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({new_AGEMA_signal_1590, LED_128_Instance_addroundkey_tmp[50]}), .c ({new_AGEMA_signal_1703, LED_128_Instance_addroundkey_out_50_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_51_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({new_AGEMA_signal_1588, LED_128_Instance_addroundkey_tmp[51]}), .c ({new_AGEMA_signal_1704, LED_128_Instance_addroundkey_out_51_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_52_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({new_AGEMA_signal_1586, LED_128_Instance_addroundkey_tmp[52]}), .c ({new_AGEMA_signal_1705, LED_128_Instance_addroundkey_out_52_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_53_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({new_AGEMA_signal_1584, LED_128_Instance_addroundkey_tmp[53]}), .c ({new_AGEMA_signal_1706, LED_128_Instance_addroundkey_out_53_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_54_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({new_AGEMA_signal_1582, LED_128_Instance_addroundkey_tmp[54]}), .c ({new_AGEMA_signal_1707, LED_128_Instance_addroundkey_out_54_}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_55_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({new_AGEMA_signal_1580, LED_128_Instance_addroundkey_tmp[55]}), .c ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_56_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({new_AGEMA_signal_1578, LED_128_Instance_addroundkey_tmp[56]}), .c ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_57_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({new_AGEMA_signal_1576, LED_128_Instance_addroundkey_tmp[57]}), .c ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_58_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({new_AGEMA_signal_1574, LED_128_Instance_addroundkey_tmp[58]}), .c ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_59_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({new_AGEMA_signal_1572, LED_128_Instance_addroundkey_tmp[59]}), .c ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_60_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({new_AGEMA_signal_1568, LED_128_Instance_addroundkey_tmp[60]}), .c ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_61_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({new_AGEMA_signal_1566, LED_128_Instance_addroundkey_tmp[61]}), .c ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_62_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({new_AGEMA_signal_1564, LED_128_Instance_addroundkey_tmp[62]}), .c ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_addroundkey_out_mux_inst_63_U1 ( .s (LED_128_Instance_MUX_addroundkey_out_n7), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({new_AGEMA_signal_1562, LED_128_Instance_addroundkey_tmp[63]}), .c ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U28 ( .a ({1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_1670, LED_128_Instance_addroundkey_out_6_}), .c ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U27 ( .a ({1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_1669, LED_128_Instance_addroundkey_out_5_}), .c ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U26 ( .a ({1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_1707, LED_128_Instance_addroundkey_out_54_}), .c ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U25 ( .a ({1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_1706, LED_128_Instance_addroundkey_out_53_}), .c ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U24 ( .a ({1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_1705, LED_128_Instance_addroundkey_out_52_}), .c ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U23 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1704, LED_128_Instance_addroundkey_out_51_}), .c ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U22 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1703, LED_128_Instance_addroundkey_out_50_}), .c ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U21 ( .a ({1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_1668, LED_128_Instance_addroundkey_out_4_}), .c ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U20 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1702, LED_128_Instance_addroundkey_out_49_}), .c ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U19 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1701, LED_128_Instance_addroundkey_out_48_}), .c ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U18 ( .a ({1'b0, 1'b1}), .b ({new_AGEMA_signal_1547, LED_128_Instance_addroundkey_out_3_}), .c ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U17 ( .a ({1'b0, roundconstant[5]}), .b ({new_AGEMA_signal_1692, LED_128_Instance_addroundkey_out_38_}), .c ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U16 ( .a ({1'b0, roundconstant[4]}), .b ({new_AGEMA_signal_1691, LED_128_Instance_addroundkey_out_37_}), .c ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U15 ( .a ({1'b0, roundconstant[3]}), .b ({new_AGEMA_signal_1659, LED_128_Instance_addroundkey_out_36_}), .c ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U14 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1658, LED_128_Instance_addroundkey_out_35_}), .c ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U13 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1657, LED_128_Instance_addroundkey_out_34_}), .c ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U12 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1690, LED_128_Instance_addroundkey_out_33_}), .c ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U11 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1656, LED_128_Instance_addroundkey_out_32_}), .c ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U10 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1667, LED_128_Instance_addroundkey_out_2_}), .c ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U9 ( .a ({1'b0, roundconstant[2]}), .b ({new_AGEMA_signal_1550, LED_128_Instance_addroundkey_out_22_}), .c ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U8 ( .a ({1'b0, roundconstant[1]}), .b ({new_AGEMA_signal_1683, LED_128_Instance_addroundkey_out_21_}), .c ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U7 ( .a ({1'b0, roundconstant[0]}), .b ({new_AGEMA_signal_1682, LED_128_Instance_addroundkey_out_20_}), .c ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U6 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1666, LED_128_Instance_addroundkey_out_1_}), .c ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U5 ( .a ({1'b0, 1'b1}), .b ({new_AGEMA_signal_1549, LED_128_Instance_addroundkey_out_19_}), .c ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U4 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1681, LED_128_Instance_addroundkey_out_18_}), .c ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U3 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1680, LED_128_Instance_addroundkey_out_17_}), .c ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U2 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1548, LED_128_Instance_addroundkey_out_16_}), .c ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_AddConstants_instance_U1 ( .a ({1'b0, 1'b0}), .b ({new_AGEMA_signal_1546, LED_128_Instance_addroundkey_out_0_}), .c ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_U3 ( .a ({new_AGEMA_signal_1800, LED_128_Instance_SBox_Instance_0_L0}), .b ({new_AGEMA_signal_1876, LED_128_Instance_SBox_Instance_0_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_U2 ( .a ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_1721, LED_128_Instance_SBox_Instance_0_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_U1 ( .a ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_1799, LED_128_Instance_SBox_Instance_0_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR1_U1 ( .a ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}), .b ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_1800, LED_128_Instance_SBox_Instance_0_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR2_U1 ( .a ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .b ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR3_U1 ( .a ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .c ({new_AGEMA_signal_1877, LED_128_Instance_SBox_Instance_0_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR4_U1 ( .a ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_1665, LED_128_Instance_addconst_out[0]}), .c ({new_AGEMA_signal_1722, LED_128_Instance_SBox_Instance_0_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR5_U1 ( .a ({new_AGEMA_signal_1722, LED_128_Instance_SBox_Instance_0_L3}), .b ({new_AGEMA_signal_1800, LED_128_Instance_SBox_Instance_0_L0}), .c ({new_AGEMA_signal_1878, LED_128_Instance_SBox_Instance_0_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR6_U1 ( .a ({new_AGEMA_signal_1661, LED_128_Instance_addconst_out[3]}), .b ({new_AGEMA_signal_1742, LED_128_Instance_addconst_out[1]}), .c ({new_AGEMA_signal_1802, LED_128_Instance_SBox_Instance_0_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR9_U1 ( .a ({new_AGEMA_signal_1801, LED_128_Instance_SBox_Instance_0_L1}), .b ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}), .c ({new_AGEMA_signal_1879, LED_128_Instance_SBox_Instance_0_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_U3 ( .a ({new_AGEMA_signal_1804, LED_128_Instance_SBox_Instance_1_L0}), .b ({new_AGEMA_signal_1881, LED_128_Instance_SBox_Instance_1_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_U2 ( .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_1745, LED_128_Instance_SBox_Instance_1_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_U1 ( .a ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_1803, LED_128_Instance_SBox_Instance_1_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR1_U1 ( .a ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}), .b ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_1804, LED_128_Instance_SBox_Instance_1_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR2_U1 ( .a ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .b ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR3_U1 ( .a ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .c ({new_AGEMA_signal_1882, LED_128_Instance_SBox_Instance_1_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR4_U1 ( .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_1733, LED_128_Instance_addconst_out[4]}), .c ({new_AGEMA_signal_1806, LED_128_Instance_SBox_Instance_1_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR5_U1 ( .a ({new_AGEMA_signal_1806, LED_128_Instance_SBox_Instance_1_L3}), .b ({new_AGEMA_signal_1804, LED_128_Instance_SBox_Instance_1_L0}), .c ({new_AGEMA_signal_1883, LED_128_Instance_SBox_Instance_1_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR6_U1 ( .a ({new_AGEMA_signal_1671, LED_128_Instance_addconst_out[7]}), .b ({new_AGEMA_signal_1727, LED_128_Instance_addconst_out[5]}), .c ({new_AGEMA_signal_1807, LED_128_Instance_SBox_Instance_1_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR9_U1 ( .a ({new_AGEMA_signal_1805, LED_128_Instance_SBox_Instance_1_L1}), .b ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}), .c ({new_AGEMA_signal_1884, LED_128_Instance_SBox_Instance_1_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_U3 ( .a ({new_AGEMA_signal_1748, LED_128_Instance_SBox_Instance_2_L0}), .b ({new_AGEMA_signal_1808, LED_128_Instance_SBox_Instance_2_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_U2 ( .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_1746, LED_128_Instance_SBox_Instance_2_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_U1 ( .a ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_1747, LED_128_Instance_SBox_Instance_2_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR1_U1 ( .a ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .b ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_1748, LED_128_Instance_SBox_Instance_2_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR2_U1 ( .a ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .b ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR3_U1 ( .a ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .c ({new_AGEMA_signal_1809, LED_128_Instance_SBox_Instance_2_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR4_U1 ( .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_1672, LED_128_Instance_addconst_out[8]}), .c ({new_AGEMA_signal_1750, LED_128_Instance_SBox_Instance_2_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR5_U1 ( .a ({new_AGEMA_signal_1750, LED_128_Instance_SBox_Instance_2_L3}), .b ({new_AGEMA_signal_1748, LED_128_Instance_SBox_Instance_2_L0}), .c ({new_AGEMA_signal_1810, LED_128_Instance_SBox_Instance_2_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR6_U1 ( .a ({new_AGEMA_signal_1675, LED_128_Instance_addconst_out[11]}), .b ({new_AGEMA_signal_1673, LED_128_Instance_addconst_out[9]}), .c ({new_AGEMA_signal_1751, LED_128_Instance_SBox_Instance_2_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR9_U1 ( .a ({new_AGEMA_signal_1749, LED_128_Instance_SBox_Instance_2_L1}), .b ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .c ({new_AGEMA_signal_1811, LED_128_Instance_SBox_Instance_2_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_U3 ( .a ({new_AGEMA_signal_1754, LED_128_Instance_SBox_Instance_3_L0}), .b ({new_AGEMA_signal_1813, LED_128_Instance_SBox_Instance_3_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_U2 ( .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_1752, LED_128_Instance_SBox_Instance_3_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_U1 ( .a ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_1753, LED_128_Instance_SBox_Instance_3_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR1_U1 ( .a ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .b ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_1754, LED_128_Instance_SBox_Instance_3_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR2_U1 ( .a ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .b ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR3_U1 ( .a ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .c ({new_AGEMA_signal_1814, LED_128_Instance_SBox_Instance_3_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR4_U1 ( .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_1676, LED_128_Instance_addconst_out[12]}), .c ({new_AGEMA_signal_1756, LED_128_Instance_SBox_Instance_3_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR5_U1 ( .a ({new_AGEMA_signal_1756, LED_128_Instance_SBox_Instance_3_L3}), .b ({new_AGEMA_signal_1754, LED_128_Instance_SBox_Instance_3_L0}), .c ({new_AGEMA_signal_1815, LED_128_Instance_SBox_Instance_3_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR6_U1 ( .a ({new_AGEMA_signal_1679, LED_128_Instance_addconst_out[15]}), .b ({new_AGEMA_signal_1677, LED_128_Instance_addconst_out[13]}), .c ({new_AGEMA_signal_1757, LED_128_Instance_SBox_Instance_3_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR9_U1 ( .a ({new_AGEMA_signal_1755, LED_128_Instance_SBox_Instance_3_L1}), .b ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .c ({new_AGEMA_signal_1816, LED_128_Instance_SBox_Instance_3_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_U3 ( .a ({new_AGEMA_signal_1819, LED_128_Instance_SBox_Instance_4_L0}), .b ({new_AGEMA_signal_1890, LED_128_Instance_SBox_Instance_4_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_U2 ( .a ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_1723, LED_128_Instance_SBox_Instance_4_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_U1 ( .a ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_1818, LED_128_Instance_SBox_Instance_4_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR1_U1 ( .a ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}), .b ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_1819, LED_128_Instance_SBox_Instance_4_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR2_U1 ( .a ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .b ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR3_U1 ( .a ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .c ({new_AGEMA_signal_1891, LED_128_Instance_SBox_Instance_4_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR4_U1 ( .a ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_1664, LED_128_Instance_addconst_out[16]}), .c ({new_AGEMA_signal_1724, LED_128_Instance_SBox_Instance_4_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR5_U1 ( .a ({new_AGEMA_signal_1724, LED_128_Instance_SBox_Instance_4_L3}), .b ({new_AGEMA_signal_1819, LED_128_Instance_SBox_Instance_4_L0}), .c ({new_AGEMA_signal_1892, LED_128_Instance_SBox_Instance_4_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR6_U1 ( .a ({new_AGEMA_signal_1663, LED_128_Instance_addconst_out[19]}), .b ({new_AGEMA_signal_1744, LED_128_Instance_addconst_out[17]}), .c ({new_AGEMA_signal_1821, LED_128_Instance_SBox_Instance_4_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR9_U1 ( .a ({new_AGEMA_signal_1820, LED_128_Instance_SBox_Instance_4_L1}), .b ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}), .c ({new_AGEMA_signal_1893, LED_128_Instance_SBox_Instance_4_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_U3 ( .a ({new_AGEMA_signal_1823, LED_128_Instance_SBox_Instance_5_L0}), .b ({new_AGEMA_signal_1895, LED_128_Instance_SBox_Instance_5_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_U2 ( .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_1758, LED_128_Instance_SBox_Instance_5_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_U1 ( .a ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_1822, LED_128_Instance_SBox_Instance_5_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR1_U1 ( .a ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}), .b ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_1823, LED_128_Instance_SBox_Instance_5_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR2_U1 ( .a ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .b ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR3_U1 ( .a ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .c ({new_AGEMA_signal_1896, LED_128_Instance_SBox_Instance_5_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR4_U1 ( .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_1741, LED_128_Instance_addconst_out[20]}), .c ({new_AGEMA_signal_1825, LED_128_Instance_SBox_Instance_5_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR5_U1 ( .a ({new_AGEMA_signal_1825, LED_128_Instance_SBox_Instance_5_L3}), .b ({new_AGEMA_signal_1823, LED_128_Instance_SBox_Instance_5_L0}), .c ({new_AGEMA_signal_1897, LED_128_Instance_SBox_Instance_5_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR6_U1 ( .a ({new_AGEMA_signal_1684, LED_128_Instance_addconst_out[23]}), .b ({new_AGEMA_signal_1740, LED_128_Instance_addconst_out[21]}), .c ({new_AGEMA_signal_1826, LED_128_Instance_SBox_Instance_5_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR9_U1 ( .a ({new_AGEMA_signal_1824, LED_128_Instance_SBox_Instance_5_L1}), .b ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}), .c ({new_AGEMA_signal_1898, LED_128_Instance_SBox_Instance_5_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_U3 ( .a ({new_AGEMA_signal_1761, LED_128_Instance_SBox_Instance_6_L0}), .b ({new_AGEMA_signal_1827, LED_128_Instance_SBox_Instance_6_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_U2 ( .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1759, LED_128_Instance_SBox_Instance_6_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_U1 ( .a ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_1760, LED_128_Instance_SBox_Instance_6_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR1_U1 ( .a ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .b ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_1761, LED_128_Instance_SBox_Instance_6_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR2_U1 ( .a ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .b ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR3_U1 ( .a ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .c ({new_AGEMA_signal_1828, LED_128_Instance_SBox_Instance_6_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR4_U1 ( .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1551, LED_128_Instance_addconst_out[24]}), .c ({new_AGEMA_signal_1763, LED_128_Instance_SBox_Instance_6_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR5_U1 ( .a ({new_AGEMA_signal_1763, LED_128_Instance_SBox_Instance_6_L3}), .b ({new_AGEMA_signal_1761, LED_128_Instance_SBox_Instance_6_L0}), .c ({new_AGEMA_signal_1829, LED_128_Instance_SBox_Instance_6_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR6_U1 ( .a ({new_AGEMA_signal_1686, LED_128_Instance_addconst_out[27]}), .b ({new_AGEMA_signal_1685, LED_128_Instance_addconst_out[25]}), .c ({new_AGEMA_signal_1764, LED_128_Instance_SBox_Instance_6_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR9_U1 ( .a ({new_AGEMA_signal_1762, LED_128_Instance_SBox_Instance_6_L1}), .b ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .c ({new_AGEMA_signal_1830, LED_128_Instance_SBox_Instance_6_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_U3 ( .a ({new_AGEMA_signal_1767, LED_128_Instance_SBox_Instance_7_L0}), .b ({new_AGEMA_signal_1832, LED_128_Instance_SBox_Instance_7_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_U2 ( .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1765, LED_128_Instance_SBox_Instance_7_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_U1 ( .a ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_1766, LED_128_Instance_SBox_Instance_7_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR1_U1 ( .a ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .b ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_1767, LED_128_Instance_SBox_Instance_7_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR2_U1 ( .a ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .b ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR3_U1 ( .a ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .c ({new_AGEMA_signal_1833, LED_128_Instance_SBox_Instance_7_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR4_U1 ( .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1655, LED_128_Instance_addconst_out[28]}), .c ({new_AGEMA_signal_1769, LED_128_Instance_SBox_Instance_7_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR5_U1 ( .a ({new_AGEMA_signal_1769, LED_128_Instance_SBox_Instance_7_L3}), .b ({new_AGEMA_signal_1767, LED_128_Instance_SBox_Instance_7_L0}), .c ({new_AGEMA_signal_1834, LED_128_Instance_SBox_Instance_7_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR6_U1 ( .a ({new_AGEMA_signal_1689, LED_128_Instance_addconst_out[31]}), .b ({new_AGEMA_signal_1687, LED_128_Instance_addconst_out[29]}), .c ({new_AGEMA_signal_1770, LED_128_Instance_SBox_Instance_7_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR9_U1 ( .a ({new_AGEMA_signal_1768, LED_128_Instance_SBox_Instance_7_L1}), .b ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .c ({new_AGEMA_signal_1835, LED_128_Instance_SBox_Instance_7_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_U3 ( .a ({new_AGEMA_signal_1838, LED_128_Instance_SBox_Instance_8_L0}), .b ({new_AGEMA_signal_1904, LED_128_Instance_SBox_Instance_8_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_U2 ( .a ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_1771, LED_128_Instance_SBox_Instance_8_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_U1 ( .a ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_1837, LED_128_Instance_SBox_Instance_8_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR1_U1 ( .a ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}), .b ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_1838, LED_128_Instance_SBox_Instance_8_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR2_U1 ( .a ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .b ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR3_U1 ( .a ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .c ({new_AGEMA_signal_1905, LED_128_Instance_SBox_Instance_8_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR4_U1 ( .a ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_1720, LED_128_Instance_addconst_out[32]}), .c ({new_AGEMA_signal_1772, LED_128_Instance_SBox_Instance_8_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR5_U1 ( .a ({new_AGEMA_signal_1772, LED_128_Instance_SBox_Instance_8_L3}), .b ({new_AGEMA_signal_1838, LED_128_Instance_SBox_Instance_8_L0}), .c ({new_AGEMA_signal_1906, LED_128_Instance_SBox_Instance_8_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR6_U1 ( .a ({new_AGEMA_signal_1718, LED_128_Instance_addconst_out[35]}), .b ({new_AGEMA_signal_1738, LED_128_Instance_addconst_out[33]}), .c ({new_AGEMA_signal_1840, LED_128_Instance_SBox_Instance_8_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR9_U1 ( .a ({new_AGEMA_signal_1839, LED_128_Instance_SBox_Instance_8_L1}), .b ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}), .c ({new_AGEMA_signal_1907, LED_128_Instance_SBox_Instance_8_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_U3 ( .a ({new_AGEMA_signal_1842, LED_128_Instance_SBox_Instance_9_L0}), .b ({new_AGEMA_signal_1909, LED_128_Instance_SBox_Instance_9_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_U2 ( .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_1725, LED_128_Instance_SBox_Instance_9_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_U1 ( .a ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_1841, LED_128_Instance_SBox_Instance_9_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR1_U1 ( .a ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}), .b ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_1842, LED_128_Instance_SBox_Instance_9_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR2_U1 ( .a ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .b ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR3_U1 ( .a ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .c ({new_AGEMA_signal_1910, LED_128_Instance_SBox_Instance_9_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR4_U1 ( .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_1717, LED_128_Instance_addconst_out[36]}), .c ({new_AGEMA_signal_1773, LED_128_Instance_SBox_Instance_9_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR5_U1 ( .a ({new_AGEMA_signal_1773, LED_128_Instance_SBox_Instance_9_L3}), .b ({new_AGEMA_signal_1842, LED_128_Instance_SBox_Instance_9_L0}), .c ({new_AGEMA_signal_1911, LED_128_Instance_SBox_Instance_9_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR6_U1 ( .a ({new_AGEMA_signal_1660, LED_128_Instance_addconst_out[39]}), .b ({new_AGEMA_signal_1737, LED_128_Instance_addconst_out[37]}), .c ({new_AGEMA_signal_1844, LED_128_Instance_SBox_Instance_9_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR9_U1 ( .a ({new_AGEMA_signal_1843, LED_128_Instance_SBox_Instance_9_L1}), .b ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}), .c ({new_AGEMA_signal_1912, LED_128_Instance_SBox_Instance_9_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_U3 ( .a ({new_AGEMA_signal_1776, LED_128_Instance_SBox_Instance_10_L0}), .b ({new_AGEMA_signal_1845, LED_128_Instance_SBox_Instance_10_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_U2 ( .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_1774, LED_128_Instance_SBox_Instance_10_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_U1 ( .a ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_1775, LED_128_Instance_SBox_Instance_10_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR1_U1 ( .a ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .b ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_1776, LED_128_Instance_SBox_Instance_10_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR2_U1 ( .a ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .b ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR3_U1 ( .a ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .c ({new_AGEMA_signal_1846, LED_128_Instance_SBox_Instance_10_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR4_U1 ( .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_1693, LED_128_Instance_addconst_out[40]}), .c ({new_AGEMA_signal_1778, LED_128_Instance_SBox_Instance_10_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR5_U1 ( .a ({new_AGEMA_signal_1778, LED_128_Instance_SBox_Instance_10_L3}), .b ({new_AGEMA_signal_1776, LED_128_Instance_SBox_Instance_10_L0}), .c ({new_AGEMA_signal_1847, LED_128_Instance_SBox_Instance_10_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR6_U1 ( .a ({new_AGEMA_signal_1696, LED_128_Instance_addconst_out[43]}), .b ({new_AGEMA_signal_1694, LED_128_Instance_addconst_out[41]}), .c ({new_AGEMA_signal_1779, LED_128_Instance_SBox_Instance_10_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR9_U1 ( .a ({new_AGEMA_signal_1777, LED_128_Instance_SBox_Instance_10_L1}), .b ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .c ({new_AGEMA_signal_1848, LED_128_Instance_SBox_Instance_10_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_U3 ( .a ({new_AGEMA_signal_1782, LED_128_Instance_SBox_Instance_11_L0}), .b ({new_AGEMA_signal_1850, LED_128_Instance_SBox_Instance_11_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_U2 ( .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_1780, LED_128_Instance_SBox_Instance_11_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_U1 ( .a ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_1781, LED_128_Instance_SBox_Instance_11_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR1_U1 ( .a ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .b ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_1782, LED_128_Instance_SBox_Instance_11_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR2_U1 ( .a ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .b ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR3_U1 ( .a ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .c ({new_AGEMA_signal_1851, LED_128_Instance_SBox_Instance_11_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR4_U1 ( .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_1697, LED_128_Instance_addconst_out[44]}), .c ({new_AGEMA_signal_1784, LED_128_Instance_SBox_Instance_11_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR5_U1 ( .a ({new_AGEMA_signal_1784, LED_128_Instance_SBox_Instance_11_L3}), .b ({new_AGEMA_signal_1782, LED_128_Instance_SBox_Instance_11_L0}), .c ({new_AGEMA_signal_1852, LED_128_Instance_SBox_Instance_11_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR6_U1 ( .a ({new_AGEMA_signal_1700, LED_128_Instance_addconst_out[47]}), .b ({new_AGEMA_signal_1698, LED_128_Instance_addconst_out[45]}), .c ({new_AGEMA_signal_1785, LED_128_Instance_SBox_Instance_11_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR9_U1 ( .a ({new_AGEMA_signal_1783, LED_128_Instance_SBox_Instance_11_L1}), .b ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .c ({new_AGEMA_signal_1853, LED_128_Instance_SBox_Instance_11_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_U3 ( .a ({new_AGEMA_signal_1857, LED_128_Instance_SBox_Instance_12_L0}), .b ({new_AGEMA_signal_1918, LED_128_Instance_SBox_Instance_12_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_U2 ( .a ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_1855, LED_128_Instance_SBox_Instance_12_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_U1 ( .a ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_1856, LED_128_Instance_SBox_Instance_12_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR1_U1 ( .a ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}), .b ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_1857, LED_128_Instance_SBox_Instance_12_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR2_U1 ( .a ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .b ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR3_U1 ( .a ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .c ({new_AGEMA_signal_1919, LED_128_Instance_SBox_Instance_12_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR4_U1 ( .a ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_1735, LED_128_Instance_addconst_out[48]}), .c ({new_AGEMA_signal_1859, LED_128_Instance_SBox_Instance_12_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR5_U1 ( .a ({new_AGEMA_signal_1859, LED_128_Instance_SBox_Instance_12_L3}), .b ({new_AGEMA_signal_1857, LED_128_Instance_SBox_Instance_12_L0}), .c ({new_AGEMA_signal_1920, LED_128_Instance_SBox_Instance_12_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR6_U1 ( .a ({new_AGEMA_signal_1731, LED_128_Instance_addconst_out[51]}), .b ({new_AGEMA_signal_1734, LED_128_Instance_addconst_out[49]}), .c ({new_AGEMA_signal_1860, LED_128_Instance_SBox_Instance_12_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR9_U1 ( .a ({new_AGEMA_signal_1858, LED_128_Instance_SBox_Instance_12_L1}), .b ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}), .c ({new_AGEMA_signal_1921, LED_128_Instance_SBox_Instance_12_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_U3 ( .a ({new_AGEMA_signal_1862, LED_128_Instance_SBox_Instance_13_L0}), .b ({new_AGEMA_signal_1923, LED_128_Instance_SBox_Instance_13_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_U2 ( .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_1786, LED_128_Instance_SBox_Instance_13_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_U1 ( .a ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_1861, LED_128_Instance_SBox_Instance_13_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR1_U1 ( .a ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}), .b ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_1862, LED_128_Instance_SBox_Instance_13_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR2_U1 ( .a ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .b ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR3_U1 ( .a ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .c ({new_AGEMA_signal_1924, LED_128_Instance_SBox_Instance_13_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR4_U1 ( .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_1730, LED_128_Instance_addconst_out[52]}), .c ({new_AGEMA_signal_1864, LED_128_Instance_SBox_Instance_13_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR5_U1 ( .a ({new_AGEMA_signal_1864, LED_128_Instance_SBox_Instance_13_L3}), .b ({new_AGEMA_signal_1862, LED_128_Instance_SBox_Instance_13_L0}), .c ({new_AGEMA_signal_1925, LED_128_Instance_SBox_Instance_13_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR6_U1 ( .a ({new_AGEMA_signal_1708, LED_128_Instance_addconst_out[55]}), .b ({new_AGEMA_signal_1729, LED_128_Instance_addconst_out[53]}), .c ({new_AGEMA_signal_1865, LED_128_Instance_SBox_Instance_13_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR9_U1 ( .a ({new_AGEMA_signal_1863, LED_128_Instance_SBox_Instance_13_L1}), .b ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}), .c ({new_AGEMA_signal_1926, LED_128_Instance_SBox_Instance_13_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_U3 ( .a ({new_AGEMA_signal_1789, LED_128_Instance_SBox_Instance_14_L0}), .b ({new_AGEMA_signal_1866, LED_128_Instance_SBox_Instance_14_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_U2 ( .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_1787, LED_128_Instance_SBox_Instance_14_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_U1 ( .a ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_1788, LED_128_Instance_SBox_Instance_14_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR1_U1 ( .a ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .b ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_1789, LED_128_Instance_SBox_Instance_14_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR2_U1 ( .a ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .b ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR3_U1 ( .a ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .c ({new_AGEMA_signal_1867, LED_128_Instance_SBox_Instance_14_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR4_U1 ( .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_1709, LED_128_Instance_addconst_out[56]}), .c ({new_AGEMA_signal_1791, LED_128_Instance_SBox_Instance_14_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR5_U1 ( .a ({new_AGEMA_signal_1791, LED_128_Instance_SBox_Instance_14_L3}), .b ({new_AGEMA_signal_1789, LED_128_Instance_SBox_Instance_14_L0}), .c ({new_AGEMA_signal_1868, LED_128_Instance_SBox_Instance_14_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR6_U1 ( .a ({new_AGEMA_signal_1712, LED_128_Instance_addconst_out[59]}), .b ({new_AGEMA_signal_1710, LED_128_Instance_addconst_out[57]}), .c ({new_AGEMA_signal_1792, LED_128_Instance_SBox_Instance_14_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR9_U1 ( .a ({new_AGEMA_signal_1790, LED_128_Instance_SBox_Instance_14_L1}), .b ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .c ({new_AGEMA_signal_1869, LED_128_Instance_SBox_Instance_14_Q7}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_U3 ( .a ({new_AGEMA_signal_1795, LED_128_Instance_SBox_Instance_15_L0}), .b ({new_AGEMA_signal_1871, LED_128_Instance_SBox_Instance_15_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_U2 ( .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_1793, LED_128_Instance_SBox_Instance_15_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_U1 ( .a ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_1794, LED_128_Instance_SBox_Instance_15_n3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR1_U1 ( .a ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .b ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_1795, LED_128_Instance_SBox_Instance_15_L0}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR2_U1 ( .a ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .b ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR3_U1 ( .a ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .c ({new_AGEMA_signal_1872, LED_128_Instance_SBox_Instance_15_L2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR4_U1 ( .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_1713, LED_128_Instance_addconst_out[60]}), .c ({new_AGEMA_signal_1797, LED_128_Instance_SBox_Instance_15_L3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR5_U1 ( .a ({new_AGEMA_signal_1797, LED_128_Instance_SBox_Instance_15_L3}), .b ({new_AGEMA_signal_1795, LED_128_Instance_SBox_Instance_15_L0}), .c ({new_AGEMA_signal_1873, LED_128_Instance_SBox_Instance_15_Q3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR6_U1 ( .a ({new_AGEMA_signal_1716, LED_128_Instance_addconst_out[63]}), .b ({new_AGEMA_signal_1714, LED_128_Instance_addconst_out[61]}), .c ({new_AGEMA_signal_1798, LED_128_Instance_SBox_Instance_15_L4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR9_U1 ( .a ({new_AGEMA_signal_1796, LED_128_Instance_SBox_Instance_15_L1}), .b ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .c ({new_AGEMA_signal_1874, LED_128_Instance_SBox_Instance_15_Q7}) ) ;
    INV_X1 LED_128_Instance_ks_reg_0__U1 ( .A (LED_128_Instance_ks_reg_0__Q), .ZN (LED_128_Instance_n4) ) ;
    INV_X1 LED_128_Instance_ks_reg_1__U1 ( .A (LED_128_Instance_n26), .ZN (LED_128_Instance_n8) ) ;
    INV_X1 LED_128_Instance_ks_reg_2__U1 ( .A (LED_128_Instance_n25), .ZN (LED_128_Instance_n1) ) ;
    INV_X1 LED_128_Instance_ks_reg_3__U1 ( .A (LED_128_Instance_n2), .ZN (LED_128_Instance_n24) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_0__U1 ( .A (roundconstant[0]), .ZN (LED_128_Instance_n6) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_1__U1 ( .A (roundconstant[1]), .ZN (LED_128_Instance_n29) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_2__U1 ( .A (roundconstant[2]), .ZN (LED_128_Instance_n5) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_3__U1 ( .A (roundconstant[3]), .ZN (LED_128_Instance_n30) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_4__U1 ( .A (roundconstant[4]), .ZN (LED_128_Instance_n28) ) ;
    INV_X1 LED_128_Instance_roundconstant_reg_5__U1 ( .A (roundconstant[5]), .ZN (LED_128_Instance_n27) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L2), .Q (new_AGEMA_signal_2580) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (CLK), .D (new_AGEMA_signal_1877), .Q (new_AGEMA_signal_2582) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L4), .Q (new_AGEMA_signal_2584) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (CLK), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_2586) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L3), .Q (new_AGEMA_signal_2588) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (CLK), .D (new_AGEMA_signal_1722), .Q (new_AGEMA_signal_2590) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L2), .Q (new_AGEMA_signal_2592) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (CLK), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_2594) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L4), .Q (new_AGEMA_signal_2596) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (CLK), .D (new_AGEMA_signal_1807), .Q (new_AGEMA_signal_2598) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L3), .Q (new_AGEMA_signal_2600) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (CLK), .D (new_AGEMA_signal_1806), .Q (new_AGEMA_signal_2602) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L2), .Q (new_AGEMA_signal_2604) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (CLK), .D (new_AGEMA_signal_1809), .Q (new_AGEMA_signal_2606) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L4), .Q (new_AGEMA_signal_2608) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (CLK), .D (new_AGEMA_signal_1751), .Q (new_AGEMA_signal_2610) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L3), .Q (new_AGEMA_signal_2612) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (CLK), .D (new_AGEMA_signal_1750), .Q (new_AGEMA_signal_2614) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L2), .Q (new_AGEMA_signal_2616) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (CLK), .D (new_AGEMA_signal_1814), .Q (new_AGEMA_signal_2618) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L4), .Q (new_AGEMA_signal_2620) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (CLK), .D (new_AGEMA_signal_1757), .Q (new_AGEMA_signal_2622) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L3), .Q (new_AGEMA_signal_2624) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (CLK), .D (new_AGEMA_signal_1756), .Q (new_AGEMA_signal_2626) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L2), .Q (new_AGEMA_signal_2628) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (CLK), .D (new_AGEMA_signal_1891), .Q (new_AGEMA_signal_2630) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L4), .Q (new_AGEMA_signal_2632) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (CLK), .D (new_AGEMA_signal_1821), .Q (new_AGEMA_signal_2634) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L3), .Q (new_AGEMA_signal_2636) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (CLK), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_2638) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L2), .Q (new_AGEMA_signal_2640) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (CLK), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_2642) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L4), .Q (new_AGEMA_signal_2644) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (CLK), .D (new_AGEMA_signal_1826), .Q (new_AGEMA_signal_2646) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L3), .Q (new_AGEMA_signal_2648) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (CLK), .D (new_AGEMA_signal_1825), .Q (new_AGEMA_signal_2650) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L2), .Q (new_AGEMA_signal_2652) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (CLK), .D (new_AGEMA_signal_1828), .Q (new_AGEMA_signal_2654) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L4), .Q (new_AGEMA_signal_2656) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (CLK), .D (new_AGEMA_signal_1764), .Q (new_AGEMA_signal_2658) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L3), .Q (new_AGEMA_signal_2660) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (CLK), .D (new_AGEMA_signal_1763), .Q (new_AGEMA_signal_2662) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L2), .Q (new_AGEMA_signal_2664) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (CLK), .D (new_AGEMA_signal_1833), .Q (new_AGEMA_signal_2666) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L4), .Q (new_AGEMA_signal_2668) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (CLK), .D (new_AGEMA_signal_1770), .Q (new_AGEMA_signal_2670) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L3), .Q (new_AGEMA_signal_2672) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (CLK), .D (new_AGEMA_signal_1769), .Q (new_AGEMA_signal_2674) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L2), .Q (new_AGEMA_signal_2676) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (CLK), .D (new_AGEMA_signal_1905), .Q (new_AGEMA_signal_2678) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L4), .Q (new_AGEMA_signal_2680) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (CLK), .D (new_AGEMA_signal_1840), .Q (new_AGEMA_signal_2682) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L3), .Q (new_AGEMA_signal_2684) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (CLK), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_2686) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L2), .Q (new_AGEMA_signal_2688) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (CLK), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_2690) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L4), .Q (new_AGEMA_signal_2692) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (CLK), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_2694) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L3), .Q (new_AGEMA_signal_2696) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (CLK), .D (new_AGEMA_signal_1773), .Q (new_AGEMA_signal_2698) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L2), .Q (new_AGEMA_signal_2700) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (CLK), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_2702) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L4), .Q (new_AGEMA_signal_2704) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (CLK), .D (new_AGEMA_signal_1779), .Q (new_AGEMA_signal_2706) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L3), .Q (new_AGEMA_signal_2708) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (CLK), .D (new_AGEMA_signal_1778), .Q (new_AGEMA_signal_2710) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L2), .Q (new_AGEMA_signal_2712) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (CLK), .D (new_AGEMA_signal_1851), .Q (new_AGEMA_signal_2714) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L4), .Q (new_AGEMA_signal_2716) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (CLK), .D (new_AGEMA_signal_1785), .Q (new_AGEMA_signal_2718) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L3), .Q (new_AGEMA_signal_2720) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (CLK), .D (new_AGEMA_signal_1784), .Q (new_AGEMA_signal_2722) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L2), .Q (new_AGEMA_signal_2724) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (CLK), .D (new_AGEMA_signal_1919), .Q (new_AGEMA_signal_2726) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L4), .Q (new_AGEMA_signal_2728) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (CLK), .D (new_AGEMA_signal_1860), .Q (new_AGEMA_signal_2730) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L3), .Q (new_AGEMA_signal_2732) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (CLK), .D (new_AGEMA_signal_1859), .Q (new_AGEMA_signal_2734) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L2), .Q (new_AGEMA_signal_2736) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (CLK), .D (new_AGEMA_signal_1924), .Q (new_AGEMA_signal_2738) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L4), .Q (new_AGEMA_signal_2740) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (CLK), .D (new_AGEMA_signal_1865), .Q (new_AGEMA_signal_2742) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L3), .Q (new_AGEMA_signal_2744) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (CLK), .D (new_AGEMA_signal_1864), .Q (new_AGEMA_signal_2746) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L2), .Q (new_AGEMA_signal_2748) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (CLK), .D (new_AGEMA_signal_1867), .Q (new_AGEMA_signal_2750) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L4), .Q (new_AGEMA_signal_2752) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (CLK), .D (new_AGEMA_signal_1792), .Q (new_AGEMA_signal_2754) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L3), .Q (new_AGEMA_signal_2756) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (CLK), .D (new_AGEMA_signal_1791), .Q (new_AGEMA_signal_2758) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L2), .Q (new_AGEMA_signal_2760) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (CLK), .D (new_AGEMA_signal_1872), .Q (new_AGEMA_signal_2762) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L4), .Q (new_AGEMA_signal_2764) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (CLK), .D (new_AGEMA_signal_1798), .Q (new_AGEMA_signal_2766) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L3), .Q (new_AGEMA_signal_2768) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (CLK), .D (new_AGEMA_signal_1797), .Q (new_AGEMA_signal_2770) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (CLK), .D (LED_128_Instance_MUX_state0_n9), .Q (new_AGEMA_signal_2772) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_0_), .Q (new_AGEMA_signal_2776) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (CLK), .D (new_AGEMA_signal_1546), .Q (new_AGEMA_signal_2780) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_1_), .Q (new_AGEMA_signal_2784) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (CLK), .D (new_AGEMA_signal_1666), .Q (new_AGEMA_signal_2788) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (CLK), .D (LED_128_Instance_MUX_state0_n8), .Q (new_AGEMA_signal_2792) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_2_), .Q (new_AGEMA_signal_2796) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (CLK), .D (new_AGEMA_signal_1667), .Q (new_AGEMA_signal_2800) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (CLK), .D (LED_128_Instance_MUX_state0_n10), .Q (new_AGEMA_signal_2804) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_3_), .Q (new_AGEMA_signal_2808) ) ;
    buf_clk new_AGEMA_reg_buffer_1360 ( .C (CLK), .D (new_AGEMA_signal_1547), .Q (new_AGEMA_signal_2812) ) ;
    buf_clk new_AGEMA_reg_buffer_1364 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_4_), .Q (new_AGEMA_signal_2816) ) ;
    buf_clk new_AGEMA_reg_buffer_1368 ( .C (CLK), .D (new_AGEMA_signal_1668), .Q (new_AGEMA_signal_2820) ) ;
    buf_clk new_AGEMA_reg_buffer_1372 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_5_), .Q (new_AGEMA_signal_2824) ) ;
    buf_clk new_AGEMA_reg_buffer_1376 ( .C (CLK), .D (new_AGEMA_signal_1669), .Q (new_AGEMA_signal_2828) ) ;
    buf_clk new_AGEMA_reg_buffer_1380 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_6_), .Q (new_AGEMA_signal_2832) ) ;
    buf_clk new_AGEMA_reg_buffer_1384 ( .C (CLK), .D (new_AGEMA_signal_1670), .Q (new_AGEMA_signal_2836) ) ;
    buf_clk new_AGEMA_reg_buffer_1388 ( .C (CLK), .D (LED_128_Instance_addconst_out[7]), .Q (new_AGEMA_signal_2840) ) ;
    buf_clk new_AGEMA_reg_buffer_1392 ( .C (CLK), .D (new_AGEMA_signal_1671), .Q (new_AGEMA_signal_2844) ) ;
    buf_clk new_AGEMA_reg_buffer_1396 ( .C (CLK), .D (LED_128_Instance_addconst_out[8]), .Q (new_AGEMA_signal_2848) ) ;
    buf_clk new_AGEMA_reg_buffer_1400 ( .C (CLK), .D (new_AGEMA_signal_1672), .Q (new_AGEMA_signal_2852) ) ;
    buf_clk new_AGEMA_reg_buffer_1404 ( .C (CLK), .D (LED_128_Instance_addconst_out[9]), .Q (new_AGEMA_signal_2856) ) ;
    buf_clk new_AGEMA_reg_buffer_1408 ( .C (CLK), .D (new_AGEMA_signal_1673), .Q (new_AGEMA_signal_2860) ) ;
    buf_clk new_AGEMA_reg_buffer_1412 ( .C (CLK), .D (LED_128_Instance_addconst_out[10]), .Q (new_AGEMA_signal_2864) ) ;
    buf_clk new_AGEMA_reg_buffer_1416 ( .C (CLK), .D (new_AGEMA_signal_1674), .Q (new_AGEMA_signal_2868) ) ;
    buf_clk new_AGEMA_reg_buffer_1420 ( .C (CLK), .D (LED_128_Instance_addconst_out[11]), .Q (new_AGEMA_signal_2872) ) ;
    buf_clk new_AGEMA_reg_buffer_1424 ( .C (CLK), .D (new_AGEMA_signal_1675), .Q (new_AGEMA_signal_2876) ) ;
    buf_clk new_AGEMA_reg_buffer_1428 ( .C (CLK), .D (LED_128_Instance_addconst_out[12]), .Q (new_AGEMA_signal_2880) ) ;
    buf_clk new_AGEMA_reg_buffer_1432 ( .C (CLK), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_2884) ) ;
    buf_clk new_AGEMA_reg_buffer_1436 ( .C (CLK), .D (LED_128_Instance_addconst_out[13]), .Q (new_AGEMA_signal_2888) ) ;
    buf_clk new_AGEMA_reg_buffer_1440 ( .C (CLK), .D (new_AGEMA_signal_1677), .Q (new_AGEMA_signal_2892) ) ;
    buf_clk new_AGEMA_reg_buffer_1444 ( .C (CLK), .D (LED_128_Instance_addconst_out[14]), .Q (new_AGEMA_signal_2896) ) ;
    buf_clk new_AGEMA_reg_buffer_1448 ( .C (CLK), .D (new_AGEMA_signal_1678), .Q (new_AGEMA_signal_2900) ) ;
    buf_clk new_AGEMA_reg_buffer_1452 ( .C (CLK), .D (LED_128_Instance_addconst_out[15]), .Q (new_AGEMA_signal_2904) ) ;
    buf_clk new_AGEMA_reg_buffer_1456 ( .C (CLK), .D (new_AGEMA_signal_1679), .Q (new_AGEMA_signal_2908) ) ;
    buf_clk new_AGEMA_reg_buffer_1460 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_16_), .Q (new_AGEMA_signal_2912) ) ;
    buf_clk new_AGEMA_reg_buffer_1464 ( .C (CLK), .D (new_AGEMA_signal_1548), .Q (new_AGEMA_signal_2916) ) ;
    buf_clk new_AGEMA_reg_buffer_1468 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_17_), .Q (new_AGEMA_signal_2920) ) ;
    buf_clk new_AGEMA_reg_buffer_1472 ( .C (CLK), .D (new_AGEMA_signal_1680), .Q (new_AGEMA_signal_2924) ) ;
    buf_clk new_AGEMA_reg_buffer_1476 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_18_), .Q (new_AGEMA_signal_2928) ) ;
    buf_clk new_AGEMA_reg_buffer_1480 ( .C (CLK), .D (new_AGEMA_signal_1681), .Q (new_AGEMA_signal_2932) ) ;
    buf_clk new_AGEMA_reg_buffer_1484 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_19_), .Q (new_AGEMA_signal_2936) ) ;
    buf_clk new_AGEMA_reg_buffer_1488 ( .C (CLK), .D (new_AGEMA_signal_1549), .Q (new_AGEMA_signal_2940) ) ;
    buf_clk new_AGEMA_reg_buffer_1492 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_20_), .Q (new_AGEMA_signal_2944) ) ;
    buf_clk new_AGEMA_reg_buffer_1496 ( .C (CLK), .D (new_AGEMA_signal_1682), .Q (new_AGEMA_signal_2948) ) ;
    buf_clk new_AGEMA_reg_buffer_1500 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_21_), .Q (new_AGEMA_signal_2952) ) ;
    buf_clk new_AGEMA_reg_buffer_1504 ( .C (CLK), .D (new_AGEMA_signal_1683), .Q (new_AGEMA_signal_2956) ) ;
    buf_clk new_AGEMA_reg_buffer_1508 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_22_), .Q (new_AGEMA_signal_2960) ) ;
    buf_clk new_AGEMA_reg_buffer_1512 ( .C (CLK), .D (new_AGEMA_signal_1550), .Q (new_AGEMA_signal_2964) ) ;
    buf_clk new_AGEMA_reg_buffer_1516 ( .C (CLK), .D (LED_128_Instance_addconst_out[23]), .Q (new_AGEMA_signal_2968) ) ;
    buf_clk new_AGEMA_reg_buffer_1520 ( .C (CLK), .D (new_AGEMA_signal_1684), .Q (new_AGEMA_signal_2972) ) ;
    buf_clk new_AGEMA_reg_buffer_1524 ( .C (CLK), .D (LED_128_Instance_addconst_out[24]), .Q (new_AGEMA_signal_2976) ) ;
    buf_clk new_AGEMA_reg_buffer_1528 ( .C (CLK), .D (new_AGEMA_signal_1551), .Q (new_AGEMA_signal_2980) ) ;
    buf_clk new_AGEMA_reg_buffer_1532 ( .C (CLK), .D (LED_128_Instance_addconst_out[25]), .Q (new_AGEMA_signal_2984) ) ;
    buf_clk new_AGEMA_reg_buffer_1536 ( .C (CLK), .D (new_AGEMA_signal_1685), .Q (new_AGEMA_signal_2988) ) ;
    buf_clk new_AGEMA_reg_buffer_1540 ( .C (CLK), .D (LED_128_Instance_addconst_out[26]), .Q (new_AGEMA_signal_2992) ) ;
    buf_clk new_AGEMA_reg_buffer_1544 ( .C (CLK), .D (new_AGEMA_signal_1552), .Q (new_AGEMA_signal_2996) ) ;
    buf_clk new_AGEMA_reg_buffer_1548 ( .C (CLK), .D (LED_128_Instance_addconst_out[27]), .Q (new_AGEMA_signal_3000) ) ;
    buf_clk new_AGEMA_reg_buffer_1552 ( .C (CLK), .D (new_AGEMA_signal_1686), .Q (new_AGEMA_signal_3004) ) ;
    buf_clk new_AGEMA_reg_buffer_1556 ( .C (CLK), .D (LED_128_Instance_addconst_out[28]), .Q (new_AGEMA_signal_3008) ) ;
    buf_clk new_AGEMA_reg_buffer_1560 ( .C (CLK), .D (new_AGEMA_signal_1655), .Q (new_AGEMA_signal_3012) ) ;
    buf_clk new_AGEMA_reg_buffer_1564 ( .C (CLK), .D (LED_128_Instance_addconst_out[29]), .Q (new_AGEMA_signal_3016) ) ;
    buf_clk new_AGEMA_reg_buffer_1568 ( .C (CLK), .D (new_AGEMA_signal_1687), .Q (new_AGEMA_signal_3020) ) ;
    buf_clk new_AGEMA_reg_buffer_1572 ( .C (CLK), .D (LED_128_Instance_addconst_out[30]), .Q (new_AGEMA_signal_3024) ) ;
    buf_clk new_AGEMA_reg_buffer_1576 ( .C (CLK), .D (new_AGEMA_signal_1688), .Q (new_AGEMA_signal_3028) ) ;
    buf_clk new_AGEMA_reg_buffer_1580 ( .C (CLK), .D (LED_128_Instance_addconst_out[31]), .Q (new_AGEMA_signal_3032) ) ;
    buf_clk new_AGEMA_reg_buffer_1584 ( .C (CLK), .D (new_AGEMA_signal_1689), .Q (new_AGEMA_signal_3036) ) ;
    buf_clk new_AGEMA_reg_buffer_1588 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_32_), .Q (new_AGEMA_signal_3040) ) ;
    buf_clk new_AGEMA_reg_buffer_1592 ( .C (CLK), .D (new_AGEMA_signal_1656), .Q (new_AGEMA_signal_3044) ) ;
    buf_clk new_AGEMA_reg_buffer_1596 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_33_), .Q (new_AGEMA_signal_3048) ) ;
    buf_clk new_AGEMA_reg_buffer_1600 ( .C (CLK), .D (new_AGEMA_signal_1690), .Q (new_AGEMA_signal_3052) ) ;
    buf_clk new_AGEMA_reg_buffer_1604 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_34_), .Q (new_AGEMA_signal_3056) ) ;
    buf_clk new_AGEMA_reg_buffer_1608 ( .C (CLK), .D (new_AGEMA_signal_1657), .Q (new_AGEMA_signal_3060) ) ;
    buf_clk new_AGEMA_reg_buffer_1612 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_35_), .Q (new_AGEMA_signal_3064) ) ;
    buf_clk new_AGEMA_reg_buffer_1616 ( .C (CLK), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_3068) ) ;
    buf_clk new_AGEMA_reg_buffer_1620 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_36_), .Q (new_AGEMA_signal_3072) ) ;
    buf_clk new_AGEMA_reg_buffer_1624 ( .C (CLK), .D (new_AGEMA_signal_1659), .Q (new_AGEMA_signal_3076) ) ;
    buf_clk new_AGEMA_reg_buffer_1628 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_37_), .Q (new_AGEMA_signal_3080) ) ;
    buf_clk new_AGEMA_reg_buffer_1632 ( .C (CLK), .D (new_AGEMA_signal_1691), .Q (new_AGEMA_signal_3084) ) ;
    buf_clk new_AGEMA_reg_buffer_1636 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_38_), .Q (new_AGEMA_signal_3088) ) ;
    buf_clk new_AGEMA_reg_buffer_1640 ( .C (CLK), .D (new_AGEMA_signal_1692), .Q (new_AGEMA_signal_3092) ) ;
    buf_clk new_AGEMA_reg_buffer_1644 ( .C (CLK), .D (LED_128_Instance_addconst_out[39]), .Q (new_AGEMA_signal_3096) ) ;
    buf_clk new_AGEMA_reg_buffer_1648 ( .C (CLK), .D (new_AGEMA_signal_1660), .Q (new_AGEMA_signal_3100) ) ;
    buf_clk new_AGEMA_reg_buffer_1652 ( .C (CLK), .D (LED_128_Instance_addconst_out[40]), .Q (new_AGEMA_signal_3104) ) ;
    buf_clk new_AGEMA_reg_buffer_1656 ( .C (CLK), .D (new_AGEMA_signal_1693), .Q (new_AGEMA_signal_3108) ) ;
    buf_clk new_AGEMA_reg_buffer_1660 ( .C (CLK), .D (LED_128_Instance_addconst_out[41]), .Q (new_AGEMA_signal_3112) ) ;
    buf_clk new_AGEMA_reg_buffer_1664 ( .C (CLK), .D (new_AGEMA_signal_1694), .Q (new_AGEMA_signal_3116) ) ;
    buf_clk new_AGEMA_reg_buffer_1668 ( .C (CLK), .D (LED_128_Instance_addconst_out[42]), .Q (new_AGEMA_signal_3120) ) ;
    buf_clk new_AGEMA_reg_buffer_1672 ( .C (CLK), .D (new_AGEMA_signal_1695), .Q (new_AGEMA_signal_3124) ) ;
    buf_clk new_AGEMA_reg_buffer_1676 ( .C (CLK), .D (LED_128_Instance_n22), .Q (new_AGEMA_signal_3128) ) ;
    buf_clk new_AGEMA_reg_buffer_1680 ( .C (CLK), .D (LED_128_Instance_addconst_out[43]), .Q (new_AGEMA_signal_3132) ) ;
    buf_clk new_AGEMA_reg_buffer_1684 ( .C (CLK), .D (new_AGEMA_signal_1696), .Q (new_AGEMA_signal_3136) ) ;
    buf_clk new_AGEMA_reg_buffer_1688 ( .C (CLK), .D (LED_128_Instance_addconst_out[44]), .Q (new_AGEMA_signal_3140) ) ;
    buf_clk new_AGEMA_reg_buffer_1692 ( .C (CLK), .D (new_AGEMA_signal_1697), .Q (new_AGEMA_signal_3144) ) ;
    buf_clk new_AGEMA_reg_buffer_1696 ( .C (CLK), .D (LED_128_Instance_addconst_out[45]), .Q (new_AGEMA_signal_3148) ) ;
    buf_clk new_AGEMA_reg_buffer_1700 ( .C (CLK), .D (new_AGEMA_signal_1698), .Q (new_AGEMA_signal_3152) ) ;
    buf_clk new_AGEMA_reg_buffer_1704 ( .C (CLK), .D (LED_128_Instance_addconst_out[46]), .Q (new_AGEMA_signal_3156) ) ;
    buf_clk new_AGEMA_reg_buffer_1708 ( .C (CLK), .D (new_AGEMA_signal_1699), .Q (new_AGEMA_signal_3160) ) ;
    buf_clk new_AGEMA_reg_buffer_1712 ( .C (CLK), .D (LED_128_Instance_addconst_out[47]), .Q (new_AGEMA_signal_3164) ) ;
    buf_clk new_AGEMA_reg_buffer_1716 ( .C (CLK), .D (new_AGEMA_signal_1700), .Q (new_AGEMA_signal_3168) ) ;
    buf_clk new_AGEMA_reg_buffer_1720 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_48_), .Q (new_AGEMA_signal_3172) ) ;
    buf_clk new_AGEMA_reg_buffer_1724 ( .C (CLK), .D (new_AGEMA_signal_1701), .Q (new_AGEMA_signal_3176) ) ;
    buf_clk new_AGEMA_reg_buffer_1728 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_49_), .Q (new_AGEMA_signal_3180) ) ;
    buf_clk new_AGEMA_reg_buffer_1732 ( .C (CLK), .D (new_AGEMA_signal_1702), .Q (new_AGEMA_signal_3184) ) ;
    buf_clk new_AGEMA_reg_buffer_1736 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_50_), .Q (new_AGEMA_signal_3188) ) ;
    buf_clk new_AGEMA_reg_buffer_1740 ( .C (CLK), .D (new_AGEMA_signal_1703), .Q (new_AGEMA_signal_3192) ) ;
    buf_clk new_AGEMA_reg_buffer_1744 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_51_), .Q (new_AGEMA_signal_3196) ) ;
    buf_clk new_AGEMA_reg_buffer_1748 ( .C (CLK), .D (new_AGEMA_signal_1704), .Q (new_AGEMA_signal_3200) ) ;
    buf_clk new_AGEMA_reg_buffer_1752 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_52_), .Q (new_AGEMA_signal_3204) ) ;
    buf_clk new_AGEMA_reg_buffer_1756 ( .C (CLK), .D (new_AGEMA_signal_1705), .Q (new_AGEMA_signal_3208) ) ;
    buf_clk new_AGEMA_reg_buffer_1760 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_53_), .Q (new_AGEMA_signal_3212) ) ;
    buf_clk new_AGEMA_reg_buffer_1764 ( .C (CLK), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_3216) ) ;
    buf_clk new_AGEMA_reg_buffer_1768 ( .C (CLK), .D (LED_128_Instance_addroundkey_out_54_), .Q (new_AGEMA_signal_3220) ) ;
    buf_clk new_AGEMA_reg_buffer_1772 ( .C (CLK), .D (new_AGEMA_signal_1707), .Q (new_AGEMA_signal_3224) ) ;
    buf_clk new_AGEMA_reg_buffer_1776 ( .C (CLK), .D (LED_128_Instance_addconst_out[55]), .Q (new_AGEMA_signal_3228) ) ;
    buf_clk new_AGEMA_reg_buffer_1780 ( .C (CLK), .D (new_AGEMA_signal_1708), .Q (new_AGEMA_signal_3232) ) ;
    buf_clk new_AGEMA_reg_buffer_1784 ( .C (CLK), .D (LED_128_Instance_addconst_out[56]), .Q (new_AGEMA_signal_3236) ) ;
    buf_clk new_AGEMA_reg_buffer_1788 ( .C (CLK), .D (new_AGEMA_signal_1709), .Q (new_AGEMA_signal_3240) ) ;
    buf_clk new_AGEMA_reg_buffer_1792 ( .C (CLK), .D (LED_128_Instance_addconst_out[57]), .Q (new_AGEMA_signal_3244) ) ;
    buf_clk new_AGEMA_reg_buffer_1796 ( .C (CLK), .D (new_AGEMA_signal_1710), .Q (new_AGEMA_signal_3248) ) ;
    buf_clk new_AGEMA_reg_buffer_1800 ( .C (CLK), .D (LED_128_Instance_addconst_out[58]), .Q (new_AGEMA_signal_3252) ) ;
    buf_clk new_AGEMA_reg_buffer_1804 ( .C (CLK), .D (new_AGEMA_signal_1711), .Q (new_AGEMA_signal_3256) ) ;
    buf_clk new_AGEMA_reg_buffer_1808 ( .C (CLK), .D (LED_128_Instance_addconst_out[59]), .Q (new_AGEMA_signal_3260) ) ;
    buf_clk new_AGEMA_reg_buffer_1812 ( .C (CLK), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_3264) ) ;
    buf_clk new_AGEMA_reg_buffer_1816 ( .C (CLK), .D (LED_128_Instance_addconst_out[60]), .Q (new_AGEMA_signal_3268) ) ;
    buf_clk new_AGEMA_reg_buffer_1820 ( .C (CLK), .D (new_AGEMA_signal_1713), .Q (new_AGEMA_signal_3272) ) ;
    buf_clk new_AGEMA_reg_buffer_1824 ( .C (CLK), .D (LED_128_Instance_addconst_out[61]), .Q (new_AGEMA_signal_3276) ) ;
    buf_clk new_AGEMA_reg_buffer_1828 ( .C (CLK), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_3280) ) ;
    buf_clk new_AGEMA_reg_buffer_1832 ( .C (CLK), .D (LED_128_Instance_addconst_out[62]), .Q (new_AGEMA_signal_3284) ) ;
    buf_clk new_AGEMA_reg_buffer_1836 ( .C (CLK), .D (new_AGEMA_signal_1715), .Q (new_AGEMA_signal_3288) ) ;
    buf_clk new_AGEMA_reg_buffer_1840 ( .C (CLK), .D (LED_128_Instance_addconst_out[63]), .Q (new_AGEMA_signal_3292) ) ;
    buf_clk new_AGEMA_reg_buffer_1844 ( .C (CLK), .D (new_AGEMA_signal_1716), .Q (new_AGEMA_signal_3296) ) ;
    buf_clk new_AGEMA_reg_buffer_1848 ( .C (CLK), .D (IN_reset), .Q (new_AGEMA_signal_3300) ) ;
    buf_clk new_AGEMA_reg_buffer_1852 ( .C (CLK), .D (IN_plaintext_s0[0]), .Q (new_AGEMA_signal_3304) ) ;
    buf_clk new_AGEMA_reg_buffer_1856 ( .C (CLK), .D (IN_plaintext_s1[0]), .Q (new_AGEMA_signal_3308) ) ;
    buf_clk new_AGEMA_reg_buffer_1860 ( .C (CLK), .D (IN_plaintext_s0[1]), .Q (new_AGEMA_signal_3312) ) ;
    buf_clk new_AGEMA_reg_buffer_1864 ( .C (CLK), .D (IN_plaintext_s1[1]), .Q (new_AGEMA_signal_3316) ) ;
    buf_clk new_AGEMA_reg_buffer_1868 ( .C (CLK), .D (IN_plaintext_s0[2]), .Q (new_AGEMA_signal_3320) ) ;
    buf_clk new_AGEMA_reg_buffer_1872 ( .C (CLK), .D (IN_plaintext_s1[2]), .Q (new_AGEMA_signal_3324) ) ;
    buf_clk new_AGEMA_reg_buffer_1876 ( .C (CLK), .D (IN_plaintext_s0[3]), .Q (new_AGEMA_signal_3328) ) ;
    buf_clk new_AGEMA_reg_buffer_1880 ( .C (CLK), .D (IN_plaintext_s1[3]), .Q (new_AGEMA_signal_3332) ) ;
    buf_clk new_AGEMA_reg_buffer_1884 ( .C (CLK), .D (IN_plaintext_s0[4]), .Q (new_AGEMA_signal_3336) ) ;
    buf_clk new_AGEMA_reg_buffer_1888 ( .C (CLK), .D (IN_plaintext_s1[4]), .Q (new_AGEMA_signal_3340) ) ;
    buf_clk new_AGEMA_reg_buffer_1892 ( .C (CLK), .D (IN_plaintext_s0[5]), .Q (new_AGEMA_signal_3344) ) ;
    buf_clk new_AGEMA_reg_buffer_1896 ( .C (CLK), .D (IN_plaintext_s1[5]), .Q (new_AGEMA_signal_3348) ) ;
    buf_clk new_AGEMA_reg_buffer_1900 ( .C (CLK), .D (IN_plaintext_s0[6]), .Q (new_AGEMA_signal_3352) ) ;
    buf_clk new_AGEMA_reg_buffer_1904 ( .C (CLK), .D (IN_plaintext_s1[6]), .Q (new_AGEMA_signal_3356) ) ;
    buf_clk new_AGEMA_reg_buffer_1908 ( .C (CLK), .D (IN_plaintext_s0[7]), .Q (new_AGEMA_signal_3360) ) ;
    buf_clk new_AGEMA_reg_buffer_1912 ( .C (CLK), .D (IN_plaintext_s1[7]), .Q (new_AGEMA_signal_3364) ) ;
    buf_clk new_AGEMA_reg_buffer_1916 ( .C (CLK), .D (IN_plaintext_s0[8]), .Q (new_AGEMA_signal_3368) ) ;
    buf_clk new_AGEMA_reg_buffer_1920 ( .C (CLK), .D (IN_plaintext_s1[8]), .Q (new_AGEMA_signal_3372) ) ;
    buf_clk new_AGEMA_reg_buffer_1924 ( .C (CLK), .D (IN_plaintext_s0[9]), .Q (new_AGEMA_signal_3376) ) ;
    buf_clk new_AGEMA_reg_buffer_1928 ( .C (CLK), .D (IN_plaintext_s1[9]), .Q (new_AGEMA_signal_3380) ) ;
    buf_clk new_AGEMA_reg_buffer_1932 ( .C (CLK), .D (IN_plaintext_s0[10]), .Q (new_AGEMA_signal_3384) ) ;
    buf_clk new_AGEMA_reg_buffer_1936 ( .C (CLK), .D (IN_plaintext_s1[10]), .Q (new_AGEMA_signal_3388) ) ;
    buf_clk new_AGEMA_reg_buffer_1940 ( .C (CLK), .D (IN_plaintext_s0[11]), .Q (new_AGEMA_signal_3392) ) ;
    buf_clk new_AGEMA_reg_buffer_1944 ( .C (CLK), .D (IN_plaintext_s1[11]), .Q (new_AGEMA_signal_3396) ) ;
    buf_clk new_AGEMA_reg_buffer_1948 ( .C (CLK), .D (IN_plaintext_s0[12]), .Q (new_AGEMA_signal_3400) ) ;
    buf_clk new_AGEMA_reg_buffer_1952 ( .C (CLK), .D (IN_plaintext_s1[12]), .Q (new_AGEMA_signal_3404) ) ;
    buf_clk new_AGEMA_reg_buffer_1956 ( .C (CLK), .D (IN_plaintext_s0[13]), .Q (new_AGEMA_signal_3408) ) ;
    buf_clk new_AGEMA_reg_buffer_1960 ( .C (CLK), .D (IN_plaintext_s1[13]), .Q (new_AGEMA_signal_3412) ) ;
    buf_clk new_AGEMA_reg_buffer_1964 ( .C (CLK), .D (IN_plaintext_s0[14]), .Q (new_AGEMA_signal_3416) ) ;
    buf_clk new_AGEMA_reg_buffer_1968 ( .C (CLK), .D (IN_plaintext_s1[14]), .Q (new_AGEMA_signal_3420) ) ;
    buf_clk new_AGEMA_reg_buffer_1972 ( .C (CLK), .D (IN_plaintext_s0[15]), .Q (new_AGEMA_signal_3424) ) ;
    buf_clk new_AGEMA_reg_buffer_1976 ( .C (CLK), .D (IN_plaintext_s1[15]), .Q (new_AGEMA_signal_3428) ) ;
    buf_clk new_AGEMA_reg_buffer_1980 ( .C (CLK), .D (IN_plaintext_s0[16]), .Q (new_AGEMA_signal_3432) ) ;
    buf_clk new_AGEMA_reg_buffer_1984 ( .C (CLK), .D (IN_plaintext_s1[16]), .Q (new_AGEMA_signal_3436) ) ;
    buf_clk new_AGEMA_reg_buffer_1988 ( .C (CLK), .D (IN_plaintext_s0[17]), .Q (new_AGEMA_signal_3440) ) ;
    buf_clk new_AGEMA_reg_buffer_1992 ( .C (CLK), .D (IN_plaintext_s1[17]), .Q (new_AGEMA_signal_3444) ) ;
    buf_clk new_AGEMA_reg_buffer_1996 ( .C (CLK), .D (IN_plaintext_s0[18]), .Q (new_AGEMA_signal_3448) ) ;
    buf_clk new_AGEMA_reg_buffer_2000 ( .C (CLK), .D (IN_plaintext_s1[18]), .Q (new_AGEMA_signal_3452) ) ;
    buf_clk new_AGEMA_reg_buffer_2004 ( .C (CLK), .D (IN_plaintext_s0[19]), .Q (new_AGEMA_signal_3456) ) ;
    buf_clk new_AGEMA_reg_buffer_2008 ( .C (CLK), .D (IN_plaintext_s1[19]), .Q (new_AGEMA_signal_3460) ) ;
    buf_clk new_AGEMA_reg_buffer_2012 ( .C (CLK), .D (IN_plaintext_s0[20]), .Q (new_AGEMA_signal_3464) ) ;
    buf_clk new_AGEMA_reg_buffer_2016 ( .C (CLK), .D (IN_plaintext_s1[20]), .Q (new_AGEMA_signal_3468) ) ;
    buf_clk new_AGEMA_reg_buffer_2020 ( .C (CLK), .D (IN_plaintext_s0[21]), .Q (new_AGEMA_signal_3472) ) ;
    buf_clk new_AGEMA_reg_buffer_2024 ( .C (CLK), .D (IN_plaintext_s1[21]), .Q (new_AGEMA_signal_3476) ) ;
    buf_clk new_AGEMA_reg_buffer_2028 ( .C (CLK), .D (IN_plaintext_s0[22]), .Q (new_AGEMA_signal_3480) ) ;
    buf_clk new_AGEMA_reg_buffer_2032 ( .C (CLK), .D (IN_plaintext_s1[22]), .Q (new_AGEMA_signal_3484) ) ;
    buf_clk new_AGEMA_reg_buffer_2036 ( .C (CLK), .D (IN_plaintext_s0[23]), .Q (new_AGEMA_signal_3488) ) ;
    buf_clk new_AGEMA_reg_buffer_2040 ( .C (CLK), .D (IN_plaintext_s1[23]), .Q (new_AGEMA_signal_3492) ) ;
    buf_clk new_AGEMA_reg_buffer_2044 ( .C (CLK), .D (IN_plaintext_s0[24]), .Q (new_AGEMA_signal_3496) ) ;
    buf_clk new_AGEMA_reg_buffer_2048 ( .C (CLK), .D (IN_plaintext_s1[24]), .Q (new_AGEMA_signal_3500) ) ;
    buf_clk new_AGEMA_reg_buffer_2052 ( .C (CLK), .D (IN_plaintext_s0[25]), .Q (new_AGEMA_signal_3504) ) ;
    buf_clk new_AGEMA_reg_buffer_2056 ( .C (CLK), .D (IN_plaintext_s1[25]), .Q (new_AGEMA_signal_3508) ) ;
    buf_clk new_AGEMA_reg_buffer_2060 ( .C (CLK), .D (IN_plaintext_s0[26]), .Q (new_AGEMA_signal_3512) ) ;
    buf_clk new_AGEMA_reg_buffer_2064 ( .C (CLK), .D (IN_plaintext_s1[26]), .Q (new_AGEMA_signal_3516) ) ;
    buf_clk new_AGEMA_reg_buffer_2068 ( .C (CLK), .D (IN_plaintext_s0[27]), .Q (new_AGEMA_signal_3520) ) ;
    buf_clk new_AGEMA_reg_buffer_2072 ( .C (CLK), .D (IN_plaintext_s1[27]), .Q (new_AGEMA_signal_3524) ) ;
    buf_clk new_AGEMA_reg_buffer_2076 ( .C (CLK), .D (IN_plaintext_s0[28]), .Q (new_AGEMA_signal_3528) ) ;
    buf_clk new_AGEMA_reg_buffer_2080 ( .C (CLK), .D (IN_plaintext_s1[28]), .Q (new_AGEMA_signal_3532) ) ;
    buf_clk new_AGEMA_reg_buffer_2084 ( .C (CLK), .D (IN_plaintext_s0[29]), .Q (new_AGEMA_signal_3536) ) ;
    buf_clk new_AGEMA_reg_buffer_2088 ( .C (CLK), .D (IN_plaintext_s1[29]), .Q (new_AGEMA_signal_3540) ) ;
    buf_clk new_AGEMA_reg_buffer_2092 ( .C (CLK), .D (IN_plaintext_s0[30]), .Q (new_AGEMA_signal_3544) ) ;
    buf_clk new_AGEMA_reg_buffer_2096 ( .C (CLK), .D (IN_plaintext_s1[30]), .Q (new_AGEMA_signal_3548) ) ;
    buf_clk new_AGEMA_reg_buffer_2100 ( .C (CLK), .D (IN_plaintext_s0[31]), .Q (new_AGEMA_signal_3552) ) ;
    buf_clk new_AGEMA_reg_buffer_2104 ( .C (CLK), .D (IN_plaintext_s1[31]), .Q (new_AGEMA_signal_3556) ) ;
    buf_clk new_AGEMA_reg_buffer_2108 ( .C (CLK), .D (IN_plaintext_s0[32]), .Q (new_AGEMA_signal_3560) ) ;
    buf_clk new_AGEMA_reg_buffer_2112 ( .C (CLK), .D (IN_plaintext_s1[32]), .Q (new_AGEMA_signal_3564) ) ;
    buf_clk new_AGEMA_reg_buffer_2116 ( .C (CLK), .D (IN_plaintext_s0[33]), .Q (new_AGEMA_signal_3568) ) ;
    buf_clk new_AGEMA_reg_buffer_2120 ( .C (CLK), .D (IN_plaintext_s1[33]), .Q (new_AGEMA_signal_3572) ) ;
    buf_clk new_AGEMA_reg_buffer_2124 ( .C (CLK), .D (IN_plaintext_s0[34]), .Q (new_AGEMA_signal_3576) ) ;
    buf_clk new_AGEMA_reg_buffer_2128 ( .C (CLK), .D (IN_plaintext_s1[34]), .Q (new_AGEMA_signal_3580) ) ;
    buf_clk new_AGEMA_reg_buffer_2132 ( .C (CLK), .D (IN_plaintext_s0[35]), .Q (new_AGEMA_signal_3584) ) ;
    buf_clk new_AGEMA_reg_buffer_2136 ( .C (CLK), .D (IN_plaintext_s1[35]), .Q (new_AGEMA_signal_3588) ) ;
    buf_clk new_AGEMA_reg_buffer_2140 ( .C (CLK), .D (IN_plaintext_s0[36]), .Q (new_AGEMA_signal_3592) ) ;
    buf_clk new_AGEMA_reg_buffer_2144 ( .C (CLK), .D (IN_plaintext_s1[36]), .Q (new_AGEMA_signal_3596) ) ;
    buf_clk new_AGEMA_reg_buffer_2148 ( .C (CLK), .D (IN_plaintext_s0[37]), .Q (new_AGEMA_signal_3600) ) ;
    buf_clk new_AGEMA_reg_buffer_2152 ( .C (CLK), .D (IN_plaintext_s1[37]), .Q (new_AGEMA_signal_3604) ) ;
    buf_clk new_AGEMA_reg_buffer_2156 ( .C (CLK), .D (IN_plaintext_s0[38]), .Q (new_AGEMA_signal_3608) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (CLK), .D (IN_plaintext_s1[38]), .Q (new_AGEMA_signal_3612) ) ;
    buf_clk new_AGEMA_reg_buffer_2164 ( .C (CLK), .D (IN_plaintext_s0[39]), .Q (new_AGEMA_signal_3616) ) ;
    buf_clk new_AGEMA_reg_buffer_2168 ( .C (CLK), .D (IN_plaintext_s1[39]), .Q (new_AGEMA_signal_3620) ) ;
    buf_clk new_AGEMA_reg_buffer_2172 ( .C (CLK), .D (IN_plaintext_s0[40]), .Q (new_AGEMA_signal_3624) ) ;
    buf_clk new_AGEMA_reg_buffer_2176 ( .C (CLK), .D (IN_plaintext_s1[40]), .Q (new_AGEMA_signal_3628) ) ;
    buf_clk new_AGEMA_reg_buffer_2180 ( .C (CLK), .D (IN_plaintext_s0[41]), .Q (new_AGEMA_signal_3632) ) ;
    buf_clk new_AGEMA_reg_buffer_2184 ( .C (CLK), .D (IN_plaintext_s1[41]), .Q (new_AGEMA_signal_3636) ) ;
    buf_clk new_AGEMA_reg_buffer_2188 ( .C (CLK), .D (IN_plaintext_s0[42]), .Q (new_AGEMA_signal_3640) ) ;
    buf_clk new_AGEMA_reg_buffer_2192 ( .C (CLK), .D (IN_plaintext_s1[42]), .Q (new_AGEMA_signal_3644) ) ;
    buf_clk new_AGEMA_reg_buffer_2196 ( .C (CLK), .D (IN_plaintext_s0[43]), .Q (new_AGEMA_signal_3648) ) ;
    buf_clk new_AGEMA_reg_buffer_2200 ( .C (CLK), .D (IN_plaintext_s1[43]), .Q (new_AGEMA_signal_3652) ) ;
    buf_clk new_AGEMA_reg_buffer_2204 ( .C (CLK), .D (IN_plaintext_s0[44]), .Q (new_AGEMA_signal_3656) ) ;
    buf_clk new_AGEMA_reg_buffer_2208 ( .C (CLK), .D (IN_plaintext_s1[44]), .Q (new_AGEMA_signal_3660) ) ;
    buf_clk new_AGEMA_reg_buffer_2212 ( .C (CLK), .D (IN_plaintext_s0[45]), .Q (new_AGEMA_signal_3664) ) ;
    buf_clk new_AGEMA_reg_buffer_2216 ( .C (CLK), .D (IN_plaintext_s1[45]), .Q (new_AGEMA_signal_3668) ) ;
    buf_clk new_AGEMA_reg_buffer_2220 ( .C (CLK), .D (IN_plaintext_s0[46]), .Q (new_AGEMA_signal_3672) ) ;
    buf_clk new_AGEMA_reg_buffer_2224 ( .C (CLK), .D (IN_plaintext_s1[46]), .Q (new_AGEMA_signal_3676) ) ;
    buf_clk new_AGEMA_reg_buffer_2228 ( .C (CLK), .D (IN_plaintext_s0[47]), .Q (new_AGEMA_signal_3680) ) ;
    buf_clk new_AGEMA_reg_buffer_2232 ( .C (CLK), .D (IN_plaintext_s1[47]), .Q (new_AGEMA_signal_3684) ) ;
    buf_clk new_AGEMA_reg_buffer_2236 ( .C (CLK), .D (IN_plaintext_s0[48]), .Q (new_AGEMA_signal_3688) ) ;
    buf_clk new_AGEMA_reg_buffer_2240 ( .C (CLK), .D (IN_plaintext_s1[48]), .Q (new_AGEMA_signal_3692) ) ;
    buf_clk new_AGEMA_reg_buffer_2244 ( .C (CLK), .D (IN_plaintext_s0[49]), .Q (new_AGEMA_signal_3696) ) ;
    buf_clk new_AGEMA_reg_buffer_2248 ( .C (CLK), .D (IN_plaintext_s1[49]), .Q (new_AGEMA_signal_3700) ) ;
    buf_clk new_AGEMA_reg_buffer_2252 ( .C (CLK), .D (IN_plaintext_s0[50]), .Q (new_AGEMA_signal_3704) ) ;
    buf_clk new_AGEMA_reg_buffer_2256 ( .C (CLK), .D (IN_plaintext_s1[50]), .Q (new_AGEMA_signal_3708) ) ;
    buf_clk new_AGEMA_reg_buffer_2260 ( .C (CLK), .D (IN_plaintext_s0[51]), .Q (new_AGEMA_signal_3712) ) ;
    buf_clk new_AGEMA_reg_buffer_2264 ( .C (CLK), .D (IN_plaintext_s1[51]), .Q (new_AGEMA_signal_3716) ) ;
    buf_clk new_AGEMA_reg_buffer_2268 ( .C (CLK), .D (IN_plaintext_s0[52]), .Q (new_AGEMA_signal_3720) ) ;
    buf_clk new_AGEMA_reg_buffer_2272 ( .C (CLK), .D (IN_plaintext_s1[52]), .Q (new_AGEMA_signal_3724) ) ;
    buf_clk new_AGEMA_reg_buffer_2276 ( .C (CLK), .D (IN_plaintext_s0[53]), .Q (new_AGEMA_signal_3728) ) ;
    buf_clk new_AGEMA_reg_buffer_2280 ( .C (CLK), .D (IN_plaintext_s1[53]), .Q (new_AGEMA_signal_3732) ) ;
    buf_clk new_AGEMA_reg_buffer_2284 ( .C (CLK), .D (IN_plaintext_s0[54]), .Q (new_AGEMA_signal_3736) ) ;
    buf_clk new_AGEMA_reg_buffer_2288 ( .C (CLK), .D (IN_plaintext_s1[54]), .Q (new_AGEMA_signal_3740) ) ;
    buf_clk new_AGEMA_reg_buffer_2292 ( .C (CLK), .D (IN_plaintext_s0[55]), .Q (new_AGEMA_signal_3744) ) ;
    buf_clk new_AGEMA_reg_buffer_2296 ( .C (CLK), .D (IN_plaintext_s1[55]), .Q (new_AGEMA_signal_3748) ) ;
    buf_clk new_AGEMA_reg_buffer_2300 ( .C (CLK), .D (IN_plaintext_s0[56]), .Q (new_AGEMA_signal_3752) ) ;
    buf_clk new_AGEMA_reg_buffer_2304 ( .C (CLK), .D (IN_plaintext_s1[56]), .Q (new_AGEMA_signal_3756) ) ;
    buf_clk new_AGEMA_reg_buffer_2308 ( .C (CLK), .D (IN_plaintext_s0[57]), .Q (new_AGEMA_signal_3760) ) ;
    buf_clk new_AGEMA_reg_buffer_2312 ( .C (CLK), .D (IN_plaintext_s1[57]), .Q (new_AGEMA_signal_3764) ) ;
    buf_clk new_AGEMA_reg_buffer_2316 ( .C (CLK), .D (IN_plaintext_s0[58]), .Q (new_AGEMA_signal_3768) ) ;
    buf_clk new_AGEMA_reg_buffer_2320 ( .C (CLK), .D (IN_plaintext_s1[58]), .Q (new_AGEMA_signal_3772) ) ;
    buf_clk new_AGEMA_reg_buffer_2324 ( .C (CLK), .D (IN_plaintext_s0[59]), .Q (new_AGEMA_signal_3776) ) ;
    buf_clk new_AGEMA_reg_buffer_2328 ( .C (CLK), .D (IN_plaintext_s1[59]), .Q (new_AGEMA_signal_3780) ) ;
    buf_clk new_AGEMA_reg_buffer_2332 ( .C (CLK), .D (IN_plaintext_s0[60]), .Q (new_AGEMA_signal_3784) ) ;
    buf_clk new_AGEMA_reg_buffer_2336 ( .C (CLK), .D (IN_plaintext_s1[60]), .Q (new_AGEMA_signal_3788) ) ;
    buf_clk new_AGEMA_reg_buffer_2340 ( .C (CLK), .D (IN_plaintext_s0[61]), .Q (new_AGEMA_signal_3792) ) ;
    buf_clk new_AGEMA_reg_buffer_2344 ( .C (CLK), .D (IN_plaintext_s1[61]), .Q (new_AGEMA_signal_3796) ) ;
    buf_clk new_AGEMA_reg_buffer_2348 ( .C (CLK), .D (IN_plaintext_s0[62]), .Q (new_AGEMA_signal_3800) ) ;
    buf_clk new_AGEMA_reg_buffer_2352 ( .C (CLK), .D (IN_plaintext_s1[62]), .Q (new_AGEMA_signal_3804) ) ;
    buf_clk new_AGEMA_reg_buffer_2356 ( .C (CLK), .D (IN_plaintext_s0[63]), .Q (new_AGEMA_signal_3808) ) ;
    buf_clk new_AGEMA_reg_buffer_2360 ( .C (CLK), .D (IN_plaintext_s1[63]), .Q (new_AGEMA_signal_3812) ) ;
    buf_clk new_AGEMA_reg_buffer_2364 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_Q3), .Q (new_AGEMA_signal_3816) ) ;
    buf_clk new_AGEMA_reg_buffer_2366 ( .C (CLK), .D (new_AGEMA_signal_1878), .Q (new_AGEMA_signal_3818) ) ;
    buf_clk new_AGEMA_reg_buffer_2368 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_Q7), .Q (new_AGEMA_signal_3820) ) ;
    buf_clk new_AGEMA_reg_buffer_2370 ( .C (CLK), .D (new_AGEMA_signal_1879), .Q (new_AGEMA_signal_3822) ) ;
    buf_clk new_AGEMA_reg_buffer_2376 ( .C (CLK), .D (LED_128_Instance_addconst_out[0]), .Q (new_AGEMA_signal_3828) ) ;
    buf_clk new_AGEMA_reg_buffer_2380 ( .C (CLK), .D (new_AGEMA_signal_1665), .Q (new_AGEMA_signal_3832) ) ;
    buf_clk new_AGEMA_reg_buffer_2384 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L1), .Q (new_AGEMA_signal_3836) ) ;
    buf_clk new_AGEMA_reg_buffer_2388 ( .C (CLK), .D (new_AGEMA_signal_1801), .Q (new_AGEMA_signal_3840) ) ;
    buf_clk new_AGEMA_reg_buffer_2396 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_Q3), .Q (new_AGEMA_signal_3848) ) ;
    buf_clk new_AGEMA_reg_buffer_2398 ( .C (CLK), .D (new_AGEMA_signal_1883), .Q (new_AGEMA_signal_3850) ) ;
    buf_clk new_AGEMA_reg_buffer_2400 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_Q7), .Q (new_AGEMA_signal_3852) ) ;
    buf_clk new_AGEMA_reg_buffer_2402 ( .C (CLK), .D (new_AGEMA_signal_1884), .Q (new_AGEMA_signal_3854) ) ;
    buf_clk new_AGEMA_reg_buffer_2408 ( .C (CLK), .D (LED_128_Instance_addconst_out[4]), .Q (new_AGEMA_signal_3860) ) ;
    buf_clk new_AGEMA_reg_buffer_2412 ( .C (CLK), .D (new_AGEMA_signal_1733), .Q (new_AGEMA_signal_3864) ) ;
    buf_clk new_AGEMA_reg_buffer_2416 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L1), .Q (new_AGEMA_signal_3868) ) ;
    buf_clk new_AGEMA_reg_buffer_2420 ( .C (CLK), .D (new_AGEMA_signal_1805), .Q (new_AGEMA_signal_3872) ) ;
    buf_clk new_AGEMA_reg_buffer_2428 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_Q3), .Q (new_AGEMA_signal_3880) ) ;
    buf_clk new_AGEMA_reg_buffer_2430 ( .C (CLK), .D (new_AGEMA_signal_1810), .Q (new_AGEMA_signal_3882) ) ;
    buf_clk new_AGEMA_reg_buffer_2432 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_Q7), .Q (new_AGEMA_signal_3884) ) ;
    buf_clk new_AGEMA_reg_buffer_2434 ( .C (CLK), .D (new_AGEMA_signal_1811), .Q (new_AGEMA_signal_3886) ) ;
    buf_clk new_AGEMA_reg_buffer_2440 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L1), .Q (new_AGEMA_signal_3892) ) ;
    buf_clk new_AGEMA_reg_buffer_2444 ( .C (CLK), .D (new_AGEMA_signal_1749), .Q (new_AGEMA_signal_3896) ) ;
    buf_clk new_AGEMA_reg_buffer_2452 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_Q3), .Q (new_AGEMA_signal_3904) ) ;
    buf_clk new_AGEMA_reg_buffer_2454 ( .C (CLK), .D (new_AGEMA_signal_1815), .Q (new_AGEMA_signal_3906) ) ;
    buf_clk new_AGEMA_reg_buffer_2456 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_Q7), .Q (new_AGEMA_signal_3908) ) ;
    buf_clk new_AGEMA_reg_buffer_2458 ( .C (CLK), .D (new_AGEMA_signal_1816), .Q (new_AGEMA_signal_3910) ) ;
    buf_clk new_AGEMA_reg_buffer_2464 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L1), .Q (new_AGEMA_signal_3916) ) ;
    buf_clk new_AGEMA_reg_buffer_2468 ( .C (CLK), .D (new_AGEMA_signal_1755), .Q (new_AGEMA_signal_3920) ) ;
    buf_clk new_AGEMA_reg_buffer_2476 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_Q3), .Q (new_AGEMA_signal_3928) ) ;
    buf_clk new_AGEMA_reg_buffer_2478 ( .C (CLK), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_3930) ) ;
    buf_clk new_AGEMA_reg_buffer_2480 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_Q7), .Q (new_AGEMA_signal_3932) ) ;
    buf_clk new_AGEMA_reg_buffer_2482 ( .C (CLK), .D (new_AGEMA_signal_1893), .Q (new_AGEMA_signal_3934) ) ;
    buf_clk new_AGEMA_reg_buffer_2488 ( .C (CLK), .D (LED_128_Instance_addconst_out[16]), .Q (new_AGEMA_signal_3940) ) ;
    buf_clk new_AGEMA_reg_buffer_2492 ( .C (CLK), .D (new_AGEMA_signal_1664), .Q (new_AGEMA_signal_3944) ) ;
    buf_clk new_AGEMA_reg_buffer_2496 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L1), .Q (new_AGEMA_signal_3948) ) ;
    buf_clk new_AGEMA_reg_buffer_2500 ( .C (CLK), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_3952) ) ;
    buf_clk new_AGEMA_reg_buffer_2508 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_Q3), .Q (new_AGEMA_signal_3960) ) ;
    buf_clk new_AGEMA_reg_buffer_2510 ( .C (CLK), .D (new_AGEMA_signal_1897), .Q (new_AGEMA_signal_3962) ) ;
    buf_clk new_AGEMA_reg_buffer_2512 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_Q7), .Q (new_AGEMA_signal_3964) ) ;
    buf_clk new_AGEMA_reg_buffer_2514 ( .C (CLK), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_3966) ) ;
    buf_clk new_AGEMA_reg_buffer_2520 ( .C (CLK), .D (LED_128_Instance_addconst_out[20]), .Q (new_AGEMA_signal_3972) ) ;
    buf_clk new_AGEMA_reg_buffer_2524 ( .C (CLK), .D (new_AGEMA_signal_1741), .Q (new_AGEMA_signal_3976) ) ;
    buf_clk new_AGEMA_reg_buffer_2528 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L1), .Q (new_AGEMA_signal_3980) ) ;
    buf_clk new_AGEMA_reg_buffer_2532 ( .C (CLK), .D (new_AGEMA_signal_1824), .Q (new_AGEMA_signal_3984) ) ;
    buf_clk new_AGEMA_reg_buffer_2540 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_Q3), .Q (new_AGEMA_signal_3992) ) ;
    buf_clk new_AGEMA_reg_buffer_2542 ( .C (CLK), .D (new_AGEMA_signal_1829), .Q (new_AGEMA_signal_3994) ) ;
    buf_clk new_AGEMA_reg_buffer_2544 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_Q7), .Q (new_AGEMA_signal_3996) ) ;
    buf_clk new_AGEMA_reg_buffer_2546 ( .C (CLK), .D (new_AGEMA_signal_1830), .Q (new_AGEMA_signal_3998) ) ;
    buf_clk new_AGEMA_reg_buffer_2552 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L1), .Q (new_AGEMA_signal_4004) ) ;
    buf_clk new_AGEMA_reg_buffer_2556 ( .C (CLK), .D (new_AGEMA_signal_1762), .Q (new_AGEMA_signal_4008) ) ;
    buf_clk new_AGEMA_reg_buffer_2564 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_Q3), .Q (new_AGEMA_signal_4016) ) ;
    buf_clk new_AGEMA_reg_buffer_2566 ( .C (CLK), .D (new_AGEMA_signal_1834), .Q (new_AGEMA_signal_4018) ) ;
    buf_clk new_AGEMA_reg_buffer_2568 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_Q7), .Q (new_AGEMA_signal_4020) ) ;
    buf_clk new_AGEMA_reg_buffer_2570 ( .C (CLK), .D (new_AGEMA_signal_1835), .Q (new_AGEMA_signal_4022) ) ;
    buf_clk new_AGEMA_reg_buffer_2576 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L1), .Q (new_AGEMA_signal_4028) ) ;
    buf_clk new_AGEMA_reg_buffer_2580 ( .C (CLK), .D (new_AGEMA_signal_1768), .Q (new_AGEMA_signal_4032) ) ;
    buf_clk new_AGEMA_reg_buffer_2588 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_Q3), .Q (new_AGEMA_signal_4040) ) ;
    buf_clk new_AGEMA_reg_buffer_2590 ( .C (CLK), .D (new_AGEMA_signal_1906), .Q (new_AGEMA_signal_4042) ) ;
    buf_clk new_AGEMA_reg_buffer_2592 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_Q7), .Q (new_AGEMA_signal_4044) ) ;
    buf_clk new_AGEMA_reg_buffer_2594 ( .C (CLK), .D (new_AGEMA_signal_1907), .Q (new_AGEMA_signal_4046) ) ;
    buf_clk new_AGEMA_reg_buffer_2600 ( .C (CLK), .D (LED_128_Instance_addconst_out[32]), .Q (new_AGEMA_signal_4052) ) ;
    buf_clk new_AGEMA_reg_buffer_2604 ( .C (CLK), .D (new_AGEMA_signal_1720), .Q (new_AGEMA_signal_4056) ) ;
    buf_clk new_AGEMA_reg_buffer_2608 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L1), .Q (new_AGEMA_signal_4060) ) ;
    buf_clk new_AGEMA_reg_buffer_2612 ( .C (CLK), .D (new_AGEMA_signal_1839), .Q (new_AGEMA_signal_4064) ) ;
    buf_clk new_AGEMA_reg_buffer_2620 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_Q3), .Q (new_AGEMA_signal_4072) ) ;
    buf_clk new_AGEMA_reg_buffer_2622 ( .C (CLK), .D (new_AGEMA_signal_1911), .Q (new_AGEMA_signal_4074) ) ;
    buf_clk new_AGEMA_reg_buffer_2624 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_Q7), .Q (new_AGEMA_signal_4076) ) ;
    buf_clk new_AGEMA_reg_buffer_2626 ( .C (CLK), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_4078) ) ;
    buf_clk new_AGEMA_reg_buffer_2632 ( .C (CLK), .D (LED_128_Instance_addconst_out[36]), .Q (new_AGEMA_signal_4084) ) ;
    buf_clk new_AGEMA_reg_buffer_2636 ( .C (CLK), .D (new_AGEMA_signal_1717), .Q (new_AGEMA_signal_4088) ) ;
    buf_clk new_AGEMA_reg_buffer_2640 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L1), .Q (new_AGEMA_signal_4092) ) ;
    buf_clk new_AGEMA_reg_buffer_2644 ( .C (CLK), .D (new_AGEMA_signal_1843), .Q (new_AGEMA_signal_4096) ) ;
    buf_clk new_AGEMA_reg_buffer_2652 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_Q3), .Q (new_AGEMA_signal_4104) ) ;
    buf_clk new_AGEMA_reg_buffer_2654 ( .C (CLK), .D (new_AGEMA_signal_1847), .Q (new_AGEMA_signal_4106) ) ;
    buf_clk new_AGEMA_reg_buffer_2656 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_Q7), .Q (new_AGEMA_signal_4108) ) ;
    buf_clk new_AGEMA_reg_buffer_2658 ( .C (CLK), .D (new_AGEMA_signal_1848), .Q (new_AGEMA_signal_4110) ) ;
    buf_clk new_AGEMA_reg_buffer_2664 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L1), .Q (new_AGEMA_signal_4116) ) ;
    buf_clk new_AGEMA_reg_buffer_2668 ( .C (CLK), .D (new_AGEMA_signal_1777), .Q (new_AGEMA_signal_4120) ) ;
    buf_clk new_AGEMA_reg_buffer_2676 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_Q3), .Q (new_AGEMA_signal_4128) ) ;
    buf_clk new_AGEMA_reg_buffer_2678 ( .C (CLK), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_4130) ) ;
    buf_clk new_AGEMA_reg_buffer_2680 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_Q7), .Q (new_AGEMA_signal_4132) ) ;
    buf_clk new_AGEMA_reg_buffer_2682 ( .C (CLK), .D (new_AGEMA_signal_1853), .Q (new_AGEMA_signal_4134) ) ;
    buf_clk new_AGEMA_reg_buffer_2688 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L1), .Q (new_AGEMA_signal_4140) ) ;
    buf_clk new_AGEMA_reg_buffer_2692 ( .C (CLK), .D (new_AGEMA_signal_1783), .Q (new_AGEMA_signal_4144) ) ;
    buf_clk new_AGEMA_reg_buffer_2700 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_Q3), .Q (new_AGEMA_signal_4152) ) ;
    buf_clk new_AGEMA_reg_buffer_2702 ( .C (CLK), .D (new_AGEMA_signal_1920), .Q (new_AGEMA_signal_4154) ) ;
    buf_clk new_AGEMA_reg_buffer_2704 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_Q7), .Q (new_AGEMA_signal_4156) ) ;
    buf_clk new_AGEMA_reg_buffer_2706 ( .C (CLK), .D (new_AGEMA_signal_1921), .Q (new_AGEMA_signal_4158) ) ;
    buf_clk new_AGEMA_reg_buffer_2712 ( .C (CLK), .D (LED_128_Instance_addconst_out[48]), .Q (new_AGEMA_signal_4164) ) ;
    buf_clk new_AGEMA_reg_buffer_2716 ( .C (CLK), .D (new_AGEMA_signal_1735), .Q (new_AGEMA_signal_4168) ) ;
    buf_clk new_AGEMA_reg_buffer_2720 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L1), .Q (new_AGEMA_signal_4172) ) ;
    buf_clk new_AGEMA_reg_buffer_2724 ( .C (CLK), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_4176) ) ;
    buf_clk new_AGEMA_reg_buffer_2732 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_Q3), .Q (new_AGEMA_signal_4184) ) ;
    buf_clk new_AGEMA_reg_buffer_2734 ( .C (CLK), .D (new_AGEMA_signal_1925), .Q (new_AGEMA_signal_4186) ) ;
    buf_clk new_AGEMA_reg_buffer_2736 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_Q7), .Q (new_AGEMA_signal_4188) ) ;
    buf_clk new_AGEMA_reg_buffer_2738 ( .C (CLK), .D (new_AGEMA_signal_1926), .Q (new_AGEMA_signal_4190) ) ;
    buf_clk new_AGEMA_reg_buffer_2744 ( .C (CLK), .D (LED_128_Instance_addconst_out[52]), .Q (new_AGEMA_signal_4196) ) ;
    buf_clk new_AGEMA_reg_buffer_2748 ( .C (CLK), .D (new_AGEMA_signal_1730), .Q (new_AGEMA_signal_4200) ) ;
    buf_clk new_AGEMA_reg_buffer_2752 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L1), .Q (new_AGEMA_signal_4204) ) ;
    buf_clk new_AGEMA_reg_buffer_2756 ( .C (CLK), .D (new_AGEMA_signal_1863), .Q (new_AGEMA_signal_4208) ) ;
    buf_clk new_AGEMA_reg_buffer_2764 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_Q3), .Q (new_AGEMA_signal_4216) ) ;
    buf_clk new_AGEMA_reg_buffer_2766 ( .C (CLK), .D (new_AGEMA_signal_1868), .Q (new_AGEMA_signal_4218) ) ;
    buf_clk new_AGEMA_reg_buffer_2768 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_Q7), .Q (new_AGEMA_signal_4220) ) ;
    buf_clk new_AGEMA_reg_buffer_2770 ( .C (CLK), .D (new_AGEMA_signal_1869), .Q (new_AGEMA_signal_4222) ) ;
    buf_clk new_AGEMA_reg_buffer_2776 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L1), .Q (new_AGEMA_signal_4228) ) ;
    buf_clk new_AGEMA_reg_buffer_2780 ( .C (CLK), .D (new_AGEMA_signal_1790), .Q (new_AGEMA_signal_4232) ) ;
    buf_clk new_AGEMA_reg_buffer_2788 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_Q3), .Q (new_AGEMA_signal_4240) ) ;
    buf_clk new_AGEMA_reg_buffer_2790 ( .C (CLK), .D (new_AGEMA_signal_1873), .Q (new_AGEMA_signal_4242) ) ;
    buf_clk new_AGEMA_reg_buffer_2792 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_Q7), .Q (new_AGEMA_signal_4244) ) ;
    buf_clk new_AGEMA_reg_buffer_2794 ( .C (CLK), .D (new_AGEMA_signal_1874), .Q (new_AGEMA_signal_4246) ) ;
    buf_clk new_AGEMA_reg_buffer_2800 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L1), .Q (new_AGEMA_signal_4252) ) ;
    buf_clk new_AGEMA_reg_buffer_2804 ( .C (CLK), .D (new_AGEMA_signal_1796), .Q (new_AGEMA_signal_4256) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (CLK), .D (LED_128_Instance_N10), .Q (new_AGEMA_signal_4328) ) ;
    buf_clk new_AGEMA_reg_buffer_2880 ( .C (CLK), .D (LED_128_Instance_N11), .Q (new_AGEMA_signal_4332) ) ;
    buf_clk new_AGEMA_reg_buffer_2884 ( .C (CLK), .D (LED_128_Instance_N12), .Q (new_AGEMA_signal_4336) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (CLK), .D (LED_128_Instance_N13), .Q (new_AGEMA_signal_4340) ) ;
    buf_clk new_AGEMA_reg_buffer_2892 ( .C (CLK), .D (LED_128_Instance_N4), .Q (new_AGEMA_signal_4344) ) ;
    buf_clk new_AGEMA_reg_buffer_2896 ( .C (CLK), .D (LED_128_Instance_N5), .Q (new_AGEMA_signal_4348) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (CLK), .D (LED_128_Instance_N6), .Q (new_AGEMA_signal_4352) ) ;
    buf_clk new_AGEMA_reg_buffer_2904 ( .C (CLK), .D (LED_128_Instance_N7), .Q (new_AGEMA_signal_4356) ) ;
    buf_clk new_AGEMA_reg_buffer_2908 ( .C (CLK), .D (LED_128_Instance_N8), .Q (new_AGEMA_signal_4360) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (CLK), .D (LED_128_Instance_N9), .Q (new_AGEMA_signal_4364) ) ;
    buf_clk new_AGEMA_reg_buffer_2916 ( .C (CLK), .D (n15), .Q (new_AGEMA_signal_4368) ) ;

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR16_U1 ( .a ({new_AGEMA_signal_1932, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_2583, new_AGEMA_signal_2581}), .c ({new_AGEMA_signal_1964, LED_128_Instance_SBox_Instance_0_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR7_U1 ( .a ({new_AGEMA_signal_1932, LED_128_Instance_SBox_Instance_0_T0}), .b ({new_AGEMA_signal_1880, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_1965, LED_128_Instance_SBox_Instance_0_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR8_U1 ( .a ({new_AGEMA_signal_2587, new_AGEMA_signal_2585}), .b ({new_AGEMA_signal_1965, LED_128_Instance_SBox_Instance_0_L5}), .c ({new_AGEMA_signal_1996, LED_128_Instance_SBox_Instance_0_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND1_U1 ( .a ({new_AGEMA_signal_1876, LED_128_Instance_SBox_Instance_0_n1}), .b ({new_AGEMA_signal_1721, LED_128_Instance_SBox_Instance_0_n2}), .clk (CLK), .r (Fresh[0]), .c ({new_AGEMA_signal_1932, LED_128_Instance_SBox_Instance_0_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND3_U1 ( .a ({new_AGEMA_signal_1799, LED_128_Instance_SBox_Instance_0_n3}), .b ({new_AGEMA_signal_1739, LED_128_Instance_addconst_out[2]}), .clk (CLK), .r (Fresh[1]), .c ({new_AGEMA_signal_1880, LED_128_Instance_SBox_Instance_0_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR15_U1 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2589}), .b ({new_AGEMA_signal_1880, LED_128_Instance_SBox_Instance_0_T2}), .c ({new_AGEMA_signal_1933, LED_128_Instance_subcells_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR16_U1 ( .a ({new_AGEMA_signal_1934, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2593}), .c ({new_AGEMA_signal_1966, LED_128_Instance_SBox_Instance_1_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR7_U1 ( .a ({new_AGEMA_signal_1934, LED_128_Instance_SBox_Instance_1_T0}), .b ({new_AGEMA_signal_1885, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_1967, LED_128_Instance_SBox_Instance_1_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR8_U1 ( .a ({new_AGEMA_signal_2599, new_AGEMA_signal_2597}), .b ({new_AGEMA_signal_1967, LED_128_Instance_SBox_Instance_1_L5}), .c ({new_AGEMA_signal_1998, LED_128_Instance_SBox_Instance_1_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND1_U1 ( .a ({new_AGEMA_signal_1881, LED_128_Instance_SBox_Instance_1_n1}), .b ({new_AGEMA_signal_1745, LED_128_Instance_SBox_Instance_1_n2}), .clk (CLK), .r (Fresh[2]), .c ({new_AGEMA_signal_1934, LED_128_Instance_SBox_Instance_1_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND3_U1 ( .a ({new_AGEMA_signal_1803, LED_128_Instance_SBox_Instance_1_n3}), .b ({new_AGEMA_signal_1726, LED_128_Instance_addconst_out[6]}), .clk (CLK), .r (Fresh[3]), .c ({new_AGEMA_signal_1885, LED_128_Instance_SBox_Instance_1_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR15_U1 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2601}), .b ({new_AGEMA_signal_1885, LED_128_Instance_SBox_Instance_1_T2}), .c ({new_AGEMA_signal_1935, LED_128_Instance_subcells_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR16_U1 ( .a ({new_AGEMA_signal_1886, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_2607, new_AGEMA_signal_2605}), .c ({new_AGEMA_signal_1936, LED_128_Instance_SBox_Instance_2_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR7_U1 ( .a ({new_AGEMA_signal_1886, LED_128_Instance_SBox_Instance_2_T0}), .b ({new_AGEMA_signal_1812, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_1937, LED_128_Instance_SBox_Instance_2_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR8_U1 ( .a ({new_AGEMA_signal_2611, new_AGEMA_signal_2609}), .b ({new_AGEMA_signal_1937, LED_128_Instance_SBox_Instance_2_L5}), .c ({new_AGEMA_signal_1968, LED_128_Instance_SBox_Instance_2_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND1_U1 ( .a ({new_AGEMA_signal_1808, LED_128_Instance_SBox_Instance_2_n1}), .b ({new_AGEMA_signal_1746, LED_128_Instance_SBox_Instance_2_n2}), .clk (CLK), .r (Fresh[4]), .c ({new_AGEMA_signal_1886, LED_128_Instance_SBox_Instance_2_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND3_U1 ( .a ({new_AGEMA_signal_1747, LED_128_Instance_SBox_Instance_2_n3}), .b ({new_AGEMA_signal_1674, LED_128_Instance_addconst_out[10]}), .clk (CLK), .r (Fresh[5]), .c ({new_AGEMA_signal_1812, LED_128_Instance_SBox_Instance_2_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR15_U1 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2613}), .b ({new_AGEMA_signal_1812, LED_128_Instance_SBox_Instance_2_T2}), .c ({new_AGEMA_signal_1887, LED_128_Instance_subcells_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR16_U1 ( .a ({new_AGEMA_signal_1888, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_2619, new_AGEMA_signal_2617}), .c ({new_AGEMA_signal_1938, LED_128_Instance_SBox_Instance_3_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR7_U1 ( .a ({new_AGEMA_signal_1888, LED_128_Instance_SBox_Instance_3_T0}), .b ({new_AGEMA_signal_1817, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_1939, LED_128_Instance_SBox_Instance_3_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR8_U1 ( .a ({new_AGEMA_signal_2623, new_AGEMA_signal_2621}), .b ({new_AGEMA_signal_1939, LED_128_Instance_SBox_Instance_3_L5}), .c ({new_AGEMA_signal_1970, LED_128_Instance_SBox_Instance_3_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND1_U1 ( .a ({new_AGEMA_signal_1813, LED_128_Instance_SBox_Instance_3_n1}), .b ({new_AGEMA_signal_1752, LED_128_Instance_SBox_Instance_3_n2}), .clk (CLK), .r (Fresh[6]), .c ({new_AGEMA_signal_1888, LED_128_Instance_SBox_Instance_3_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND3_U1 ( .a ({new_AGEMA_signal_1753, LED_128_Instance_SBox_Instance_3_n3}), .b ({new_AGEMA_signal_1678, LED_128_Instance_addconst_out[14]}), .clk (CLK), .r (Fresh[7]), .c ({new_AGEMA_signal_1817, LED_128_Instance_SBox_Instance_3_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR15_U1 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2625}), .b ({new_AGEMA_signal_1817, LED_128_Instance_SBox_Instance_3_T2}), .c ({new_AGEMA_signal_1889, LED_128_Instance_subcells_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR16_U1 ( .a ({new_AGEMA_signal_1940, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_2631, new_AGEMA_signal_2629}), .c ({new_AGEMA_signal_1972, LED_128_Instance_SBox_Instance_4_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR7_U1 ( .a ({new_AGEMA_signal_1940, LED_128_Instance_SBox_Instance_4_T0}), .b ({new_AGEMA_signal_1894, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_1973, LED_128_Instance_SBox_Instance_4_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR8_U1 ( .a ({new_AGEMA_signal_2635, new_AGEMA_signal_2633}), .b ({new_AGEMA_signal_1973, LED_128_Instance_SBox_Instance_4_L5}), .c ({new_AGEMA_signal_2004, LED_128_Instance_SBox_Instance_4_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND1_U1 ( .a ({new_AGEMA_signal_1890, LED_128_Instance_SBox_Instance_4_n1}), .b ({new_AGEMA_signal_1723, LED_128_Instance_SBox_Instance_4_n2}), .clk (CLK), .r (Fresh[8]), .c ({new_AGEMA_signal_1940, LED_128_Instance_SBox_Instance_4_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND3_U1 ( .a ({new_AGEMA_signal_1818, LED_128_Instance_SBox_Instance_4_n3}), .b ({new_AGEMA_signal_1743, LED_128_Instance_addconst_out[18]}), .clk (CLK), .r (Fresh[9]), .c ({new_AGEMA_signal_1894, LED_128_Instance_SBox_Instance_4_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR15_U1 ( .a ({new_AGEMA_signal_2639, new_AGEMA_signal_2637}), .b ({new_AGEMA_signal_1894, LED_128_Instance_SBox_Instance_4_T2}), .c ({new_AGEMA_signal_1941, LED_128_Instance_subcells_out[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR16_U1 ( .a ({new_AGEMA_signal_1942, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_2643, new_AGEMA_signal_2641}), .c ({new_AGEMA_signal_1974, LED_128_Instance_SBox_Instance_5_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR7_U1 ( .a ({new_AGEMA_signal_1942, LED_128_Instance_SBox_Instance_5_T0}), .b ({new_AGEMA_signal_1899, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_1975, LED_128_Instance_SBox_Instance_5_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR8_U1 ( .a ({new_AGEMA_signal_2647, new_AGEMA_signal_2645}), .b ({new_AGEMA_signal_1975, LED_128_Instance_SBox_Instance_5_L5}), .c ({new_AGEMA_signal_2006, LED_128_Instance_SBox_Instance_5_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND1_U1 ( .a ({new_AGEMA_signal_1895, LED_128_Instance_SBox_Instance_5_n1}), .b ({new_AGEMA_signal_1758, LED_128_Instance_SBox_Instance_5_n2}), .clk (CLK), .r (Fresh[10]), .c ({new_AGEMA_signal_1942, LED_128_Instance_SBox_Instance_5_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND3_U1 ( .a ({new_AGEMA_signal_1822, LED_128_Instance_SBox_Instance_5_n3}), .b ({new_AGEMA_signal_1662, LED_128_Instance_addconst_out[22]}), .clk (CLK), .r (Fresh[11]), .c ({new_AGEMA_signal_1899, LED_128_Instance_SBox_Instance_5_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR15_U1 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2649}), .b ({new_AGEMA_signal_1899, LED_128_Instance_SBox_Instance_5_T2}), .c ({new_AGEMA_signal_1943, LED_128_Instance_subcells_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR16_U1 ( .a ({new_AGEMA_signal_1900, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_2655, new_AGEMA_signal_2653}), .c ({new_AGEMA_signal_1944, LED_128_Instance_SBox_Instance_6_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR7_U1 ( .a ({new_AGEMA_signal_1900, LED_128_Instance_SBox_Instance_6_T0}), .b ({new_AGEMA_signal_1831, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_1945, LED_128_Instance_SBox_Instance_6_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR8_U1 ( .a ({new_AGEMA_signal_2659, new_AGEMA_signal_2657}), .b ({new_AGEMA_signal_1945, LED_128_Instance_SBox_Instance_6_L5}), .c ({new_AGEMA_signal_1976, LED_128_Instance_SBox_Instance_6_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND1_U1 ( .a ({new_AGEMA_signal_1827, LED_128_Instance_SBox_Instance_6_n1}), .b ({new_AGEMA_signal_1759, LED_128_Instance_SBox_Instance_6_n2}), .clk (CLK), .r (Fresh[12]), .c ({new_AGEMA_signal_1900, LED_128_Instance_SBox_Instance_6_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND3_U1 ( .a ({new_AGEMA_signal_1760, LED_128_Instance_SBox_Instance_6_n3}), .b ({new_AGEMA_signal_1552, LED_128_Instance_addconst_out[26]}), .clk (CLK), .r (Fresh[13]), .c ({new_AGEMA_signal_1831, LED_128_Instance_SBox_Instance_6_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR15_U1 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2661}), .b ({new_AGEMA_signal_1831, LED_128_Instance_SBox_Instance_6_T2}), .c ({new_AGEMA_signal_1901, LED_128_Instance_subcells_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR16_U1 ( .a ({new_AGEMA_signal_1902, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_2667, new_AGEMA_signal_2665}), .c ({new_AGEMA_signal_1946, LED_128_Instance_SBox_Instance_7_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR7_U1 ( .a ({new_AGEMA_signal_1902, LED_128_Instance_SBox_Instance_7_T0}), .b ({new_AGEMA_signal_1836, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_1947, LED_128_Instance_SBox_Instance_7_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR8_U1 ( .a ({new_AGEMA_signal_2671, new_AGEMA_signal_2669}), .b ({new_AGEMA_signal_1947, LED_128_Instance_SBox_Instance_7_L5}), .c ({new_AGEMA_signal_1978, LED_128_Instance_SBox_Instance_7_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND1_U1 ( .a ({new_AGEMA_signal_1832, LED_128_Instance_SBox_Instance_7_n1}), .b ({new_AGEMA_signal_1765, LED_128_Instance_SBox_Instance_7_n2}), .clk (CLK), .r (Fresh[14]), .c ({new_AGEMA_signal_1902, LED_128_Instance_SBox_Instance_7_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND3_U1 ( .a ({new_AGEMA_signal_1766, LED_128_Instance_SBox_Instance_7_n3}), .b ({new_AGEMA_signal_1688, LED_128_Instance_addconst_out[30]}), .clk (CLK), .r (Fresh[15]), .c ({new_AGEMA_signal_1836, LED_128_Instance_SBox_Instance_7_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR15_U1 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2673}), .b ({new_AGEMA_signal_1836, LED_128_Instance_SBox_Instance_7_T2}), .c ({new_AGEMA_signal_1903, LED_128_Instance_subcells_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR16_U1 ( .a ({new_AGEMA_signal_1948, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_2679, new_AGEMA_signal_2677}), .c ({new_AGEMA_signal_1980, LED_128_Instance_SBox_Instance_8_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR7_U1 ( .a ({new_AGEMA_signal_1948, LED_128_Instance_SBox_Instance_8_T0}), .b ({new_AGEMA_signal_1908, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_1981, LED_128_Instance_SBox_Instance_8_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR8_U1 ( .a ({new_AGEMA_signal_2683, new_AGEMA_signal_2681}), .b ({new_AGEMA_signal_1981, LED_128_Instance_SBox_Instance_8_L5}), .c ({new_AGEMA_signal_2012, LED_128_Instance_SBox_Instance_8_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND1_U1 ( .a ({new_AGEMA_signal_1904, LED_128_Instance_SBox_Instance_8_n1}), .b ({new_AGEMA_signal_1771, LED_128_Instance_SBox_Instance_8_n2}), .clk (CLK), .r (Fresh[16]), .c ({new_AGEMA_signal_1948, LED_128_Instance_SBox_Instance_8_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND3_U1 ( .a ({new_AGEMA_signal_1837, LED_128_Instance_SBox_Instance_8_n3}), .b ({new_AGEMA_signal_1719, LED_128_Instance_addconst_out[34]}), .clk (CLK), .r (Fresh[17]), .c ({new_AGEMA_signal_1908, LED_128_Instance_SBox_Instance_8_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR15_U1 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2685}), .b ({new_AGEMA_signal_1908, LED_128_Instance_SBox_Instance_8_T2}), .c ({new_AGEMA_signal_1949, LED_128_Instance_subcells_out[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR16_U1 ( .a ({new_AGEMA_signal_1950, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_2691, new_AGEMA_signal_2689}), .c ({new_AGEMA_signal_1982, LED_128_Instance_SBox_Instance_9_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR7_U1 ( .a ({new_AGEMA_signal_1950, LED_128_Instance_SBox_Instance_9_T0}), .b ({new_AGEMA_signal_1913, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_1983, LED_128_Instance_SBox_Instance_9_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR8_U1 ( .a ({new_AGEMA_signal_2695, new_AGEMA_signal_2693}), .b ({new_AGEMA_signal_1983, LED_128_Instance_SBox_Instance_9_L5}), .c ({new_AGEMA_signal_2014, LED_128_Instance_SBox_Instance_9_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND1_U1 ( .a ({new_AGEMA_signal_1909, LED_128_Instance_SBox_Instance_9_n1}), .b ({new_AGEMA_signal_1725, LED_128_Instance_SBox_Instance_9_n2}), .clk (CLK), .r (Fresh[18]), .c ({new_AGEMA_signal_1950, LED_128_Instance_SBox_Instance_9_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND3_U1 ( .a ({new_AGEMA_signal_1841, LED_128_Instance_SBox_Instance_9_n3}), .b ({new_AGEMA_signal_1736, LED_128_Instance_addconst_out[38]}), .clk (CLK), .r (Fresh[19]), .c ({new_AGEMA_signal_1913, LED_128_Instance_SBox_Instance_9_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR15_U1 ( .a ({new_AGEMA_signal_2699, new_AGEMA_signal_2697}), .b ({new_AGEMA_signal_1913, LED_128_Instance_SBox_Instance_9_T2}), .c ({new_AGEMA_signal_1951, LED_128_Instance_subcells_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR16_U1 ( .a ({new_AGEMA_signal_1914, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_2703, new_AGEMA_signal_2701}), .c ({new_AGEMA_signal_1952, LED_128_Instance_SBox_Instance_10_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR7_U1 ( .a ({new_AGEMA_signal_1914, LED_128_Instance_SBox_Instance_10_T0}), .b ({new_AGEMA_signal_1849, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_1953, LED_128_Instance_SBox_Instance_10_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR8_U1 ( .a ({new_AGEMA_signal_2707, new_AGEMA_signal_2705}), .b ({new_AGEMA_signal_1953, LED_128_Instance_SBox_Instance_10_L5}), .c ({new_AGEMA_signal_1984, LED_128_Instance_SBox_Instance_10_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND1_U1 ( .a ({new_AGEMA_signal_1845, LED_128_Instance_SBox_Instance_10_n1}), .b ({new_AGEMA_signal_1774, LED_128_Instance_SBox_Instance_10_n2}), .clk (CLK), .r (Fresh[20]), .c ({new_AGEMA_signal_1914, LED_128_Instance_SBox_Instance_10_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND3_U1 ( .a ({new_AGEMA_signal_1775, LED_128_Instance_SBox_Instance_10_n3}), .b ({new_AGEMA_signal_1695, LED_128_Instance_addconst_out[42]}), .clk (CLK), .r (Fresh[21]), .c ({new_AGEMA_signal_1849, LED_128_Instance_SBox_Instance_10_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR15_U1 ( .a ({new_AGEMA_signal_2711, new_AGEMA_signal_2709}), .b ({new_AGEMA_signal_1849, LED_128_Instance_SBox_Instance_10_T2}), .c ({new_AGEMA_signal_1915, LED_128_Instance_subcells_out[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR16_U1 ( .a ({new_AGEMA_signal_1916, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_2715, new_AGEMA_signal_2713}), .c ({new_AGEMA_signal_1954, LED_128_Instance_SBox_Instance_11_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR7_U1 ( .a ({new_AGEMA_signal_1916, LED_128_Instance_SBox_Instance_11_T0}), .b ({new_AGEMA_signal_1854, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_1955, LED_128_Instance_SBox_Instance_11_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR8_U1 ( .a ({new_AGEMA_signal_2719, new_AGEMA_signal_2717}), .b ({new_AGEMA_signal_1955, LED_128_Instance_SBox_Instance_11_L5}), .c ({new_AGEMA_signal_1986, LED_128_Instance_SBox_Instance_11_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND1_U1 ( .a ({new_AGEMA_signal_1850, LED_128_Instance_SBox_Instance_11_n1}), .b ({new_AGEMA_signal_1780, LED_128_Instance_SBox_Instance_11_n2}), .clk (CLK), .r (Fresh[22]), .c ({new_AGEMA_signal_1916, LED_128_Instance_SBox_Instance_11_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND3_U1 ( .a ({new_AGEMA_signal_1781, LED_128_Instance_SBox_Instance_11_n3}), .b ({new_AGEMA_signal_1699, LED_128_Instance_addconst_out[46]}), .clk (CLK), .r (Fresh[23]), .c ({new_AGEMA_signal_1854, LED_128_Instance_SBox_Instance_11_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR15_U1 ( .a ({new_AGEMA_signal_2723, new_AGEMA_signal_2721}), .b ({new_AGEMA_signal_1854, LED_128_Instance_SBox_Instance_11_T2}), .c ({new_AGEMA_signal_1917, LED_128_Instance_subcells_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR16_U1 ( .a ({new_AGEMA_signal_1956, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2725}), .c ({new_AGEMA_signal_1988, LED_128_Instance_SBox_Instance_12_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR7_U1 ( .a ({new_AGEMA_signal_1956, LED_128_Instance_SBox_Instance_12_T0}), .b ({new_AGEMA_signal_1922, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_1989, LED_128_Instance_SBox_Instance_12_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR8_U1 ( .a ({new_AGEMA_signal_2731, new_AGEMA_signal_2729}), .b ({new_AGEMA_signal_1989, LED_128_Instance_SBox_Instance_12_L5}), .c ({new_AGEMA_signal_2020, LED_128_Instance_SBox_Instance_12_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND1_U1 ( .a ({new_AGEMA_signal_1918, LED_128_Instance_SBox_Instance_12_n1}), .b ({new_AGEMA_signal_1855, LED_128_Instance_SBox_Instance_12_n2}), .clk (CLK), .r (Fresh[24]), .c ({new_AGEMA_signal_1956, LED_128_Instance_SBox_Instance_12_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND3_U1 ( .a ({new_AGEMA_signal_1856, LED_128_Instance_SBox_Instance_12_n3}), .b ({new_AGEMA_signal_1732, LED_128_Instance_addconst_out[50]}), .clk (CLK), .r (Fresh[25]), .c ({new_AGEMA_signal_1922, LED_128_Instance_SBox_Instance_12_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR15_U1 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2733}), .b ({new_AGEMA_signal_1922, LED_128_Instance_SBox_Instance_12_T2}), .c ({new_AGEMA_signal_1957, LED_128_Instance_subcells_out[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR16_U1 ( .a ({new_AGEMA_signal_1958, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2737}), .c ({new_AGEMA_signal_1990, LED_128_Instance_SBox_Instance_13_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR7_U1 ( .a ({new_AGEMA_signal_1958, LED_128_Instance_SBox_Instance_13_T0}), .b ({new_AGEMA_signal_1927, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_1991, LED_128_Instance_SBox_Instance_13_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR8_U1 ( .a ({new_AGEMA_signal_2743, new_AGEMA_signal_2741}), .b ({new_AGEMA_signal_1991, LED_128_Instance_SBox_Instance_13_L5}), .c ({new_AGEMA_signal_2022, LED_128_Instance_SBox_Instance_13_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND1_U1 ( .a ({new_AGEMA_signal_1923, LED_128_Instance_SBox_Instance_13_n1}), .b ({new_AGEMA_signal_1786, LED_128_Instance_SBox_Instance_13_n2}), .clk (CLK), .r (Fresh[26]), .c ({new_AGEMA_signal_1958, LED_128_Instance_SBox_Instance_13_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND3_U1 ( .a ({new_AGEMA_signal_1861, LED_128_Instance_SBox_Instance_13_n3}), .b ({new_AGEMA_signal_1728, LED_128_Instance_addconst_out[54]}), .clk (CLK), .r (Fresh[27]), .c ({new_AGEMA_signal_1927, LED_128_Instance_SBox_Instance_13_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR15_U1 ( .a ({new_AGEMA_signal_2747, new_AGEMA_signal_2745}), .b ({new_AGEMA_signal_1927, LED_128_Instance_SBox_Instance_13_T2}), .c ({new_AGEMA_signal_1959, LED_128_Instance_subcells_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR16_U1 ( .a ({new_AGEMA_signal_1928, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2749}), .c ({new_AGEMA_signal_1960, LED_128_Instance_SBox_Instance_14_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR7_U1 ( .a ({new_AGEMA_signal_1928, LED_128_Instance_SBox_Instance_14_T0}), .b ({new_AGEMA_signal_1870, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_1961, LED_128_Instance_SBox_Instance_14_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR8_U1 ( .a ({new_AGEMA_signal_2755, new_AGEMA_signal_2753}), .b ({new_AGEMA_signal_1961, LED_128_Instance_SBox_Instance_14_L5}), .c ({new_AGEMA_signal_1992, LED_128_Instance_SBox_Instance_14_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND1_U1 ( .a ({new_AGEMA_signal_1866, LED_128_Instance_SBox_Instance_14_n1}), .b ({new_AGEMA_signal_1787, LED_128_Instance_SBox_Instance_14_n2}), .clk (CLK), .r (Fresh[28]), .c ({new_AGEMA_signal_1928, LED_128_Instance_SBox_Instance_14_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND3_U1 ( .a ({new_AGEMA_signal_1788, LED_128_Instance_SBox_Instance_14_n3}), .b ({new_AGEMA_signal_1711, LED_128_Instance_addconst_out[58]}), .clk (CLK), .r (Fresh[29]), .c ({new_AGEMA_signal_1870, LED_128_Instance_SBox_Instance_14_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR15_U1 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2757}), .b ({new_AGEMA_signal_1870, LED_128_Instance_SBox_Instance_14_T2}), .c ({new_AGEMA_signal_1929, LED_128_Instance_subcells_out[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR16_U1 ( .a ({new_AGEMA_signal_1930, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2761}), .c ({new_AGEMA_signal_1962, LED_128_Instance_SBox_Instance_15_Q2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR7_U1 ( .a ({new_AGEMA_signal_1930, LED_128_Instance_SBox_Instance_15_T0}), .b ({new_AGEMA_signal_1875, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_1963, LED_128_Instance_SBox_Instance_15_L5}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR8_U1 ( .a ({new_AGEMA_signal_2767, new_AGEMA_signal_2765}), .b ({new_AGEMA_signal_1963, LED_128_Instance_SBox_Instance_15_L5}), .c ({new_AGEMA_signal_1994, LED_128_Instance_SBox_Instance_15_Q6}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND1_U1 ( .a ({new_AGEMA_signal_1871, LED_128_Instance_SBox_Instance_15_n1}), .b ({new_AGEMA_signal_1793, LED_128_Instance_SBox_Instance_15_n2}), .clk (CLK), .r (Fresh[30]), .c ({new_AGEMA_signal_1930, LED_128_Instance_SBox_Instance_15_T0}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND3_U1 ( .a ({new_AGEMA_signal_1794, LED_128_Instance_SBox_Instance_15_n3}), .b ({new_AGEMA_signal_1715, LED_128_Instance_addconst_out[62]}), .clk (CLK), .r (Fresh[31]), .c ({new_AGEMA_signal_1875, LED_128_Instance_SBox_Instance_15_T2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR15_U1 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2769}), .b ({new_AGEMA_signal_1875, LED_128_Instance_SBox_Instance_15_T2}), .c ({new_AGEMA_signal_1931, LED_128_Instance_subcells_out[60]}) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (CLK), .D (new_AGEMA_signal_2580), .Q (new_AGEMA_signal_2581) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (CLK), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_2583) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (CLK), .D (new_AGEMA_signal_2584), .Q (new_AGEMA_signal_2585) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (CLK), .D (new_AGEMA_signal_2586), .Q (new_AGEMA_signal_2587) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (CLK), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_2589) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (CLK), .D (new_AGEMA_signal_2590), .Q (new_AGEMA_signal_2591) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (CLK), .D (new_AGEMA_signal_2592), .Q (new_AGEMA_signal_2593) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (CLK), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_2595) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (CLK), .D (new_AGEMA_signal_2596), .Q (new_AGEMA_signal_2597) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (CLK), .D (new_AGEMA_signal_2598), .Q (new_AGEMA_signal_2599) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (CLK), .D (new_AGEMA_signal_2600), .Q (new_AGEMA_signal_2601) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (CLK), .D (new_AGEMA_signal_2602), .Q (new_AGEMA_signal_2603) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (CLK), .D (new_AGEMA_signal_2604), .Q (new_AGEMA_signal_2605) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (CLK), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_2607) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (CLK), .D (new_AGEMA_signal_2608), .Q (new_AGEMA_signal_2609) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (CLK), .D (new_AGEMA_signal_2610), .Q (new_AGEMA_signal_2611) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (CLK), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_2613) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (CLK), .D (new_AGEMA_signal_2614), .Q (new_AGEMA_signal_2615) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (CLK), .D (new_AGEMA_signal_2616), .Q (new_AGEMA_signal_2617) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (CLK), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_2619) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (CLK), .D (new_AGEMA_signal_2620), .Q (new_AGEMA_signal_2621) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (CLK), .D (new_AGEMA_signal_2622), .Q (new_AGEMA_signal_2623) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (CLK), .D (new_AGEMA_signal_2624), .Q (new_AGEMA_signal_2625) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (CLK), .D (new_AGEMA_signal_2626), .Q (new_AGEMA_signal_2627) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (CLK), .D (new_AGEMA_signal_2628), .Q (new_AGEMA_signal_2629) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (CLK), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_2631) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (CLK), .D (new_AGEMA_signal_2632), .Q (new_AGEMA_signal_2633) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (CLK), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_2635) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (CLK), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_2637) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (CLK), .D (new_AGEMA_signal_2638), .Q (new_AGEMA_signal_2639) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (CLK), .D (new_AGEMA_signal_2640), .Q (new_AGEMA_signal_2641) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (CLK), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_2643) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (CLK), .D (new_AGEMA_signal_2644), .Q (new_AGEMA_signal_2645) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (CLK), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_2647) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (CLK), .D (new_AGEMA_signal_2648), .Q (new_AGEMA_signal_2649) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (CLK), .D (new_AGEMA_signal_2650), .Q (new_AGEMA_signal_2651) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (CLK), .D (new_AGEMA_signal_2652), .Q (new_AGEMA_signal_2653) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (CLK), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_2655) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (CLK), .D (new_AGEMA_signal_2656), .Q (new_AGEMA_signal_2657) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (CLK), .D (new_AGEMA_signal_2658), .Q (new_AGEMA_signal_2659) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (CLK), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_2661) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (CLK), .D (new_AGEMA_signal_2662), .Q (new_AGEMA_signal_2663) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (CLK), .D (new_AGEMA_signal_2664), .Q (new_AGEMA_signal_2665) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (CLK), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_2667) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (CLK), .D (new_AGEMA_signal_2668), .Q (new_AGEMA_signal_2669) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (CLK), .D (new_AGEMA_signal_2670), .Q (new_AGEMA_signal_2671) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (CLK), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_2673) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (CLK), .D (new_AGEMA_signal_2674), .Q (new_AGEMA_signal_2675) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (CLK), .D (new_AGEMA_signal_2676), .Q (new_AGEMA_signal_2677) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (CLK), .D (new_AGEMA_signal_2678), .Q (new_AGEMA_signal_2679) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (CLK), .D (new_AGEMA_signal_2680), .Q (new_AGEMA_signal_2681) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (CLK), .D (new_AGEMA_signal_2682), .Q (new_AGEMA_signal_2683) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (CLK), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_2685) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (CLK), .D (new_AGEMA_signal_2686), .Q (new_AGEMA_signal_2687) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (CLK), .D (new_AGEMA_signal_2688), .Q (new_AGEMA_signal_2689) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (CLK), .D (new_AGEMA_signal_2690), .Q (new_AGEMA_signal_2691) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (CLK), .D (new_AGEMA_signal_2692), .Q (new_AGEMA_signal_2693) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (CLK), .D (new_AGEMA_signal_2694), .Q (new_AGEMA_signal_2695) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (CLK), .D (new_AGEMA_signal_2696), .Q (new_AGEMA_signal_2697) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (CLK), .D (new_AGEMA_signal_2698), .Q (new_AGEMA_signal_2699) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (CLK), .D (new_AGEMA_signal_2700), .Q (new_AGEMA_signal_2701) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (CLK), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_2703) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (CLK), .D (new_AGEMA_signal_2704), .Q (new_AGEMA_signal_2705) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (CLK), .D (new_AGEMA_signal_2706), .Q (new_AGEMA_signal_2707) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (CLK), .D (new_AGEMA_signal_2708), .Q (new_AGEMA_signal_2709) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (CLK), .D (new_AGEMA_signal_2710), .Q (new_AGEMA_signal_2711) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (CLK), .D (new_AGEMA_signal_2712), .Q (new_AGEMA_signal_2713) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (CLK), .D (new_AGEMA_signal_2714), .Q (new_AGEMA_signal_2715) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (CLK), .D (new_AGEMA_signal_2716), .Q (new_AGEMA_signal_2717) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (CLK), .D (new_AGEMA_signal_2718), .Q (new_AGEMA_signal_2719) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (CLK), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_2721) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (CLK), .D (new_AGEMA_signal_2722), .Q (new_AGEMA_signal_2723) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (CLK), .D (new_AGEMA_signal_2724), .Q (new_AGEMA_signal_2725) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (CLK), .D (new_AGEMA_signal_2726), .Q (new_AGEMA_signal_2727) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (CLK), .D (new_AGEMA_signal_2728), .Q (new_AGEMA_signal_2729) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (CLK), .D (new_AGEMA_signal_2730), .Q (new_AGEMA_signal_2731) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (CLK), .D (new_AGEMA_signal_2732), .Q (new_AGEMA_signal_2733) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (CLK), .D (new_AGEMA_signal_2734), .Q (new_AGEMA_signal_2735) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (CLK), .D (new_AGEMA_signal_2736), .Q (new_AGEMA_signal_2737) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (CLK), .D (new_AGEMA_signal_2738), .Q (new_AGEMA_signal_2739) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (CLK), .D (new_AGEMA_signal_2740), .Q (new_AGEMA_signal_2741) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (CLK), .D (new_AGEMA_signal_2742), .Q (new_AGEMA_signal_2743) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (CLK), .D (new_AGEMA_signal_2744), .Q (new_AGEMA_signal_2745) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (CLK), .D (new_AGEMA_signal_2746), .Q (new_AGEMA_signal_2747) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (CLK), .D (new_AGEMA_signal_2748), .Q (new_AGEMA_signal_2749) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (CLK), .D (new_AGEMA_signal_2750), .Q (new_AGEMA_signal_2751) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (CLK), .D (new_AGEMA_signal_2752), .Q (new_AGEMA_signal_2753) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (CLK), .D (new_AGEMA_signal_2754), .Q (new_AGEMA_signal_2755) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (CLK), .D (new_AGEMA_signal_2756), .Q (new_AGEMA_signal_2757) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (CLK), .D (new_AGEMA_signal_2758), .Q (new_AGEMA_signal_2759) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (CLK), .D (new_AGEMA_signal_2760), .Q (new_AGEMA_signal_2761) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (CLK), .D (new_AGEMA_signal_2762), .Q (new_AGEMA_signal_2763) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (CLK), .D (new_AGEMA_signal_2764), .Q (new_AGEMA_signal_2765) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (CLK), .D (new_AGEMA_signal_2766), .Q (new_AGEMA_signal_2767) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (CLK), .D (new_AGEMA_signal_2768), .Q (new_AGEMA_signal_2769) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (CLK), .D (new_AGEMA_signal_2770), .Q (new_AGEMA_signal_2771) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (CLK), .D (new_AGEMA_signal_2772), .Q (new_AGEMA_signal_2773) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (CLK), .D (new_AGEMA_signal_2776), .Q (new_AGEMA_signal_2777) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (CLK), .D (new_AGEMA_signal_2780), .Q (new_AGEMA_signal_2781) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (CLK), .D (new_AGEMA_signal_2784), .Q (new_AGEMA_signal_2785) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (CLK), .D (new_AGEMA_signal_2788), .Q (new_AGEMA_signal_2789) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (CLK), .D (new_AGEMA_signal_2792), .Q (new_AGEMA_signal_2793) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (CLK), .D (new_AGEMA_signal_2796), .Q (new_AGEMA_signal_2797) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (CLK), .D (new_AGEMA_signal_2800), .Q (new_AGEMA_signal_2801) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (CLK), .D (new_AGEMA_signal_2804), .Q (new_AGEMA_signal_2805) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (CLK), .D (new_AGEMA_signal_2808), .Q (new_AGEMA_signal_2809) ) ;
    buf_clk new_AGEMA_reg_buffer_1361 ( .C (CLK), .D (new_AGEMA_signal_2812), .Q (new_AGEMA_signal_2813) ) ;
    buf_clk new_AGEMA_reg_buffer_1365 ( .C (CLK), .D (new_AGEMA_signal_2816), .Q (new_AGEMA_signal_2817) ) ;
    buf_clk new_AGEMA_reg_buffer_1369 ( .C (CLK), .D (new_AGEMA_signal_2820), .Q (new_AGEMA_signal_2821) ) ;
    buf_clk new_AGEMA_reg_buffer_1373 ( .C (CLK), .D (new_AGEMA_signal_2824), .Q (new_AGEMA_signal_2825) ) ;
    buf_clk new_AGEMA_reg_buffer_1377 ( .C (CLK), .D (new_AGEMA_signal_2828), .Q (new_AGEMA_signal_2829) ) ;
    buf_clk new_AGEMA_reg_buffer_1381 ( .C (CLK), .D (new_AGEMA_signal_2832), .Q (new_AGEMA_signal_2833) ) ;
    buf_clk new_AGEMA_reg_buffer_1385 ( .C (CLK), .D (new_AGEMA_signal_2836), .Q (new_AGEMA_signal_2837) ) ;
    buf_clk new_AGEMA_reg_buffer_1389 ( .C (CLK), .D (new_AGEMA_signal_2840), .Q (new_AGEMA_signal_2841) ) ;
    buf_clk new_AGEMA_reg_buffer_1393 ( .C (CLK), .D (new_AGEMA_signal_2844), .Q (new_AGEMA_signal_2845) ) ;
    buf_clk new_AGEMA_reg_buffer_1397 ( .C (CLK), .D (new_AGEMA_signal_2848), .Q (new_AGEMA_signal_2849) ) ;
    buf_clk new_AGEMA_reg_buffer_1401 ( .C (CLK), .D (new_AGEMA_signal_2852), .Q (new_AGEMA_signal_2853) ) ;
    buf_clk new_AGEMA_reg_buffer_1405 ( .C (CLK), .D (new_AGEMA_signal_2856), .Q (new_AGEMA_signal_2857) ) ;
    buf_clk new_AGEMA_reg_buffer_1409 ( .C (CLK), .D (new_AGEMA_signal_2860), .Q (new_AGEMA_signal_2861) ) ;
    buf_clk new_AGEMA_reg_buffer_1413 ( .C (CLK), .D (new_AGEMA_signal_2864), .Q (new_AGEMA_signal_2865) ) ;
    buf_clk new_AGEMA_reg_buffer_1417 ( .C (CLK), .D (new_AGEMA_signal_2868), .Q (new_AGEMA_signal_2869) ) ;
    buf_clk new_AGEMA_reg_buffer_1421 ( .C (CLK), .D (new_AGEMA_signal_2872), .Q (new_AGEMA_signal_2873) ) ;
    buf_clk new_AGEMA_reg_buffer_1425 ( .C (CLK), .D (new_AGEMA_signal_2876), .Q (new_AGEMA_signal_2877) ) ;
    buf_clk new_AGEMA_reg_buffer_1429 ( .C (CLK), .D (new_AGEMA_signal_2880), .Q (new_AGEMA_signal_2881) ) ;
    buf_clk new_AGEMA_reg_buffer_1433 ( .C (CLK), .D (new_AGEMA_signal_2884), .Q (new_AGEMA_signal_2885) ) ;
    buf_clk new_AGEMA_reg_buffer_1437 ( .C (CLK), .D (new_AGEMA_signal_2888), .Q (new_AGEMA_signal_2889) ) ;
    buf_clk new_AGEMA_reg_buffer_1441 ( .C (CLK), .D (new_AGEMA_signal_2892), .Q (new_AGEMA_signal_2893) ) ;
    buf_clk new_AGEMA_reg_buffer_1445 ( .C (CLK), .D (new_AGEMA_signal_2896), .Q (new_AGEMA_signal_2897) ) ;
    buf_clk new_AGEMA_reg_buffer_1449 ( .C (CLK), .D (new_AGEMA_signal_2900), .Q (new_AGEMA_signal_2901) ) ;
    buf_clk new_AGEMA_reg_buffer_1453 ( .C (CLK), .D (new_AGEMA_signal_2904), .Q (new_AGEMA_signal_2905) ) ;
    buf_clk new_AGEMA_reg_buffer_1457 ( .C (CLK), .D (new_AGEMA_signal_2908), .Q (new_AGEMA_signal_2909) ) ;
    buf_clk new_AGEMA_reg_buffer_1461 ( .C (CLK), .D (new_AGEMA_signal_2912), .Q (new_AGEMA_signal_2913) ) ;
    buf_clk new_AGEMA_reg_buffer_1465 ( .C (CLK), .D (new_AGEMA_signal_2916), .Q (new_AGEMA_signal_2917) ) ;
    buf_clk new_AGEMA_reg_buffer_1469 ( .C (CLK), .D (new_AGEMA_signal_2920), .Q (new_AGEMA_signal_2921) ) ;
    buf_clk new_AGEMA_reg_buffer_1473 ( .C (CLK), .D (new_AGEMA_signal_2924), .Q (new_AGEMA_signal_2925) ) ;
    buf_clk new_AGEMA_reg_buffer_1477 ( .C (CLK), .D (new_AGEMA_signal_2928), .Q (new_AGEMA_signal_2929) ) ;
    buf_clk new_AGEMA_reg_buffer_1481 ( .C (CLK), .D (new_AGEMA_signal_2932), .Q (new_AGEMA_signal_2933) ) ;
    buf_clk new_AGEMA_reg_buffer_1485 ( .C (CLK), .D (new_AGEMA_signal_2936), .Q (new_AGEMA_signal_2937) ) ;
    buf_clk new_AGEMA_reg_buffer_1489 ( .C (CLK), .D (new_AGEMA_signal_2940), .Q (new_AGEMA_signal_2941) ) ;
    buf_clk new_AGEMA_reg_buffer_1493 ( .C (CLK), .D (new_AGEMA_signal_2944), .Q (new_AGEMA_signal_2945) ) ;
    buf_clk new_AGEMA_reg_buffer_1497 ( .C (CLK), .D (new_AGEMA_signal_2948), .Q (new_AGEMA_signal_2949) ) ;
    buf_clk new_AGEMA_reg_buffer_1501 ( .C (CLK), .D (new_AGEMA_signal_2952), .Q (new_AGEMA_signal_2953) ) ;
    buf_clk new_AGEMA_reg_buffer_1505 ( .C (CLK), .D (new_AGEMA_signal_2956), .Q (new_AGEMA_signal_2957) ) ;
    buf_clk new_AGEMA_reg_buffer_1509 ( .C (CLK), .D (new_AGEMA_signal_2960), .Q (new_AGEMA_signal_2961) ) ;
    buf_clk new_AGEMA_reg_buffer_1513 ( .C (CLK), .D (new_AGEMA_signal_2964), .Q (new_AGEMA_signal_2965) ) ;
    buf_clk new_AGEMA_reg_buffer_1517 ( .C (CLK), .D (new_AGEMA_signal_2968), .Q (new_AGEMA_signal_2969) ) ;
    buf_clk new_AGEMA_reg_buffer_1521 ( .C (CLK), .D (new_AGEMA_signal_2972), .Q (new_AGEMA_signal_2973) ) ;
    buf_clk new_AGEMA_reg_buffer_1525 ( .C (CLK), .D (new_AGEMA_signal_2976), .Q (new_AGEMA_signal_2977) ) ;
    buf_clk new_AGEMA_reg_buffer_1529 ( .C (CLK), .D (new_AGEMA_signal_2980), .Q (new_AGEMA_signal_2981) ) ;
    buf_clk new_AGEMA_reg_buffer_1533 ( .C (CLK), .D (new_AGEMA_signal_2984), .Q (new_AGEMA_signal_2985) ) ;
    buf_clk new_AGEMA_reg_buffer_1537 ( .C (CLK), .D (new_AGEMA_signal_2988), .Q (new_AGEMA_signal_2989) ) ;
    buf_clk new_AGEMA_reg_buffer_1541 ( .C (CLK), .D (new_AGEMA_signal_2992), .Q (new_AGEMA_signal_2993) ) ;
    buf_clk new_AGEMA_reg_buffer_1545 ( .C (CLK), .D (new_AGEMA_signal_2996), .Q (new_AGEMA_signal_2997) ) ;
    buf_clk new_AGEMA_reg_buffer_1549 ( .C (CLK), .D (new_AGEMA_signal_3000), .Q (new_AGEMA_signal_3001) ) ;
    buf_clk new_AGEMA_reg_buffer_1553 ( .C (CLK), .D (new_AGEMA_signal_3004), .Q (new_AGEMA_signal_3005) ) ;
    buf_clk new_AGEMA_reg_buffer_1557 ( .C (CLK), .D (new_AGEMA_signal_3008), .Q (new_AGEMA_signal_3009) ) ;
    buf_clk new_AGEMA_reg_buffer_1561 ( .C (CLK), .D (new_AGEMA_signal_3012), .Q (new_AGEMA_signal_3013) ) ;
    buf_clk new_AGEMA_reg_buffer_1565 ( .C (CLK), .D (new_AGEMA_signal_3016), .Q (new_AGEMA_signal_3017) ) ;
    buf_clk new_AGEMA_reg_buffer_1569 ( .C (CLK), .D (new_AGEMA_signal_3020), .Q (new_AGEMA_signal_3021) ) ;
    buf_clk new_AGEMA_reg_buffer_1573 ( .C (CLK), .D (new_AGEMA_signal_3024), .Q (new_AGEMA_signal_3025) ) ;
    buf_clk new_AGEMA_reg_buffer_1577 ( .C (CLK), .D (new_AGEMA_signal_3028), .Q (new_AGEMA_signal_3029) ) ;
    buf_clk new_AGEMA_reg_buffer_1581 ( .C (CLK), .D (new_AGEMA_signal_3032), .Q (new_AGEMA_signal_3033) ) ;
    buf_clk new_AGEMA_reg_buffer_1585 ( .C (CLK), .D (new_AGEMA_signal_3036), .Q (new_AGEMA_signal_3037) ) ;
    buf_clk new_AGEMA_reg_buffer_1589 ( .C (CLK), .D (new_AGEMA_signal_3040), .Q (new_AGEMA_signal_3041) ) ;
    buf_clk new_AGEMA_reg_buffer_1593 ( .C (CLK), .D (new_AGEMA_signal_3044), .Q (new_AGEMA_signal_3045) ) ;
    buf_clk new_AGEMA_reg_buffer_1597 ( .C (CLK), .D (new_AGEMA_signal_3048), .Q (new_AGEMA_signal_3049) ) ;
    buf_clk new_AGEMA_reg_buffer_1601 ( .C (CLK), .D (new_AGEMA_signal_3052), .Q (new_AGEMA_signal_3053) ) ;
    buf_clk new_AGEMA_reg_buffer_1605 ( .C (CLK), .D (new_AGEMA_signal_3056), .Q (new_AGEMA_signal_3057) ) ;
    buf_clk new_AGEMA_reg_buffer_1609 ( .C (CLK), .D (new_AGEMA_signal_3060), .Q (new_AGEMA_signal_3061) ) ;
    buf_clk new_AGEMA_reg_buffer_1613 ( .C (CLK), .D (new_AGEMA_signal_3064), .Q (new_AGEMA_signal_3065) ) ;
    buf_clk new_AGEMA_reg_buffer_1617 ( .C (CLK), .D (new_AGEMA_signal_3068), .Q (new_AGEMA_signal_3069) ) ;
    buf_clk new_AGEMA_reg_buffer_1621 ( .C (CLK), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_3073) ) ;
    buf_clk new_AGEMA_reg_buffer_1625 ( .C (CLK), .D (new_AGEMA_signal_3076), .Q (new_AGEMA_signal_3077) ) ;
    buf_clk new_AGEMA_reg_buffer_1629 ( .C (CLK), .D (new_AGEMA_signal_3080), .Q (new_AGEMA_signal_3081) ) ;
    buf_clk new_AGEMA_reg_buffer_1633 ( .C (CLK), .D (new_AGEMA_signal_3084), .Q (new_AGEMA_signal_3085) ) ;
    buf_clk new_AGEMA_reg_buffer_1637 ( .C (CLK), .D (new_AGEMA_signal_3088), .Q (new_AGEMA_signal_3089) ) ;
    buf_clk new_AGEMA_reg_buffer_1641 ( .C (CLK), .D (new_AGEMA_signal_3092), .Q (new_AGEMA_signal_3093) ) ;
    buf_clk new_AGEMA_reg_buffer_1645 ( .C (CLK), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_3097) ) ;
    buf_clk new_AGEMA_reg_buffer_1649 ( .C (CLK), .D (new_AGEMA_signal_3100), .Q (new_AGEMA_signal_3101) ) ;
    buf_clk new_AGEMA_reg_buffer_1653 ( .C (CLK), .D (new_AGEMA_signal_3104), .Q (new_AGEMA_signal_3105) ) ;
    buf_clk new_AGEMA_reg_buffer_1657 ( .C (CLK), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_3109) ) ;
    buf_clk new_AGEMA_reg_buffer_1661 ( .C (CLK), .D (new_AGEMA_signal_3112), .Q (new_AGEMA_signal_3113) ) ;
    buf_clk new_AGEMA_reg_buffer_1665 ( .C (CLK), .D (new_AGEMA_signal_3116), .Q (new_AGEMA_signal_3117) ) ;
    buf_clk new_AGEMA_reg_buffer_1669 ( .C (CLK), .D (new_AGEMA_signal_3120), .Q (new_AGEMA_signal_3121) ) ;
    buf_clk new_AGEMA_reg_buffer_1673 ( .C (CLK), .D (new_AGEMA_signal_3124), .Q (new_AGEMA_signal_3125) ) ;
    buf_clk new_AGEMA_reg_buffer_1677 ( .C (CLK), .D (new_AGEMA_signal_3128), .Q (new_AGEMA_signal_3129) ) ;
    buf_clk new_AGEMA_reg_buffer_1681 ( .C (CLK), .D (new_AGEMA_signal_3132), .Q (new_AGEMA_signal_3133) ) ;
    buf_clk new_AGEMA_reg_buffer_1685 ( .C (CLK), .D (new_AGEMA_signal_3136), .Q (new_AGEMA_signal_3137) ) ;
    buf_clk new_AGEMA_reg_buffer_1689 ( .C (CLK), .D (new_AGEMA_signal_3140), .Q (new_AGEMA_signal_3141) ) ;
    buf_clk new_AGEMA_reg_buffer_1693 ( .C (CLK), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_3145) ) ;
    buf_clk new_AGEMA_reg_buffer_1697 ( .C (CLK), .D (new_AGEMA_signal_3148), .Q (new_AGEMA_signal_3149) ) ;
    buf_clk new_AGEMA_reg_buffer_1701 ( .C (CLK), .D (new_AGEMA_signal_3152), .Q (new_AGEMA_signal_3153) ) ;
    buf_clk new_AGEMA_reg_buffer_1705 ( .C (CLK), .D (new_AGEMA_signal_3156), .Q (new_AGEMA_signal_3157) ) ;
    buf_clk new_AGEMA_reg_buffer_1709 ( .C (CLK), .D (new_AGEMA_signal_3160), .Q (new_AGEMA_signal_3161) ) ;
    buf_clk new_AGEMA_reg_buffer_1713 ( .C (CLK), .D (new_AGEMA_signal_3164), .Q (new_AGEMA_signal_3165) ) ;
    buf_clk new_AGEMA_reg_buffer_1717 ( .C (CLK), .D (new_AGEMA_signal_3168), .Q (new_AGEMA_signal_3169) ) ;
    buf_clk new_AGEMA_reg_buffer_1721 ( .C (CLK), .D (new_AGEMA_signal_3172), .Q (new_AGEMA_signal_3173) ) ;
    buf_clk new_AGEMA_reg_buffer_1725 ( .C (CLK), .D (new_AGEMA_signal_3176), .Q (new_AGEMA_signal_3177) ) ;
    buf_clk new_AGEMA_reg_buffer_1729 ( .C (CLK), .D (new_AGEMA_signal_3180), .Q (new_AGEMA_signal_3181) ) ;
    buf_clk new_AGEMA_reg_buffer_1733 ( .C (CLK), .D (new_AGEMA_signal_3184), .Q (new_AGEMA_signal_3185) ) ;
    buf_clk new_AGEMA_reg_buffer_1737 ( .C (CLK), .D (new_AGEMA_signal_3188), .Q (new_AGEMA_signal_3189) ) ;
    buf_clk new_AGEMA_reg_buffer_1741 ( .C (CLK), .D (new_AGEMA_signal_3192), .Q (new_AGEMA_signal_3193) ) ;
    buf_clk new_AGEMA_reg_buffer_1745 ( .C (CLK), .D (new_AGEMA_signal_3196), .Q (new_AGEMA_signal_3197) ) ;
    buf_clk new_AGEMA_reg_buffer_1749 ( .C (CLK), .D (new_AGEMA_signal_3200), .Q (new_AGEMA_signal_3201) ) ;
    buf_clk new_AGEMA_reg_buffer_1753 ( .C (CLK), .D (new_AGEMA_signal_3204), .Q (new_AGEMA_signal_3205) ) ;
    buf_clk new_AGEMA_reg_buffer_1757 ( .C (CLK), .D (new_AGEMA_signal_3208), .Q (new_AGEMA_signal_3209) ) ;
    buf_clk new_AGEMA_reg_buffer_1761 ( .C (CLK), .D (new_AGEMA_signal_3212), .Q (new_AGEMA_signal_3213) ) ;
    buf_clk new_AGEMA_reg_buffer_1765 ( .C (CLK), .D (new_AGEMA_signal_3216), .Q (new_AGEMA_signal_3217) ) ;
    buf_clk new_AGEMA_reg_buffer_1769 ( .C (CLK), .D (new_AGEMA_signal_3220), .Q (new_AGEMA_signal_3221) ) ;
    buf_clk new_AGEMA_reg_buffer_1773 ( .C (CLK), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_3225) ) ;
    buf_clk new_AGEMA_reg_buffer_1777 ( .C (CLK), .D (new_AGEMA_signal_3228), .Q (new_AGEMA_signal_3229) ) ;
    buf_clk new_AGEMA_reg_buffer_1781 ( .C (CLK), .D (new_AGEMA_signal_3232), .Q (new_AGEMA_signal_3233) ) ;
    buf_clk new_AGEMA_reg_buffer_1785 ( .C (CLK), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_3237) ) ;
    buf_clk new_AGEMA_reg_buffer_1789 ( .C (CLK), .D (new_AGEMA_signal_3240), .Q (new_AGEMA_signal_3241) ) ;
    buf_clk new_AGEMA_reg_buffer_1793 ( .C (CLK), .D (new_AGEMA_signal_3244), .Q (new_AGEMA_signal_3245) ) ;
    buf_clk new_AGEMA_reg_buffer_1797 ( .C (CLK), .D (new_AGEMA_signal_3248), .Q (new_AGEMA_signal_3249) ) ;
    buf_clk new_AGEMA_reg_buffer_1801 ( .C (CLK), .D (new_AGEMA_signal_3252), .Q (new_AGEMA_signal_3253) ) ;
    buf_clk new_AGEMA_reg_buffer_1805 ( .C (CLK), .D (new_AGEMA_signal_3256), .Q (new_AGEMA_signal_3257) ) ;
    buf_clk new_AGEMA_reg_buffer_1809 ( .C (CLK), .D (new_AGEMA_signal_3260), .Q (new_AGEMA_signal_3261) ) ;
    buf_clk new_AGEMA_reg_buffer_1813 ( .C (CLK), .D (new_AGEMA_signal_3264), .Q (new_AGEMA_signal_3265) ) ;
    buf_clk new_AGEMA_reg_buffer_1817 ( .C (CLK), .D (new_AGEMA_signal_3268), .Q (new_AGEMA_signal_3269) ) ;
    buf_clk new_AGEMA_reg_buffer_1821 ( .C (CLK), .D (new_AGEMA_signal_3272), .Q (new_AGEMA_signal_3273) ) ;
    buf_clk new_AGEMA_reg_buffer_1825 ( .C (CLK), .D (new_AGEMA_signal_3276), .Q (new_AGEMA_signal_3277) ) ;
    buf_clk new_AGEMA_reg_buffer_1829 ( .C (CLK), .D (new_AGEMA_signal_3280), .Q (new_AGEMA_signal_3281) ) ;
    buf_clk new_AGEMA_reg_buffer_1833 ( .C (CLK), .D (new_AGEMA_signal_3284), .Q (new_AGEMA_signal_3285) ) ;
    buf_clk new_AGEMA_reg_buffer_1837 ( .C (CLK), .D (new_AGEMA_signal_3288), .Q (new_AGEMA_signal_3289) ) ;
    buf_clk new_AGEMA_reg_buffer_1841 ( .C (CLK), .D (new_AGEMA_signal_3292), .Q (new_AGEMA_signal_3293) ) ;
    buf_clk new_AGEMA_reg_buffer_1845 ( .C (CLK), .D (new_AGEMA_signal_3296), .Q (new_AGEMA_signal_3297) ) ;
    buf_clk new_AGEMA_reg_buffer_1849 ( .C (CLK), .D (new_AGEMA_signal_3300), .Q (new_AGEMA_signal_3301) ) ;
    buf_clk new_AGEMA_reg_buffer_1853 ( .C (CLK), .D (new_AGEMA_signal_3304), .Q (new_AGEMA_signal_3305) ) ;
    buf_clk new_AGEMA_reg_buffer_1857 ( .C (CLK), .D (new_AGEMA_signal_3308), .Q (new_AGEMA_signal_3309) ) ;
    buf_clk new_AGEMA_reg_buffer_1861 ( .C (CLK), .D (new_AGEMA_signal_3312), .Q (new_AGEMA_signal_3313) ) ;
    buf_clk new_AGEMA_reg_buffer_1865 ( .C (CLK), .D (new_AGEMA_signal_3316), .Q (new_AGEMA_signal_3317) ) ;
    buf_clk new_AGEMA_reg_buffer_1869 ( .C (CLK), .D (new_AGEMA_signal_3320), .Q (new_AGEMA_signal_3321) ) ;
    buf_clk new_AGEMA_reg_buffer_1873 ( .C (CLK), .D (new_AGEMA_signal_3324), .Q (new_AGEMA_signal_3325) ) ;
    buf_clk new_AGEMA_reg_buffer_1877 ( .C (CLK), .D (new_AGEMA_signal_3328), .Q (new_AGEMA_signal_3329) ) ;
    buf_clk new_AGEMA_reg_buffer_1881 ( .C (CLK), .D (new_AGEMA_signal_3332), .Q (new_AGEMA_signal_3333) ) ;
    buf_clk new_AGEMA_reg_buffer_1885 ( .C (CLK), .D (new_AGEMA_signal_3336), .Q (new_AGEMA_signal_3337) ) ;
    buf_clk new_AGEMA_reg_buffer_1889 ( .C (CLK), .D (new_AGEMA_signal_3340), .Q (new_AGEMA_signal_3341) ) ;
    buf_clk new_AGEMA_reg_buffer_1893 ( .C (CLK), .D (new_AGEMA_signal_3344), .Q (new_AGEMA_signal_3345) ) ;
    buf_clk new_AGEMA_reg_buffer_1897 ( .C (CLK), .D (new_AGEMA_signal_3348), .Q (new_AGEMA_signal_3349) ) ;
    buf_clk new_AGEMA_reg_buffer_1901 ( .C (CLK), .D (new_AGEMA_signal_3352), .Q (new_AGEMA_signal_3353) ) ;
    buf_clk new_AGEMA_reg_buffer_1905 ( .C (CLK), .D (new_AGEMA_signal_3356), .Q (new_AGEMA_signal_3357) ) ;
    buf_clk new_AGEMA_reg_buffer_1909 ( .C (CLK), .D (new_AGEMA_signal_3360), .Q (new_AGEMA_signal_3361) ) ;
    buf_clk new_AGEMA_reg_buffer_1913 ( .C (CLK), .D (new_AGEMA_signal_3364), .Q (new_AGEMA_signal_3365) ) ;
    buf_clk new_AGEMA_reg_buffer_1917 ( .C (CLK), .D (new_AGEMA_signal_3368), .Q (new_AGEMA_signal_3369) ) ;
    buf_clk new_AGEMA_reg_buffer_1921 ( .C (CLK), .D (new_AGEMA_signal_3372), .Q (new_AGEMA_signal_3373) ) ;
    buf_clk new_AGEMA_reg_buffer_1925 ( .C (CLK), .D (new_AGEMA_signal_3376), .Q (new_AGEMA_signal_3377) ) ;
    buf_clk new_AGEMA_reg_buffer_1929 ( .C (CLK), .D (new_AGEMA_signal_3380), .Q (new_AGEMA_signal_3381) ) ;
    buf_clk new_AGEMA_reg_buffer_1933 ( .C (CLK), .D (new_AGEMA_signal_3384), .Q (new_AGEMA_signal_3385) ) ;
    buf_clk new_AGEMA_reg_buffer_1937 ( .C (CLK), .D (new_AGEMA_signal_3388), .Q (new_AGEMA_signal_3389) ) ;
    buf_clk new_AGEMA_reg_buffer_1941 ( .C (CLK), .D (new_AGEMA_signal_3392), .Q (new_AGEMA_signal_3393) ) ;
    buf_clk new_AGEMA_reg_buffer_1945 ( .C (CLK), .D (new_AGEMA_signal_3396), .Q (new_AGEMA_signal_3397) ) ;
    buf_clk new_AGEMA_reg_buffer_1949 ( .C (CLK), .D (new_AGEMA_signal_3400), .Q (new_AGEMA_signal_3401) ) ;
    buf_clk new_AGEMA_reg_buffer_1953 ( .C (CLK), .D (new_AGEMA_signal_3404), .Q (new_AGEMA_signal_3405) ) ;
    buf_clk new_AGEMA_reg_buffer_1957 ( .C (CLK), .D (new_AGEMA_signal_3408), .Q (new_AGEMA_signal_3409) ) ;
    buf_clk new_AGEMA_reg_buffer_1961 ( .C (CLK), .D (new_AGEMA_signal_3412), .Q (new_AGEMA_signal_3413) ) ;
    buf_clk new_AGEMA_reg_buffer_1965 ( .C (CLK), .D (new_AGEMA_signal_3416), .Q (new_AGEMA_signal_3417) ) ;
    buf_clk new_AGEMA_reg_buffer_1969 ( .C (CLK), .D (new_AGEMA_signal_3420), .Q (new_AGEMA_signal_3421) ) ;
    buf_clk new_AGEMA_reg_buffer_1973 ( .C (CLK), .D (new_AGEMA_signal_3424), .Q (new_AGEMA_signal_3425) ) ;
    buf_clk new_AGEMA_reg_buffer_1977 ( .C (CLK), .D (new_AGEMA_signal_3428), .Q (new_AGEMA_signal_3429) ) ;
    buf_clk new_AGEMA_reg_buffer_1981 ( .C (CLK), .D (new_AGEMA_signal_3432), .Q (new_AGEMA_signal_3433) ) ;
    buf_clk new_AGEMA_reg_buffer_1985 ( .C (CLK), .D (new_AGEMA_signal_3436), .Q (new_AGEMA_signal_3437) ) ;
    buf_clk new_AGEMA_reg_buffer_1989 ( .C (CLK), .D (new_AGEMA_signal_3440), .Q (new_AGEMA_signal_3441) ) ;
    buf_clk new_AGEMA_reg_buffer_1993 ( .C (CLK), .D (new_AGEMA_signal_3444), .Q (new_AGEMA_signal_3445) ) ;
    buf_clk new_AGEMA_reg_buffer_1997 ( .C (CLK), .D (new_AGEMA_signal_3448), .Q (new_AGEMA_signal_3449) ) ;
    buf_clk new_AGEMA_reg_buffer_2001 ( .C (CLK), .D (new_AGEMA_signal_3452), .Q (new_AGEMA_signal_3453) ) ;
    buf_clk new_AGEMA_reg_buffer_2005 ( .C (CLK), .D (new_AGEMA_signal_3456), .Q (new_AGEMA_signal_3457) ) ;
    buf_clk new_AGEMA_reg_buffer_2009 ( .C (CLK), .D (new_AGEMA_signal_3460), .Q (new_AGEMA_signal_3461) ) ;
    buf_clk new_AGEMA_reg_buffer_2013 ( .C (CLK), .D (new_AGEMA_signal_3464), .Q (new_AGEMA_signal_3465) ) ;
    buf_clk new_AGEMA_reg_buffer_2017 ( .C (CLK), .D (new_AGEMA_signal_3468), .Q (new_AGEMA_signal_3469) ) ;
    buf_clk new_AGEMA_reg_buffer_2021 ( .C (CLK), .D (new_AGEMA_signal_3472), .Q (new_AGEMA_signal_3473) ) ;
    buf_clk new_AGEMA_reg_buffer_2025 ( .C (CLK), .D (new_AGEMA_signal_3476), .Q (new_AGEMA_signal_3477) ) ;
    buf_clk new_AGEMA_reg_buffer_2029 ( .C (CLK), .D (new_AGEMA_signal_3480), .Q (new_AGEMA_signal_3481) ) ;
    buf_clk new_AGEMA_reg_buffer_2033 ( .C (CLK), .D (new_AGEMA_signal_3484), .Q (new_AGEMA_signal_3485) ) ;
    buf_clk new_AGEMA_reg_buffer_2037 ( .C (CLK), .D (new_AGEMA_signal_3488), .Q (new_AGEMA_signal_3489) ) ;
    buf_clk new_AGEMA_reg_buffer_2041 ( .C (CLK), .D (new_AGEMA_signal_3492), .Q (new_AGEMA_signal_3493) ) ;
    buf_clk new_AGEMA_reg_buffer_2045 ( .C (CLK), .D (new_AGEMA_signal_3496), .Q (new_AGEMA_signal_3497) ) ;
    buf_clk new_AGEMA_reg_buffer_2049 ( .C (CLK), .D (new_AGEMA_signal_3500), .Q (new_AGEMA_signal_3501) ) ;
    buf_clk new_AGEMA_reg_buffer_2053 ( .C (CLK), .D (new_AGEMA_signal_3504), .Q (new_AGEMA_signal_3505) ) ;
    buf_clk new_AGEMA_reg_buffer_2057 ( .C (CLK), .D (new_AGEMA_signal_3508), .Q (new_AGEMA_signal_3509) ) ;
    buf_clk new_AGEMA_reg_buffer_2061 ( .C (CLK), .D (new_AGEMA_signal_3512), .Q (new_AGEMA_signal_3513) ) ;
    buf_clk new_AGEMA_reg_buffer_2065 ( .C (CLK), .D (new_AGEMA_signal_3516), .Q (new_AGEMA_signal_3517) ) ;
    buf_clk new_AGEMA_reg_buffer_2069 ( .C (CLK), .D (new_AGEMA_signal_3520), .Q (new_AGEMA_signal_3521) ) ;
    buf_clk new_AGEMA_reg_buffer_2073 ( .C (CLK), .D (new_AGEMA_signal_3524), .Q (new_AGEMA_signal_3525) ) ;
    buf_clk new_AGEMA_reg_buffer_2077 ( .C (CLK), .D (new_AGEMA_signal_3528), .Q (new_AGEMA_signal_3529) ) ;
    buf_clk new_AGEMA_reg_buffer_2081 ( .C (CLK), .D (new_AGEMA_signal_3532), .Q (new_AGEMA_signal_3533) ) ;
    buf_clk new_AGEMA_reg_buffer_2085 ( .C (CLK), .D (new_AGEMA_signal_3536), .Q (new_AGEMA_signal_3537) ) ;
    buf_clk new_AGEMA_reg_buffer_2089 ( .C (CLK), .D (new_AGEMA_signal_3540), .Q (new_AGEMA_signal_3541) ) ;
    buf_clk new_AGEMA_reg_buffer_2093 ( .C (CLK), .D (new_AGEMA_signal_3544), .Q (new_AGEMA_signal_3545) ) ;
    buf_clk new_AGEMA_reg_buffer_2097 ( .C (CLK), .D (new_AGEMA_signal_3548), .Q (new_AGEMA_signal_3549) ) ;
    buf_clk new_AGEMA_reg_buffer_2101 ( .C (CLK), .D (new_AGEMA_signal_3552), .Q (new_AGEMA_signal_3553) ) ;
    buf_clk new_AGEMA_reg_buffer_2105 ( .C (CLK), .D (new_AGEMA_signal_3556), .Q (new_AGEMA_signal_3557) ) ;
    buf_clk new_AGEMA_reg_buffer_2109 ( .C (CLK), .D (new_AGEMA_signal_3560), .Q (new_AGEMA_signal_3561) ) ;
    buf_clk new_AGEMA_reg_buffer_2113 ( .C (CLK), .D (new_AGEMA_signal_3564), .Q (new_AGEMA_signal_3565) ) ;
    buf_clk new_AGEMA_reg_buffer_2117 ( .C (CLK), .D (new_AGEMA_signal_3568), .Q (new_AGEMA_signal_3569) ) ;
    buf_clk new_AGEMA_reg_buffer_2121 ( .C (CLK), .D (new_AGEMA_signal_3572), .Q (new_AGEMA_signal_3573) ) ;
    buf_clk new_AGEMA_reg_buffer_2125 ( .C (CLK), .D (new_AGEMA_signal_3576), .Q (new_AGEMA_signal_3577) ) ;
    buf_clk new_AGEMA_reg_buffer_2129 ( .C (CLK), .D (new_AGEMA_signal_3580), .Q (new_AGEMA_signal_3581) ) ;
    buf_clk new_AGEMA_reg_buffer_2133 ( .C (CLK), .D (new_AGEMA_signal_3584), .Q (new_AGEMA_signal_3585) ) ;
    buf_clk new_AGEMA_reg_buffer_2137 ( .C (CLK), .D (new_AGEMA_signal_3588), .Q (new_AGEMA_signal_3589) ) ;
    buf_clk new_AGEMA_reg_buffer_2141 ( .C (CLK), .D (new_AGEMA_signal_3592), .Q (new_AGEMA_signal_3593) ) ;
    buf_clk new_AGEMA_reg_buffer_2145 ( .C (CLK), .D (new_AGEMA_signal_3596), .Q (new_AGEMA_signal_3597) ) ;
    buf_clk new_AGEMA_reg_buffer_2149 ( .C (CLK), .D (new_AGEMA_signal_3600), .Q (new_AGEMA_signal_3601) ) ;
    buf_clk new_AGEMA_reg_buffer_2153 ( .C (CLK), .D (new_AGEMA_signal_3604), .Q (new_AGEMA_signal_3605) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (CLK), .D (new_AGEMA_signal_3608), .Q (new_AGEMA_signal_3609) ) ;
    buf_clk new_AGEMA_reg_buffer_2161 ( .C (CLK), .D (new_AGEMA_signal_3612), .Q (new_AGEMA_signal_3613) ) ;
    buf_clk new_AGEMA_reg_buffer_2165 ( .C (CLK), .D (new_AGEMA_signal_3616), .Q (new_AGEMA_signal_3617) ) ;
    buf_clk new_AGEMA_reg_buffer_2169 ( .C (CLK), .D (new_AGEMA_signal_3620), .Q (new_AGEMA_signal_3621) ) ;
    buf_clk new_AGEMA_reg_buffer_2173 ( .C (CLK), .D (new_AGEMA_signal_3624), .Q (new_AGEMA_signal_3625) ) ;
    buf_clk new_AGEMA_reg_buffer_2177 ( .C (CLK), .D (new_AGEMA_signal_3628), .Q (new_AGEMA_signal_3629) ) ;
    buf_clk new_AGEMA_reg_buffer_2181 ( .C (CLK), .D (new_AGEMA_signal_3632), .Q (new_AGEMA_signal_3633) ) ;
    buf_clk new_AGEMA_reg_buffer_2185 ( .C (CLK), .D (new_AGEMA_signal_3636), .Q (new_AGEMA_signal_3637) ) ;
    buf_clk new_AGEMA_reg_buffer_2189 ( .C (CLK), .D (new_AGEMA_signal_3640), .Q (new_AGEMA_signal_3641) ) ;
    buf_clk new_AGEMA_reg_buffer_2193 ( .C (CLK), .D (new_AGEMA_signal_3644), .Q (new_AGEMA_signal_3645) ) ;
    buf_clk new_AGEMA_reg_buffer_2197 ( .C (CLK), .D (new_AGEMA_signal_3648), .Q (new_AGEMA_signal_3649) ) ;
    buf_clk new_AGEMA_reg_buffer_2201 ( .C (CLK), .D (new_AGEMA_signal_3652), .Q (new_AGEMA_signal_3653) ) ;
    buf_clk new_AGEMA_reg_buffer_2205 ( .C (CLK), .D (new_AGEMA_signal_3656), .Q (new_AGEMA_signal_3657) ) ;
    buf_clk new_AGEMA_reg_buffer_2209 ( .C (CLK), .D (new_AGEMA_signal_3660), .Q (new_AGEMA_signal_3661) ) ;
    buf_clk new_AGEMA_reg_buffer_2213 ( .C (CLK), .D (new_AGEMA_signal_3664), .Q (new_AGEMA_signal_3665) ) ;
    buf_clk new_AGEMA_reg_buffer_2217 ( .C (CLK), .D (new_AGEMA_signal_3668), .Q (new_AGEMA_signal_3669) ) ;
    buf_clk new_AGEMA_reg_buffer_2221 ( .C (CLK), .D (new_AGEMA_signal_3672), .Q (new_AGEMA_signal_3673) ) ;
    buf_clk new_AGEMA_reg_buffer_2225 ( .C (CLK), .D (new_AGEMA_signal_3676), .Q (new_AGEMA_signal_3677) ) ;
    buf_clk new_AGEMA_reg_buffer_2229 ( .C (CLK), .D (new_AGEMA_signal_3680), .Q (new_AGEMA_signal_3681) ) ;
    buf_clk new_AGEMA_reg_buffer_2233 ( .C (CLK), .D (new_AGEMA_signal_3684), .Q (new_AGEMA_signal_3685) ) ;
    buf_clk new_AGEMA_reg_buffer_2237 ( .C (CLK), .D (new_AGEMA_signal_3688), .Q (new_AGEMA_signal_3689) ) ;
    buf_clk new_AGEMA_reg_buffer_2241 ( .C (CLK), .D (new_AGEMA_signal_3692), .Q (new_AGEMA_signal_3693) ) ;
    buf_clk new_AGEMA_reg_buffer_2245 ( .C (CLK), .D (new_AGEMA_signal_3696), .Q (new_AGEMA_signal_3697) ) ;
    buf_clk new_AGEMA_reg_buffer_2249 ( .C (CLK), .D (new_AGEMA_signal_3700), .Q (new_AGEMA_signal_3701) ) ;
    buf_clk new_AGEMA_reg_buffer_2253 ( .C (CLK), .D (new_AGEMA_signal_3704), .Q (new_AGEMA_signal_3705) ) ;
    buf_clk new_AGEMA_reg_buffer_2257 ( .C (CLK), .D (new_AGEMA_signal_3708), .Q (new_AGEMA_signal_3709) ) ;
    buf_clk new_AGEMA_reg_buffer_2261 ( .C (CLK), .D (new_AGEMA_signal_3712), .Q (new_AGEMA_signal_3713) ) ;
    buf_clk new_AGEMA_reg_buffer_2265 ( .C (CLK), .D (new_AGEMA_signal_3716), .Q (new_AGEMA_signal_3717) ) ;
    buf_clk new_AGEMA_reg_buffer_2269 ( .C (CLK), .D (new_AGEMA_signal_3720), .Q (new_AGEMA_signal_3721) ) ;
    buf_clk new_AGEMA_reg_buffer_2273 ( .C (CLK), .D (new_AGEMA_signal_3724), .Q (new_AGEMA_signal_3725) ) ;
    buf_clk new_AGEMA_reg_buffer_2277 ( .C (CLK), .D (new_AGEMA_signal_3728), .Q (new_AGEMA_signal_3729) ) ;
    buf_clk new_AGEMA_reg_buffer_2281 ( .C (CLK), .D (new_AGEMA_signal_3732), .Q (new_AGEMA_signal_3733) ) ;
    buf_clk new_AGEMA_reg_buffer_2285 ( .C (CLK), .D (new_AGEMA_signal_3736), .Q (new_AGEMA_signal_3737) ) ;
    buf_clk new_AGEMA_reg_buffer_2289 ( .C (CLK), .D (new_AGEMA_signal_3740), .Q (new_AGEMA_signal_3741) ) ;
    buf_clk new_AGEMA_reg_buffer_2293 ( .C (CLK), .D (new_AGEMA_signal_3744), .Q (new_AGEMA_signal_3745) ) ;
    buf_clk new_AGEMA_reg_buffer_2297 ( .C (CLK), .D (new_AGEMA_signal_3748), .Q (new_AGEMA_signal_3749) ) ;
    buf_clk new_AGEMA_reg_buffer_2301 ( .C (CLK), .D (new_AGEMA_signal_3752), .Q (new_AGEMA_signal_3753) ) ;
    buf_clk new_AGEMA_reg_buffer_2305 ( .C (CLK), .D (new_AGEMA_signal_3756), .Q (new_AGEMA_signal_3757) ) ;
    buf_clk new_AGEMA_reg_buffer_2309 ( .C (CLK), .D (new_AGEMA_signal_3760), .Q (new_AGEMA_signal_3761) ) ;
    buf_clk new_AGEMA_reg_buffer_2313 ( .C (CLK), .D (new_AGEMA_signal_3764), .Q (new_AGEMA_signal_3765) ) ;
    buf_clk new_AGEMA_reg_buffer_2317 ( .C (CLK), .D (new_AGEMA_signal_3768), .Q (new_AGEMA_signal_3769) ) ;
    buf_clk new_AGEMA_reg_buffer_2321 ( .C (CLK), .D (new_AGEMA_signal_3772), .Q (new_AGEMA_signal_3773) ) ;
    buf_clk new_AGEMA_reg_buffer_2325 ( .C (CLK), .D (new_AGEMA_signal_3776), .Q (new_AGEMA_signal_3777) ) ;
    buf_clk new_AGEMA_reg_buffer_2329 ( .C (CLK), .D (new_AGEMA_signal_3780), .Q (new_AGEMA_signal_3781) ) ;
    buf_clk new_AGEMA_reg_buffer_2333 ( .C (CLK), .D (new_AGEMA_signal_3784), .Q (new_AGEMA_signal_3785) ) ;
    buf_clk new_AGEMA_reg_buffer_2337 ( .C (CLK), .D (new_AGEMA_signal_3788), .Q (new_AGEMA_signal_3789) ) ;
    buf_clk new_AGEMA_reg_buffer_2341 ( .C (CLK), .D (new_AGEMA_signal_3792), .Q (new_AGEMA_signal_3793) ) ;
    buf_clk new_AGEMA_reg_buffer_2345 ( .C (CLK), .D (new_AGEMA_signal_3796), .Q (new_AGEMA_signal_3797) ) ;
    buf_clk new_AGEMA_reg_buffer_2349 ( .C (CLK), .D (new_AGEMA_signal_3800), .Q (new_AGEMA_signal_3801) ) ;
    buf_clk new_AGEMA_reg_buffer_2353 ( .C (CLK), .D (new_AGEMA_signal_3804), .Q (new_AGEMA_signal_3805) ) ;
    buf_clk new_AGEMA_reg_buffer_2357 ( .C (CLK), .D (new_AGEMA_signal_3808), .Q (new_AGEMA_signal_3809) ) ;
    buf_clk new_AGEMA_reg_buffer_2361 ( .C (CLK), .D (new_AGEMA_signal_3812), .Q (new_AGEMA_signal_3813) ) ;
    buf_clk new_AGEMA_reg_buffer_2365 ( .C (CLK), .D (new_AGEMA_signal_3816), .Q (new_AGEMA_signal_3817) ) ;
    buf_clk new_AGEMA_reg_buffer_2367 ( .C (CLK), .D (new_AGEMA_signal_3818), .Q (new_AGEMA_signal_3819) ) ;
    buf_clk new_AGEMA_reg_buffer_2369 ( .C (CLK), .D (new_AGEMA_signal_3820), .Q (new_AGEMA_signal_3821) ) ;
    buf_clk new_AGEMA_reg_buffer_2371 ( .C (CLK), .D (new_AGEMA_signal_3822), .Q (new_AGEMA_signal_3823) ) ;
    buf_clk new_AGEMA_reg_buffer_2377 ( .C (CLK), .D (new_AGEMA_signal_3828), .Q (new_AGEMA_signal_3829) ) ;
    buf_clk new_AGEMA_reg_buffer_2381 ( .C (CLK), .D (new_AGEMA_signal_3832), .Q (new_AGEMA_signal_3833) ) ;
    buf_clk new_AGEMA_reg_buffer_2385 ( .C (CLK), .D (new_AGEMA_signal_3836), .Q (new_AGEMA_signal_3837) ) ;
    buf_clk new_AGEMA_reg_buffer_2389 ( .C (CLK), .D (new_AGEMA_signal_3840), .Q (new_AGEMA_signal_3841) ) ;
    buf_clk new_AGEMA_reg_buffer_2397 ( .C (CLK), .D (new_AGEMA_signal_3848), .Q (new_AGEMA_signal_3849) ) ;
    buf_clk new_AGEMA_reg_buffer_2399 ( .C (CLK), .D (new_AGEMA_signal_3850), .Q (new_AGEMA_signal_3851) ) ;
    buf_clk new_AGEMA_reg_buffer_2401 ( .C (CLK), .D (new_AGEMA_signal_3852), .Q (new_AGEMA_signal_3853) ) ;
    buf_clk new_AGEMA_reg_buffer_2403 ( .C (CLK), .D (new_AGEMA_signal_3854), .Q (new_AGEMA_signal_3855) ) ;
    buf_clk new_AGEMA_reg_buffer_2409 ( .C (CLK), .D (new_AGEMA_signal_3860), .Q (new_AGEMA_signal_3861) ) ;
    buf_clk new_AGEMA_reg_buffer_2413 ( .C (CLK), .D (new_AGEMA_signal_3864), .Q (new_AGEMA_signal_3865) ) ;
    buf_clk new_AGEMA_reg_buffer_2417 ( .C (CLK), .D (new_AGEMA_signal_3868), .Q (new_AGEMA_signal_3869) ) ;
    buf_clk new_AGEMA_reg_buffer_2421 ( .C (CLK), .D (new_AGEMA_signal_3872), .Q (new_AGEMA_signal_3873) ) ;
    buf_clk new_AGEMA_reg_buffer_2429 ( .C (CLK), .D (new_AGEMA_signal_3880), .Q (new_AGEMA_signal_3881) ) ;
    buf_clk new_AGEMA_reg_buffer_2431 ( .C (CLK), .D (new_AGEMA_signal_3882), .Q (new_AGEMA_signal_3883) ) ;
    buf_clk new_AGEMA_reg_buffer_2433 ( .C (CLK), .D (new_AGEMA_signal_3884), .Q (new_AGEMA_signal_3885) ) ;
    buf_clk new_AGEMA_reg_buffer_2435 ( .C (CLK), .D (new_AGEMA_signal_3886), .Q (new_AGEMA_signal_3887) ) ;
    buf_clk new_AGEMA_reg_buffer_2441 ( .C (CLK), .D (new_AGEMA_signal_3892), .Q (new_AGEMA_signal_3893) ) ;
    buf_clk new_AGEMA_reg_buffer_2445 ( .C (CLK), .D (new_AGEMA_signal_3896), .Q (new_AGEMA_signal_3897) ) ;
    buf_clk new_AGEMA_reg_buffer_2453 ( .C (CLK), .D (new_AGEMA_signal_3904), .Q (new_AGEMA_signal_3905) ) ;
    buf_clk new_AGEMA_reg_buffer_2455 ( .C (CLK), .D (new_AGEMA_signal_3906), .Q (new_AGEMA_signal_3907) ) ;
    buf_clk new_AGEMA_reg_buffer_2457 ( .C (CLK), .D (new_AGEMA_signal_3908), .Q (new_AGEMA_signal_3909) ) ;
    buf_clk new_AGEMA_reg_buffer_2459 ( .C (CLK), .D (new_AGEMA_signal_3910), .Q (new_AGEMA_signal_3911) ) ;
    buf_clk new_AGEMA_reg_buffer_2465 ( .C (CLK), .D (new_AGEMA_signal_3916), .Q (new_AGEMA_signal_3917) ) ;
    buf_clk new_AGEMA_reg_buffer_2469 ( .C (CLK), .D (new_AGEMA_signal_3920), .Q (new_AGEMA_signal_3921) ) ;
    buf_clk new_AGEMA_reg_buffer_2477 ( .C (CLK), .D (new_AGEMA_signal_3928), .Q (new_AGEMA_signal_3929) ) ;
    buf_clk new_AGEMA_reg_buffer_2479 ( .C (CLK), .D (new_AGEMA_signal_3930), .Q (new_AGEMA_signal_3931) ) ;
    buf_clk new_AGEMA_reg_buffer_2481 ( .C (CLK), .D (new_AGEMA_signal_3932), .Q (new_AGEMA_signal_3933) ) ;
    buf_clk new_AGEMA_reg_buffer_2483 ( .C (CLK), .D (new_AGEMA_signal_3934), .Q (new_AGEMA_signal_3935) ) ;
    buf_clk new_AGEMA_reg_buffer_2489 ( .C (CLK), .D (new_AGEMA_signal_3940), .Q (new_AGEMA_signal_3941) ) ;
    buf_clk new_AGEMA_reg_buffer_2493 ( .C (CLK), .D (new_AGEMA_signal_3944), .Q (new_AGEMA_signal_3945) ) ;
    buf_clk new_AGEMA_reg_buffer_2497 ( .C (CLK), .D (new_AGEMA_signal_3948), .Q (new_AGEMA_signal_3949) ) ;
    buf_clk new_AGEMA_reg_buffer_2501 ( .C (CLK), .D (new_AGEMA_signal_3952), .Q (new_AGEMA_signal_3953) ) ;
    buf_clk new_AGEMA_reg_buffer_2509 ( .C (CLK), .D (new_AGEMA_signal_3960), .Q (new_AGEMA_signal_3961) ) ;
    buf_clk new_AGEMA_reg_buffer_2511 ( .C (CLK), .D (new_AGEMA_signal_3962), .Q (new_AGEMA_signal_3963) ) ;
    buf_clk new_AGEMA_reg_buffer_2513 ( .C (CLK), .D (new_AGEMA_signal_3964), .Q (new_AGEMA_signal_3965) ) ;
    buf_clk new_AGEMA_reg_buffer_2515 ( .C (CLK), .D (new_AGEMA_signal_3966), .Q (new_AGEMA_signal_3967) ) ;
    buf_clk new_AGEMA_reg_buffer_2521 ( .C (CLK), .D (new_AGEMA_signal_3972), .Q (new_AGEMA_signal_3973) ) ;
    buf_clk new_AGEMA_reg_buffer_2525 ( .C (CLK), .D (new_AGEMA_signal_3976), .Q (new_AGEMA_signal_3977) ) ;
    buf_clk new_AGEMA_reg_buffer_2529 ( .C (CLK), .D (new_AGEMA_signal_3980), .Q (new_AGEMA_signal_3981) ) ;
    buf_clk new_AGEMA_reg_buffer_2533 ( .C (CLK), .D (new_AGEMA_signal_3984), .Q (new_AGEMA_signal_3985) ) ;
    buf_clk new_AGEMA_reg_buffer_2541 ( .C (CLK), .D (new_AGEMA_signal_3992), .Q (new_AGEMA_signal_3993) ) ;
    buf_clk new_AGEMA_reg_buffer_2543 ( .C (CLK), .D (new_AGEMA_signal_3994), .Q (new_AGEMA_signal_3995) ) ;
    buf_clk new_AGEMA_reg_buffer_2545 ( .C (CLK), .D (new_AGEMA_signal_3996), .Q (new_AGEMA_signal_3997) ) ;
    buf_clk new_AGEMA_reg_buffer_2547 ( .C (CLK), .D (new_AGEMA_signal_3998), .Q (new_AGEMA_signal_3999) ) ;
    buf_clk new_AGEMA_reg_buffer_2553 ( .C (CLK), .D (new_AGEMA_signal_4004), .Q (new_AGEMA_signal_4005) ) ;
    buf_clk new_AGEMA_reg_buffer_2557 ( .C (CLK), .D (new_AGEMA_signal_4008), .Q (new_AGEMA_signal_4009) ) ;
    buf_clk new_AGEMA_reg_buffer_2565 ( .C (CLK), .D (new_AGEMA_signal_4016), .Q (new_AGEMA_signal_4017) ) ;
    buf_clk new_AGEMA_reg_buffer_2567 ( .C (CLK), .D (new_AGEMA_signal_4018), .Q (new_AGEMA_signal_4019) ) ;
    buf_clk new_AGEMA_reg_buffer_2569 ( .C (CLK), .D (new_AGEMA_signal_4020), .Q (new_AGEMA_signal_4021) ) ;
    buf_clk new_AGEMA_reg_buffer_2571 ( .C (CLK), .D (new_AGEMA_signal_4022), .Q (new_AGEMA_signal_4023) ) ;
    buf_clk new_AGEMA_reg_buffer_2577 ( .C (CLK), .D (new_AGEMA_signal_4028), .Q (new_AGEMA_signal_4029) ) ;
    buf_clk new_AGEMA_reg_buffer_2581 ( .C (CLK), .D (new_AGEMA_signal_4032), .Q (new_AGEMA_signal_4033) ) ;
    buf_clk new_AGEMA_reg_buffer_2589 ( .C (CLK), .D (new_AGEMA_signal_4040), .Q (new_AGEMA_signal_4041) ) ;
    buf_clk new_AGEMA_reg_buffer_2591 ( .C (CLK), .D (new_AGEMA_signal_4042), .Q (new_AGEMA_signal_4043) ) ;
    buf_clk new_AGEMA_reg_buffer_2593 ( .C (CLK), .D (new_AGEMA_signal_4044), .Q (new_AGEMA_signal_4045) ) ;
    buf_clk new_AGEMA_reg_buffer_2595 ( .C (CLK), .D (new_AGEMA_signal_4046), .Q (new_AGEMA_signal_4047) ) ;
    buf_clk new_AGEMA_reg_buffer_2601 ( .C (CLK), .D (new_AGEMA_signal_4052), .Q (new_AGEMA_signal_4053) ) ;
    buf_clk new_AGEMA_reg_buffer_2605 ( .C (CLK), .D (new_AGEMA_signal_4056), .Q (new_AGEMA_signal_4057) ) ;
    buf_clk new_AGEMA_reg_buffer_2609 ( .C (CLK), .D (new_AGEMA_signal_4060), .Q (new_AGEMA_signal_4061) ) ;
    buf_clk new_AGEMA_reg_buffer_2613 ( .C (CLK), .D (new_AGEMA_signal_4064), .Q (new_AGEMA_signal_4065) ) ;
    buf_clk new_AGEMA_reg_buffer_2621 ( .C (CLK), .D (new_AGEMA_signal_4072), .Q (new_AGEMA_signal_4073) ) ;
    buf_clk new_AGEMA_reg_buffer_2623 ( .C (CLK), .D (new_AGEMA_signal_4074), .Q (new_AGEMA_signal_4075) ) ;
    buf_clk new_AGEMA_reg_buffer_2625 ( .C (CLK), .D (new_AGEMA_signal_4076), .Q (new_AGEMA_signal_4077) ) ;
    buf_clk new_AGEMA_reg_buffer_2627 ( .C (CLK), .D (new_AGEMA_signal_4078), .Q (new_AGEMA_signal_4079) ) ;
    buf_clk new_AGEMA_reg_buffer_2633 ( .C (CLK), .D (new_AGEMA_signal_4084), .Q (new_AGEMA_signal_4085) ) ;
    buf_clk new_AGEMA_reg_buffer_2637 ( .C (CLK), .D (new_AGEMA_signal_4088), .Q (new_AGEMA_signal_4089) ) ;
    buf_clk new_AGEMA_reg_buffer_2641 ( .C (CLK), .D (new_AGEMA_signal_4092), .Q (new_AGEMA_signal_4093) ) ;
    buf_clk new_AGEMA_reg_buffer_2645 ( .C (CLK), .D (new_AGEMA_signal_4096), .Q (new_AGEMA_signal_4097) ) ;
    buf_clk new_AGEMA_reg_buffer_2653 ( .C (CLK), .D (new_AGEMA_signal_4104), .Q (new_AGEMA_signal_4105) ) ;
    buf_clk new_AGEMA_reg_buffer_2655 ( .C (CLK), .D (new_AGEMA_signal_4106), .Q (new_AGEMA_signal_4107) ) ;
    buf_clk new_AGEMA_reg_buffer_2657 ( .C (CLK), .D (new_AGEMA_signal_4108), .Q (new_AGEMA_signal_4109) ) ;
    buf_clk new_AGEMA_reg_buffer_2659 ( .C (CLK), .D (new_AGEMA_signal_4110), .Q (new_AGEMA_signal_4111) ) ;
    buf_clk new_AGEMA_reg_buffer_2665 ( .C (CLK), .D (new_AGEMA_signal_4116), .Q (new_AGEMA_signal_4117) ) ;
    buf_clk new_AGEMA_reg_buffer_2669 ( .C (CLK), .D (new_AGEMA_signal_4120), .Q (new_AGEMA_signal_4121) ) ;
    buf_clk new_AGEMA_reg_buffer_2677 ( .C (CLK), .D (new_AGEMA_signal_4128), .Q (new_AGEMA_signal_4129) ) ;
    buf_clk new_AGEMA_reg_buffer_2679 ( .C (CLK), .D (new_AGEMA_signal_4130), .Q (new_AGEMA_signal_4131) ) ;
    buf_clk new_AGEMA_reg_buffer_2681 ( .C (CLK), .D (new_AGEMA_signal_4132), .Q (new_AGEMA_signal_4133) ) ;
    buf_clk new_AGEMA_reg_buffer_2683 ( .C (CLK), .D (new_AGEMA_signal_4134), .Q (new_AGEMA_signal_4135) ) ;
    buf_clk new_AGEMA_reg_buffer_2689 ( .C (CLK), .D (new_AGEMA_signal_4140), .Q (new_AGEMA_signal_4141) ) ;
    buf_clk new_AGEMA_reg_buffer_2693 ( .C (CLK), .D (new_AGEMA_signal_4144), .Q (new_AGEMA_signal_4145) ) ;
    buf_clk new_AGEMA_reg_buffer_2701 ( .C (CLK), .D (new_AGEMA_signal_4152), .Q (new_AGEMA_signal_4153) ) ;
    buf_clk new_AGEMA_reg_buffer_2703 ( .C (CLK), .D (new_AGEMA_signal_4154), .Q (new_AGEMA_signal_4155) ) ;
    buf_clk new_AGEMA_reg_buffer_2705 ( .C (CLK), .D (new_AGEMA_signal_4156), .Q (new_AGEMA_signal_4157) ) ;
    buf_clk new_AGEMA_reg_buffer_2707 ( .C (CLK), .D (new_AGEMA_signal_4158), .Q (new_AGEMA_signal_4159) ) ;
    buf_clk new_AGEMA_reg_buffer_2713 ( .C (CLK), .D (new_AGEMA_signal_4164), .Q (new_AGEMA_signal_4165) ) ;
    buf_clk new_AGEMA_reg_buffer_2717 ( .C (CLK), .D (new_AGEMA_signal_4168), .Q (new_AGEMA_signal_4169) ) ;
    buf_clk new_AGEMA_reg_buffer_2721 ( .C (CLK), .D (new_AGEMA_signal_4172), .Q (new_AGEMA_signal_4173) ) ;
    buf_clk new_AGEMA_reg_buffer_2725 ( .C (CLK), .D (new_AGEMA_signal_4176), .Q (new_AGEMA_signal_4177) ) ;
    buf_clk new_AGEMA_reg_buffer_2733 ( .C (CLK), .D (new_AGEMA_signal_4184), .Q (new_AGEMA_signal_4185) ) ;
    buf_clk new_AGEMA_reg_buffer_2735 ( .C (CLK), .D (new_AGEMA_signal_4186), .Q (new_AGEMA_signal_4187) ) ;
    buf_clk new_AGEMA_reg_buffer_2737 ( .C (CLK), .D (new_AGEMA_signal_4188), .Q (new_AGEMA_signal_4189) ) ;
    buf_clk new_AGEMA_reg_buffer_2739 ( .C (CLK), .D (new_AGEMA_signal_4190), .Q (new_AGEMA_signal_4191) ) ;
    buf_clk new_AGEMA_reg_buffer_2745 ( .C (CLK), .D (new_AGEMA_signal_4196), .Q (new_AGEMA_signal_4197) ) ;
    buf_clk new_AGEMA_reg_buffer_2749 ( .C (CLK), .D (new_AGEMA_signal_4200), .Q (new_AGEMA_signal_4201) ) ;
    buf_clk new_AGEMA_reg_buffer_2753 ( .C (CLK), .D (new_AGEMA_signal_4204), .Q (new_AGEMA_signal_4205) ) ;
    buf_clk new_AGEMA_reg_buffer_2757 ( .C (CLK), .D (new_AGEMA_signal_4208), .Q (new_AGEMA_signal_4209) ) ;
    buf_clk new_AGEMA_reg_buffer_2765 ( .C (CLK), .D (new_AGEMA_signal_4216), .Q (new_AGEMA_signal_4217) ) ;
    buf_clk new_AGEMA_reg_buffer_2767 ( .C (CLK), .D (new_AGEMA_signal_4218), .Q (new_AGEMA_signal_4219) ) ;
    buf_clk new_AGEMA_reg_buffer_2769 ( .C (CLK), .D (new_AGEMA_signal_4220), .Q (new_AGEMA_signal_4221) ) ;
    buf_clk new_AGEMA_reg_buffer_2771 ( .C (CLK), .D (new_AGEMA_signal_4222), .Q (new_AGEMA_signal_4223) ) ;
    buf_clk new_AGEMA_reg_buffer_2777 ( .C (CLK), .D (new_AGEMA_signal_4228), .Q (new_AGEMA_signal_4229) ) ;
    buf_clk new_AGEMA_reg_buffer_2781 ( .C (CLK), .D (new_AGEMA_signal_4232), .Q (new_AGEMA_signal_4233) ) ;
    buf_clk new_AGEMA_reg_buffer_2789 ( .C (CLK), .D (new_AGEMA_signal_4240), .Q (new_AGEMA_signal_4241) ) ;
    buf_clk new_AGEMA_reg_buffer_2791 ( .C (CLK), .D (new_AGEMA_signal_4242), .Q (new_AGEMA_signal_4243) ) ;
    buf_clk new_AGEMA_reg_buffer_2793 ( .C (CLK), .D (new_AGEMA_signal_4244), .Q (new_AGEMA_signal_4245) ) ;
    buf_clk new_AGEMA_reg_buffer_2795 ( .C (CLK), .D (new_AGEMA_signal_4246), .Q (new_AGEMA_signal_4247) ) ;
    buf_clk new_AGEMA_reg_buffer_2801 ( .C (CLK), .D (new_AGEMA_signal_4252), .Q (new_AGEMA_signal_4253) ) ;
    buf_clk new_AGEMA_reg_buffer_2805 ( .C (CLK), .D (new_AGEMA_signal_4256), .Q (new_AGEMA_signal_4257) ) ;
    buf_clk new_AGEMA_reg_buffer_2877 ( .C (CLK), .D (new_AGEMA_signal_4328), .Q (new_AGEMA_signal_4329) ) ;
    buf_clk new_AGEMA_reg_buffer_2881 ( .C (CLK), .D (new_AGEMA_signal_4332), .Q (new_AGEMA_signal_4333) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (CLK), .D (new_AGEMA_signal_4336), .Q (new_AGEMA_signal_4337) ) ;
    buf_clk new_AGEMA_reg_buffer_2889 ( .C (CLK), .D (new_AGEMA_signal_4340), .Q (new_AGEMA_signal_4341) ) ;
    buf_clk new_AGEMA_reg_buffer_2893 ( .C (CLK), .D (new_AGEMA_signal_4344), .Q (new_AGEMA_signal_4345) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (CLK), .D (new_AGEMA_signal_4348), .Q (new_AGEMA_signal_4349) ) ;
    buf_clk new_AGEMA_reg_buffer_2901 ( .C (CLK), .D (new_AGEMA_signal_4352), .Q (new_AGEMA_signal_4353) ) ;
    buf_clk new_AGEMA_reg_buffer_2905 ( .C (CLK), .D (new_AGEMA_signal_4356), .Q (new_AGEMA_signal_4357) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (CLK), .D (new_AGEMA_signal_4360), .Q (new_AGEMA_signal_4361) ) ;
    buf_clk new_AGEMA_reg_buffer_2913 ( .C (CLK), .D (new_AGEMA_signal_4364), .Q (new_AGEMA_signal_4365) ) ;
    buf_clk new_AGEMA_reg_buffer_2917 ( .C (CLK), .D (new_AGEMA_signal_4368), .Q (new_AGEMA_signal_4369) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (CLK), .D (new_AGEMA_signal_2773), .Q (new_AGEMA_signal_2774) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (CLK), .D (new_AGEMA_signal_2777), .Q (new_AGEMA_signal_2778) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (CLK), .D (new_AGEMA_signal_2781), .Q (new_AGEMA_signal_2782) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (CLK), .D (new_AGEMA_signal_2785), .Q (new_AGEMA_signal_2786) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (CLK), .D (new_AGEMA_signal_2789), .Q (new_AGEMA_signal_2790) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (CLK), .D (new_AGEMA_signal_2793), .Q (new_AGEMA_signal_2794) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (CLK), .D (new_AGEMA_signal_2797), .Q (new_AGEMA_signal_2798) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (CLK), .D (new_AGEMA_signal_2801), .Q (new_AGEMA_signal_2802) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (CLK), .D (new_AGEMA_signal_2805), .Q (new_AGEMA_signal_2806) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (CLK), .D (new_AGEMA_signal_2809), .Q (new_AGEMA_signal_2810) ) ;
    buf_clk new_AGEMA_reg_buffer_1362 ( .C (CLK), .D (new_AGEMA_signal_2813), .Q (new_AGEMA_signal_2814) ) ;
    buf_clk new_AGEMA_reg_buffer_1366 ( .C (CLK), .D (new_AGEMA_signal_2817), .Q (new_AGEMA_signal_2818) ) ;
    buf_clk new_AGEMA_reg_buffer_1370 ( .C (CLK), .D (new_AGEMA_signal_2821), .Q (new_AGEMA_signal_2822) ) ;
    buf_clk new_AGEMA_reg_buffer_1374 ( .C (CLK), .D (new_AGEMA_signal_2825), .Q (new_AGEMA_signal_2826) ) ;
    buf_clk new_AGEMA_reg_buffer_1378 ( .C (CLK), .D (new_AGEMA_signal_2829), .Q (new_AGEMA_signal_2830) ) ;
    buf_clk new_AGEMA_reg_buffer_1382 ( .C (CLK), .D (new_AGEMA_signal_2833), .Q (new_AGEMA_signal_2834) ) ;
    buf_clk new_AGEMA_reg_buffer_1386 ( .C (CLK), .D (new_AGEMA_signal_2837), .Q (new_AGEMA_signal_2838) ) ;
    buf_clk new_AGEMA_reg_buffer_1390 ( .C (CLK), .D (new_AGEMA_signal_2841), .Q (new_AGEMA_signal_2842) ) ;
    buf_clk new_AGEMA_reg_buffer_1394 ( .C (CLK), .D (new_AGEMA_signal_2845), .Q (new_AGEMA_signal_2846) ) ;
    buf_clk new_AGEMA_reg_buffer_1398 ( .C (CLK), .D (new_AGEMA_signal_2849), .Q (new_AGEMA_signal_2850) ) ;
    buf_clk new_AGEMA_reg_buffer_1402 ( .C (CLK), .D (new_AGEMA_signal_2853), .Q (new_AGEMA_signal_2854) ) ;
    buf_clk new_AGEMA_reg_buffer_1406 ( .C (CLK), .D (new_AGEMA_signal_2857), .Q (new_AGEMA_signal_2858) ) ;
    buf_clk new_AGEMA_reg_buffer_1410 ( .C (CLK), .D (new_AGEMA_signal_2861), .Q (new_AGEMA_signal_2862) ) ;
    buf_clk new_AGEMA_reg_buffer_1414 ( .C (CLK), .D (new_AGEMA_signal_2865), .Q (new_AGEMA_signal_2866) ) ;
    buf_clk new_AGEMA_reg_buffer_1418 ( .C (CLK), .D (new_AGEMA_signal_2869), .Q (new_AGEMA_signal_2870) ) ;
    buf_clk new_AGEMA_reg_buffer_1422 ( .C (CLK), .D (new_AGEMA_signal_2873), .Q (new_AGEMA_signal_2874) ) ;
    buf_clk new_AGEMA_reg_buffer_1426 ( .C (CLK), .D (new_AGEMA_signal_2877), .Q (new_AGEMA_signal_2878) ) ;
    buf_clk new_AGEMA_reg_buffer_1430 ( .C (CLK), .D (new_AGEMA_signal_2881), .Q (new_AGEMA_signal_2882) ) ;
    buf_clk new_AGEMA_reg_buffer_1434 ( .C (CLK), .D (new_AGEMA_signal_2885), .Q (new_AGEMA_signal_2886) ) ;
    buf_clk new_AGEMA_reg_buffer_1438 ( .C (CLK), .D (new_AGEMA_signal_2889), .Q (new_AGEMA_signal_2890) ) ;
    buf_clk new_AGEMA_reg_buffer_1442 ( .C (CLK), .D (new_AGEMA_signal_2893), .Q (new_AGEMA_signal_2894) ) ;
    buf_clk new_AGEMA_reg_buffer_1446 ( .C (CLK), .D (new_AGEMA_signal_2897), .Q (new_AGEMA_signal_2898) ) ;
    buf_clk new_AGEMA_reg_buffer_1450 ( .C (CLK), .D (new_AGEMA_signal_2901), .Q (new_AGEMA_signal_2902) ) ;
    buf_clk new_AGEMA_reg_buffer_1454 ( .C (CLK), .D (new_AGEMA_signal_2905), .Q (new_AGEMA_signal_2906) ) ;
    buf_clk new_AGEMA_reg_buffer_1458 ( .C (CLK), .D (new_AGEMA_signal_2909), .Q (new_AGEMA_signal_2910) ) ;
    buf_clk new_AGEMA_reg_buffer_1462 ( .C (CLK), .D (new_AGEMA_signal_2913), .Q (new_AGEMA_signal_2914) ) ;
    buf_clk new_AGEMA_reg_buffer_1466 ( .C (CLK), .D (new_AGEMA_signal_2917), .Q (new_AGEMA_signal_2918) ) ;
    buf_clk new_AGEMA_reg_buffer_1470 ( .C (CLK), .D (new_AGEMA_signal_2921), .Q (new_AGEMA_signal_2922) ) ;
    buf_clk new_AGEMA_reg_buffer_1474 ( .C (CLK), .D (new_AGEMA_signal_2925), .Q (new_AGEMA_signal_2926) ) ;
    buf_clk new_AGEMA_reg_buffer_1478 ( .C (CLK), .D (new_AGEMA_signal_2929), .Q (new_AGEMA_signal_2930) ) ;
    buf_clk new_AGEMA_reg_buffer_1482 ( .C (CLK), .D (new_AGEMA_signal_2933), .Q (new_AGEMA_signal_2934) ) ;
    buf_clk new_AGEMA_reg_buffer_1486 ( .C (CLK), .D (new_AGEMA_signal_2937), .Q (new_AGEMA_signal_2938) ) ;
    buf_clk new_AGEMA_reg_buffer_1490 ( .C (CLK), .D (new_AGEMA_signal_2941), .Q (new_AGEMA_signal_2942) ) ;
    buf_clk new_AGEMA_reg_buffer_1494 ( .C (CLK), .D (new_AGEMA_signal_2945), .Q (new_AGEMA_signal_2946) ) ;
    buf_clk new_AGEMA_reg_buffer_1498 ( .C (CLK), .D (new_AGEMA_signal_2949), .Q (new_AGEMA_signal_2950) ) ;
    buf_clk new_AGEMA_reg_buffer_1502 ( .C (CLK), .D (new_AGEMA_signal_2953), .Q (new_AGEMA_signal_2954) ) ;
    buf_clk new_AGEMA_reg_buffer_1506 ( .C (CLK), .D (new_AGEMA_signal_2957), .Q (new_AGEMA_signal_2958) ) ;
    buf_clk new_AGEMA_reg_buffer_1510 ( .C (CLK), .D (new_AGEMA_signal_2961), .Q (new_AGEMA_signal_2962) ) ;
    buf_clk new_AGEMA_reg_buffer_1514 ( .C (CLK), .D (new_AGEMA_signal_2965), .Q (new_AGEMA_signal_2966) ) ;
    buf_clk new_AGEMA_reg_buffer_1518 ( .C (CLK), .D (new_AGEMA_signal_2969), .Q (new_AGEMA_signal_2970) ) ;
    buf_clk new_AGEMA_reg_buffer_1522 ( .C (CLK), .D (new_AGEMA_signal_2973), .Q (new_AGEMA_signal_2974) ) ;
    buf_clk new_AGEMA_reg_buffer_1526 ( .C (CLK), .D (new_AGEMA_signal_2977), .Q (new_AGEMA_signal_2978) ) ;
    buf_clk new_AGEMA_reg_buffer_1530 ( .C (CLK), .D (new_AGEMA_signal_2981), .Q (new_AGEMA_signal_2982) ) ;
    buf_clk new_AGEMA_reg_buffer_1534 ( .C (CLK), .D (new_AGEMA_signal_2985), .Q (new_AGEMA_signal_2986) ) ;
    buf_clk new_AGEMA_reg_buffer_1538 ( .C (CLK), .D (new_AGEMA_signal_2989), .Q (new_AGEMA_signal_2990) ) ;
    buf_clk new_AGEMA_reg_buffer_1542 ( .C (CLK), .D (new_AGEMA_signal_2993), .Q (new_AGEMA_signal_2994) ) ;
    buf_clk new_AGEMA_reg_buffer_1546 ( .C (CLK), .D (new_AGEMA_signal_2997), .Q (new_AGEMA_signal_2998) ) ;
    buf_clk new_AGEMA_reg_buffer_1550 ( .C (CLK), .D (new_AGEMA_signal_3001), .Q (new_AGEMA_signal_3002) ) ;
    buf_clk new_AGEMA_reg_buffer_1554 ( .C (CLK), .D (new_AGEMA_signal_3005), .Q (new_AGEMA_signal_3006) ) ;
    buf_clk new_AGEMA_reg_buffer_1558 ( .C (CLK), .D (new_AGEMA_signal_3009), .Q (new_AGEMA_signal_3010) ) ;
    buf_clk new_AGEMA_reg_buffer_1562 ( .C (CLK), .D (new_AGEMA_signal_3013), .Q (new_AGEMA_signal_3014) ) ;
    buf_clk new_AGEMA_reg_buffer_1566 ( .C (CLK), .D (new_AGEMA_signal_3017), .Q (new_AGEMA_signal_3018) ) ;
    buf_clk new_AGEMA_reg_buffer_1570 ( .C (CLK), .D (new_AGEMA_signal_3021), .Q (new_AGEMA_signal_3022) ) ;
    buf_clk new_AGEMA_reg_buffer_1574 ( .C (CLK), .D (new_AGEMA_signal_3025), .Q (new_AGEMA_signal_3026) ) ;
    buf_clk new_AGEMA_reg_buffer_1578 ( .C (CLK), .D (new_AGEMA_signal_3029), .Q (new_AGEMA_signal_3030) ) ;
    buf_clk new_AGEMA_reg_buffer_1582 ( .C (CLK), .D (new_AGEMA_signal_3033), .Q (new_AGEMA_signal_3034) ) ;
    buf_clk new_AGEMA_reg_buffer_1586 ( .C (CLK), .D (new_AGEMA_signal_3037), .Q (new_AGEMA_signal_3038) ) ;
    buf_clk new_AGEMA_reg_buffer_1590 ( .C (CLK), .D (new_AGEMA_signal_3041), .Q (new_AGEMA_signal_3042) ) ;
    buf_clk new_AGEMA_reg_buffer_1594 ( .C (CLK), .D (new_AGEMA_signal_3045), .Q (new_AGEMA_signal_3046) ) ;
    buf_clk new_AGEMA_reg_buffer_1598 ( .C (CLK), .D (new_AGEMA_signal_3049), .Q (new_AGEMA_signal_3050) ) ;
    buf_clk new_AGEMA_reg_buffer_1602 ( .C (CLK), .D (new_AGEMA_signal_3053), .Q (new_AGEMA_signal_3054) ) ;
    buf_clk new_AGEMA_reg_buffer_1606 ( .C (CLK), .D (new_AGEMA_signal_3057), .Q (new_AGEMA_signal_3058) ) ;
    buf_clk new_AGEMA_reg_buffer_1610 ( .C (CLK), .D (new_AGEMA_signal_3061), .Q (new_AGEMA_signal_3062) ) ;
    buf_clk new_AGEMA_reg_buffer_1614 ( .C (CLK), .D (new_AGEMA_signal_3065), .Q (new_AGEMA_signal_3066) ) ;
    buf_clk new_AGEMA_reg_buffer_1618 ( .C (CLK), .D (new_AGEMA_signal_3069), .Q (new_AGEMA_signal_3070) ) ;
    buf_clk new_AGEMA_reg_buffer_1622 ( .C (CLK), .D (new_AGEMA_signal_3073), .Q (new_AGEMA_signal_3074) ) ;
    buf_clk new_AGEMA_reg_buffer_1626 ( .C (CLK), .D (new_AGEMA_signal_3077), .Q (new_AGEMA_signal_3078) ) ;
    buf_clk new_AGEMA_reg_buffer_1630 ( .C (CLK), .D (new_AGEMA_signal_3081), .Q (new_AGEMA_signal_3082) ) ;
    buf_clk new_AGEMA_reg_buffer_1634 ( .C (CLK), .D (new_AGEMA_signal_3085), .Q (new_AGEMA_signal_3086) ) ;
    buf_clk new_AGEMA_reg_buffer_1638 ( .C (CLK), .D (new_AGEMA_signal_3089), .Q (new_AGEMA_signal_3090) ) ;
    buf_clk new_AGEMA_reg_buffer_1642 ( .C (CLK), .D (new_AGEMA_signal_3093), .Q (new_AGEMA_signal_3094) ) ;
    buf_clk new_AGEMA_reg_buffer_1646 ( .C (CLK), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_3098) ) ;
    buf_clk new_AGEMA_reg_buffer_1650 ( .C (CLK), .D (new_AGEMA_signal_3101), .Q (new_AGEMA_signal_3102) ) ;
    buf_clk new_AGEMA_reg_buffer_1654 ( .C (CLK), .D (new_AGEMA_signal_3105), .Q (new_AGEMA_signal_3106) ) ;
    buf_clk new_AGEMA_reg_buffer_1658 ( .C (CLK), .D (new_AGEMA_signal_3109), .Q (new_AGEMA_signal_3110) ) ;
    buf_clk new_AGEMA_reg_buffer_1662 ( .C (CLK), .D (new_AGEMA_signal_3113), .Q (new_AGEMA_signal_3114) ) ;
    buf_clk new_AGEMA_reg_buffer_1666 ( .C (CLK), .D (new_AGEMA_signal_3117), .Q (new_AGEMA_signal_3118) ) ;
    buf_clk new_AGEMA_reg_buffer_1670 ( .C (CLK), .D (new_AGEMA_signal_3121), .Q (new_AGEMA_signal_3122) ) ;
    buf_clk new_AGEMA_reg_buffer_1674 ( .C (CLK), .D (new_AGEMA_signal_3125), .Q (new_AGEMA_signal_3126) ) ;
    buf_clk new_AGEMA_reg_buffer_1678 ( .C (CLK), .D (new_AGEMA_signal_3129), .Q (new_AGEMA_signal_3130) ) ;
    buf_clk new_AGEMA_reg_buffer_1682 ( .C (CLK), .D (new_AGEMA_signal_3133), .Q (new_AGEMA_signal_3134) ) ;
    buf_clk new_AGEMA_reg_buffer_1686 ( .C (CLK), .D (new_AGEMA_signal_3137), .Q (new_AGEMA_signal_3138) ) ;
    buf_clk new_AGEMA_reg_buffer_1690 ( .C (CLK), .D (new_AGEMA_signal_3141), .Q (new_AGEMA_signal_3142) ) ;
    buf_clk new_AGEMA_reg_buffer_1694 ( .C (CLK), .D (new_AGEMA_signal_3145), .Q (new_AGEMA_signal_3146) ) ;
    buf_clk new_AGEMA_reg_buffer_1698 ( .C (CLK), .D (new_AGEMA_signal_3149), .Q (new_AGEMA_signal_3150) ) ;
    buf_clk new_AGEMA_reg_buffer_1702 ( .C (CLK), .D (new_AGEMA_signal_3153), .Q (new_AGEMA_signal_3154) ) ;
    buf_clk new_AGEMA_reg_buffer_1706 ( .C (CLK), .D (new_AGEMA_signal_3157), .Q (new_AGEMA_signal_3158) ) ;
    buf_clk new_AGEMA_reg_buffer_1710 ( .C (CLK), .D (new_AGEMA_signal_3161), .Q (new_AGEMA_signal_3162) ) ;
    buf_clk new_AGEMA_reg_buffer_1714 ( .C (CLK), .D (new_AGEMA_signal_3165), .Q (new_AGEMA_signal_3166) ) ;
    buf_clk new_AGEMA_reg_buffer_1718 ( .C (CLK), .D (new_AGEMA_signal_3169), .Q (new_AGEMA_signal_3170) ) ;
    buf_clk new_AGEMA_reg_buffer_1722 ( .C (CLK), .D (new_AGEMA_signal_3173), .Q (new_AGEMA_signal_3174) ) ;
    buf_clk new_AGEMA_reg_buffer_1726 ( .C (CLK), .D (new_AGEMA_signal_3177), .Q (new_AGEMA_signal_3178) ) ;
    buf_clk new_AGEMA_reg_buffer_1730 ( .C (CLK), .D (new_AGEMA_signal_3181), .Q (new_AGEMA_signal_3182) ) ;
    buf_clk new_AGEMA_reg_buffer_1734 ( .C (CLK), .D (new_AGEMA_signal_3185), .Q (new_AGEMA_signal_3186) ) ;
    buf_clk new_AGEMA_reg_buffer_1738 ( .C (CLK), .D (new_AGEMA_signal_3189), .Q (new_AGEMA_signal_3190) ) ;
    buf_clk new_AGEMA_reg_buffer_1742 ( .C (CLK), .D (new_AGEMA_signal_3193), .Q (new_AGEMA_signal_3194) ) ;
    buf_clk new_AGEMA_reg_buffer_1746 ( .C (CLK), .D (new_AGEMA_signal_3197), .Q (new_AGEMA_signal_3198) ) ;
    buf_clk new_AGEMA_reg_buffer_1750 ( .C (CLK), .D (new_AGEMA_signal_3201), .Q (new_AGEMA_signal_3202) ) ;
    buf_clk new_AGEMA_reg_buffer_1754 ( .C (CLK), .D (new_AGEMA_signal_3205), .Q (new_AGEMA_signal_3206) ) ;
    buf_clk new_AGEMA_reg_buffer_1758 ( .C (CLK), .D (new_AGEMA_signal_3209), .Q (new_AGEMA_signal_3210) ) ;
    buf_clk new_AGEMA_reg_buffer_1762 ( .C (CLK), .D (new_AGEMA_signal_3213), .Q (new_AGEMA_signal_3214) ) ;
    buf_clk new_AGEMA_reg_buffer_1766 ( .C (CLK), .D (new_AGEMA_signal_3217), .Q (new_AGEMA_signal_3218) ) ;
    buf_clk new_AGEMA_reg_buffer_1770 ( .C (CLK), .D (new_AGEMA_signal_3221), .Q (new_AGEMA_signal_3222) ) ;
    buf_clk new_AGEMA_reg_buffer_1774 ( .C (CLK), .D (new_AGEMA_signal_3225), .Q (new_AGEMA_signal_3226) ) ;
    buf_clk new_AGEMA_reg_buffer_1778 ( .C (CLK), .D (new_AGEMA_signal_3229), .Q (new_AGEMA_signal_3230) ) ;
    buf_clk new_AGEMA_reg_buffer_1782 ( .C (CLK), .D (new_AGEMA_signal_3233), .Q (new_AGEMA_signal_3234) ) ;
    buf_clk new_AGEMA_reg_buffer_1786 ( .C (CLK), .D (new_AGEMA_signal_3237), .Q (new_AGEMA_signal_3238) ) ;
    buf_clk new_AGEMA_reg_buffer_1790 ( .C (CLK), .D (new_AGEMA_signal_3241), .Q (new_AGEMA_signal_3242) ) ;
    buf_clk new_AGEMA_reg_buffer_1794 ( .C (CLK), .D (new_AGEMA_signal_3245), .Q (new_AGEMA_signal_3246) ) ;
    buf_clk new_AGEMA_reg_buffer_1798 ( .C (CLK), .D (new_AGEMA_signal_3249), .Q (new_AGEMA_signal_3250) ) ;
    buf_clk new_AGEMA_reg_buffer_1802 ( .C (CLK), .D (new_AGEMA_signal_3253), .Q (new_AGEMA_signal_3254) ) ;
    buf_clk new_AGEMA_reg_buffer_1806 ( .C (CLK), .D (new_AGEMA_signal_3257), .Q (new_AGEMA_signal_3258) ) ;
    buf_clk new_AGEMA_reg_buffer_1810 ( .C (CLK), .D (new_AGEMA_signal_3261), .Q (new_AGEMA_signal_3262) ) ;
    buf_clk new_AGEMA_reg_buffer_1814 ( .C (CLK), .D (new_AGEMA_signal_3265), .Q (new_AGEMA_signal_3266) ) ;
    buf_clk new_AGEMA_reg_buffer_1818 ( .C (CLK), .D (new_AGEMA_signal_3269), .Q (new_AGEMA_signal_3270) ) ;
    buf_clk new_AGEMA_reg_buffer_1822 ( .C (CLK), .D (new_AGEMA_signal_3273), .Q (new_AGEMA_signal_3274) ) ;
    buf_clk new_AGEMA_reg_buffer_1826 ( .C (CLK), .D (new_AGEMA_signal_3277), .Q (new_AGEMA_signal_3278) ) ;
    buf_clk new_AGEMA_reg_buffer_1830 ( .C (CLK), .D (new_AGEMA_signal_3281), .Q (new_AGEMA_signal_3282) ) ;
    buf_clk new_AGEMA_reg_buffer_1834 ( .C (CLK), .D (new_AGEMA_signal_3285), .Q (new_AGEMA_signal_3286) ) ;
    buf_clk new_AGEMA_reg_buffer_1838 ( .C (CLK), .D (new_AGEMA_signal_3289), .Q (new_AGEMA_signal_3290) ) ;
    buf_clk new_AGEMA_reg_buffer_1842 ( .C (CLK), .D (new_AGEMA_signal_3293), .Q (new_AGEMA_signal_3294) ) ;
    buf_clk new_AGEMA_reg_buffer_1846 ( .C (CLK), .D (new_AGEMA_signal_3297), .Q (new_AGEMA_signal_3298) ) ;
    buf_clk new_AGEMA_reg_buffer_1850 ( .C (CLK), .D (new_AGEMA_signal_3301), .Q (new_AGEMA_signal_3302) ) ;
    buf_clk new_AGEMA_reg_buffer_1854 ( .C (CLK), .D (new_AGEMA_signal_3305), .Q (new_AGEMA_signal_3306) ) ;
    buf_clk new_AGEMA_reg_buffer_1858 ( .C (CLK), .D (new_AGEMA_signal_3309), .Q (new_AGEMA_signal_3310) ) ;
    buf_clk new_AGEMA_reg_buffer_1862 ( .C (CLK), .D (new_AGEMA_signal_3313), .Q (new_AGEMA_signal_3314) ) ;
    buf_clk new_AGEMA_reg_buffer_1866 ( .C (CLK), .D (new_AGEMA_signal_3317), .Q (new_AGEMA_signal_3318) ) ;
    buf_clk new_AGEMA_reg_buffer_1870 ( .C (CLK), .D (new_AGEMA_signal_3321), .Q (new_AGEMA_signal_3322) ) ;
    buf_clk new_AGEMA_reg_buffer_1874 ( .C (CLK), .D (new_AGEMA_signal_3325), .Q (new_AGEMA_signal_3326) ) ;
    buf_clk new_AGEMA_reg_buffer_1878 ( .C (CLK), .D (new_AGEMA_signal_3329), .Q (new_AGEMA_signal_3330) ) ;
    buf_clk new_AGEMA_reg_buffer_1882 ( .C (CLK), .D (new_AGEMA_signal_3333), .Q (new_AGEMA_signal_3334) ) ;
    buf_clk new_AGEMA_reg_buffer_1886 ( .C (CLK), .D (new_AGEMA_signal_3337), .Q (new_AGEMA_signal_3338) ) ;
    buf_clk new_AGEMA_reg_buffer_1890 ( .C (CLK), .D (new_AGEMA_signal_3341), .Q (new_AGEMA_signal_3342) ) ;
    buf_clk new_AGEMA_reg_buffer_1894 ( .C (CLK), .D (new_AGEMA_signal_3345), .Q (new_AGEMA_signal_3346) ) ;
    buf_clk new_AGEMA_reg_buffer_1898 ( .C (CLK), .D (new_AGEMA_signal_3349), .Q (new_AGEMA_signal_3350) ) ;
    buf_clk new_AGEMA_reg_buffer_1902 ( .C (CLK), .D (new_AGEMA_signal_3353), .Q (new_AGEMA_signal_3354) ) ;
    buf_clk new_AGEMA_reg_buffer_1906 ( .C (CLK), .D (new_AGEMA_signal_3357), .Q (new_AGEMA_signal_3358) ) ;
    buf_clk new_AGEMA_reg_buffer_1910 ( .C (CLK), .D (new_AGEMA_signal_3361), .Q (new_AGEMA_signal_3362) ) ;
    buf_clk new_AGEMA_reg_buffer_1914 ( .C (CLK), .D (new_AGEMA_signal_3365), .Q (new_AGEMA_signal_3366) ) ;
    buf_clk new_AGEMA_reg_buffer_1918 ( .C (CLK), .D (new_AGEMA_signal_3369), .Q (new_AGEMA_signal_3370) ) ;
    buf_clk new_AGEMA_reg_buffer_1922 ( .C (CLK), .D (new_AGEMA_signal_3373), .Q (new_AGEMA_signal_3374) ) ;
    buf_clk new_AGEMA_reg_buffer_1926 ( .C (CLK), .D (new_AGEMA_signal_3377), .Q (new_AGEMA_signal_3378) ) ;
    buf_clk new_AGEMA_reg_buffer_1930 ( .C (CLK), .D (new_AGEMA_signal_3381), .Q (new_AGEMA_signal_3382) ) ;
    buf_clk new_AGEMA_reg_buffer_1934 ( .C (CLK), .D (new_AGEMA_signal_3385), .Q (new_AGEMA_signal_3386) ) ;
    buf_clk new_AGEMA_reg_buffer_1938 ( .C (CLK), .D (new_AGEMA_signal_3389), .Q (new_AGEMA_signal_3390) ) ;
    buf_clk new_AGEMA_reg_buffer_1942 ( .C (CLK), .D (new_AGEMA_signal_3393), .Q (new_AGEMA_signal_3394) ) ;
    buf_clk new_AGEMA_reg_buffer_1946 ( .C (CLK), .D (new_AGEMA_signal_3397), .Q (new_AGEMA_signal_3398) ) ;
    buf_clk new_AGEMA_reg_buffer_1950 ( .C (CLK), .D (new_AGEMA_signal_3401), .Q (new_AGEMA_signal_3402) ) ;
    buf_clk new_AGEMA_reg_buffer_1954 ( .C (CLK), .D (new_AGEMA_signal_3405), .Q (new_AGEMA_signal_3406) ) ;
    buf_clk new_AGEMA_reg_buffer_1958 ( .C (CLK), .D (new_AGEMA_signal_3409), .Q (new_AGEMA_signal_3410) ) ;
    buf_clk new_AGEMA_reg_buffer_1962 ( .C (CLK), .D (new_AGEMA_signal_3413), .Q (new_AGEMA_signal_3414) ) ;
    buf_clk new_AGEMA_reg_buffer_1966 ( .C (CLK), .D (new_AGEMA_signal_3417), .Q (new_AGEMA_signal_3418) ) ;
    buf_clk new_AGEMA_reg_buffer_1970 ( .C (CLK), .D (new_AGEMA_signal_3421), .Q (new_AGEMA_signal_3422) ) ;
    buf_clk new_AGEMA_reg_buffer_1974 ( .C (CLK), .D (new_AGEMA_signal_3425), .Q (new_AGEMA_signal_3426) ) ;
    buf_clk new_AGEMA_reg_buffer_1978 ( .C (CLK), .D (new_AGEMA_signal_3429), .Q (new_AGEMA_signal_3430) ) ;
    buf_clk new_AGEMA_reg_buffer_1982 ( .C (CLK), .D (new_AGEMA_signal_3433), .Q (new_AGEMA_signal_3434) ) ;
    buf_clk new_AGEMA_reg_buffer_1986 ( .C (CLK), .D (new_AGEMA_signal_3437), .Q (new_AGEMA_signal_3438) ) ;
    buf_clk new_AGEMA_reg_buffer_1990 ( .C (CLK), .D (new_AGEMA_signal_3441), .Q (new_AGEMA_signal_3442) ) ;
    buf_clk new_AGEMA_reg_buffer_1994 ( .C (CLK), .D (new_AGEMA_signal_3445), .Q (new_AGEMA_signal_3446) ) ;
    buf_clk new_AGEMA_reg_buffer_1998 ( .C (CLK), .D (new_AGEMA_signal_3449), .Q (new_AGEMA_signal_3450) ) ;
    buf_clk new_AGEMA_reg_buffer_2002 ( .C (CLK), .D (new_AGEMA_signal_3453), .Q (new_AGEMA_signal_3454) ) ;
    buf_clk new_AGEMA_reg_buffer_2006 ( .C (CLK), .D (new_AGEMA_signal_3457), .Q (new_AGEMA_signal_3458) ) ;
    buf_clk new_AGEMA_reg_buffer_2010 ( .C (CLK), .D (new_AGEMA_signal_3461), .Q (new_AGEMA_signal_3462) ) ;
    buf_clk new_AGEMA_reg_buffer_2014 ( .C (CLK), .D (new_AGEMA_signal_3465), .Q (new_AGEMA_signal_3466) ) ;
    buf_clk new_AGEMA_reg_buffer_2018 ( .C (CLK), .D (new_AGEMA_signal_3469), .Q (new_AGEMA_signal_3470) ) ;
    buf_clk new_AGEMA_reg_buffer_2022 ( .C (CLK), .D (new_AGEMA_signal_3473), .Q (new_AGEMA_signal_3474) ) ;
    buf_clk new_AGEMA_reg_buffer_2026 ( .C (CLK), .D (new_AGEMA_signal_3477), .Q (new_AGEMA_signal_3478) ) ;
    buf_clk new_AGEMA_reg_buffer_2030 ( .C (CLK), .D (new_AGEMA_signal_3481), .Q (new_AGEMA_signal_3482) ) ;
    buf_clk new_AGEMA_reg_buffer_2034 ( .C (CLK), .D (new_AGEMA_signal_3485), .Q (new_AGEMA_signal_3486) ) ;
    buf_clk new_AGEMA_reg_buffer_2038 ( .C (CLK), .D (new_AGEMA_signal_3489), .Q (new_AGEMA_signal_3490) ) ;
    buf_clk new_AGEMA_reg_buffer_2042 ( .C (CLK), .D (new_AGEMA_signal_3493), .Q (new_AGEMA_signal_3494) ) ;
    buf_clk new_AGEMA_reg_buffer_2046 ( .C (CLK), .D (new_AGEMA_signal_3497), .Q (new_AGEMA_signal_3498) ) ;
    buf_clk new_AGEMA_reg_buffer_2050 ( .C (CLK), .D (new_AGEMA_signal_3501), .Q (new_AGEMA_signal_3502) ) ;
    buf_clk new_AGEMA_reg_buffer_2054 ( .C (CLK), .D (new_AGEMA_signal_3505), .Q (new_AGEMA_signal_3506) ) ;
    buf_clk new_AGEMA_reg_buffer_2058 ( .C (CLK), .D (new_AGEMA_signal_3509), .Q (new_AGEMA_signal_3510) ) ;
    buf_clk new_AGEMA_reg_buffer_2062 ( .C (CLK), .D (new_AGEMA_signal_3513), .Q (new_AGEMA_signal_3514) ) ;
    buf_clk new_AGEMA_reg_buffer_2066 ( .C (CLK), .D (new_AGEMA_signal_3517), .Q (new_AGEMA_signal_3518) ) ;
    buf_clk new_AGEMA_reg_buffer_2070 ( .C (CLK), .D (new_AGEMA_signal_3521), .Q (new_AGEMA_signal_3522) ) ;
    buf_clk new_AGEMA_reg_buffer_2074 ( .C (CLK), .D (new_AGEMA_signal_3525), .Q (new_AGEMA_signal_3526) ) ;
    buf_clk new_AGEMA_reg_buffer_2078 ( .C (CLK), .D (new_AGEMA_signal_3529), .Q (new_AGEMA_signal_3530) ) ;
    buf_clk new_AGEMA_reg_buffer_2082 ( .C (CLK), .D (new_AGEMA_signal_3533), .Q (new_AGEMA_signal_3534) ) ;
    buf_clk new_AGEMA_reg_buffer_2086 ( .C (CLK), .D (new_AGEMA_signal_3537), .Q (new_AGEMA_signal_3538) ) ;
    buf_clk new_AGEMA_reg_buffer_2090 ( .C (CLK), .D (new_AGEMA_signal_3541), .Q (new_AGEMA_signal_3542) ) ;
    buf_clk new_AGEMA_reg_buffer_2094 ( .C (CLK), .D (new_AGEMA_signal_3545), .Q (new_AGEMA_signal_3546) ) ;
    buf_clk new_AGEMA_reg_buffer_2098 ( .C (CLK), .D (new_AGEMA_signal_3549), .Q (new_AGEMA_signal_3550) ) ;
    buf_clk new_AGEMA_reg_buffer_2102 ( .C (CLK), .D (new_AGEMA_signal_3553), .Q (new_AGEMA_signal_3554) ) ;
    buf_clk new_AGEMA_reg_buffer_2106 ( .C (CLK), .D (new_AGEMA_signal_3557), .Q (new_AGEMA_signal_3558) ) ;
    buf_clk new_AGEMA_reg_buffer_2110 ( .C (CLK), .D (new_AGEMA_signal_3561), .Q (new_AGEMA_signal_3562) ) ;
    buf_clk new_AGEMA_reg_buffer_2114 ( .C (CLK), .D (new_AGEMA_signal_3565), .Q (new_AGEMA_signal_3566) ) ;
    buf_clk new_AGEMA_reg_buffer_2118 ( .C (CLK), .D (new_AGEMA_signal_3569), .Q (new_AGEMA_signal_3570) ) ;
    buf_clk new_AGEMA_reg_buffer_2122 ( .C (CLK), .D (new_AGEMA_signal_3573), .Q (new_AGEMA_signal_3574) ) ;
    buf_clk new_AGEMA_reg_buffer_2126 ( .C (CLK), .D (new_AGEMA_signal_3577), .Q (new_AGEMA_signal_3578) ) ;
    buf_clk new_AGEMA_reg_buffer_2130 ( .C (CLK), .D (new_AGEMA_signal_3581), .Q (new_AGEMA_signal_3582) ) ;
    buf_clk new_AGEMA_reg_buffer_2134 ( .C (CLK), .D (new_AGEMA_signal_3585), .Q (new_AGEMA_signal_3586) ) ;
    buf_clk new_AGEMA_reg_buffer_2138 ( .C (CLK), .D (new_AGEMA_signal_3589), .Q (new_AGEMA_signal_3590) ) ;
    buf_clk new_AGEMA_reg_buffer_2142 ( .C (CLK), .D (new_AGEMA_signal_3593), .Q (new_AGEMA_signal_3594) ) ;
    buf_clk new_AGEMA_reg_buffer_2146 ( .C (CLK), .D (new_AGEMA_signal_3597), .Q (new_AGEMA_signal_3598) ) ;
    buf_clk new_AGEMA_reg_buffer_2150 ( .C (CLK), .D (new_AGEMA_signal_3601), .Q (new_AGEMA_signal_3602) ) ;
    buf_clk new_AGEMA_reg_buffer_2154 ( .C (CLK), .D (new_AGEMA_signal_3605), .Q (new_AGEMA_signal_3606) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (CLK), .D (new_AGEMA_signal_3609), .Q (new_AGEMA_signal_3610) ) ;
    buf_clk new_AGEMA_reg_buffer_2162 ( .C (CLK), .D (new_AGEMA_signal_3613), .Q (new_AGEMA_signal_3614) ) ;
    buf_clk new_AGEMA_reg_buffer_2166 ( .C (CLK), .D (new_AGEMA_signal_3617), .Q (new_AGEMA_signal_3618) ) ;
    buf_clk new_AGEMA_reg_buffer_2170 ( .C (CLK), .D (new_AGEMA_signal_3621), .Q (new_AGEMA_signal_3622) ) ;
    buf_clk new_AGEMA_reg_buffer_2174 ( .C (CLK), .D (new_AGEMA_signal_3625), .Q (new_AGEMA_signal_3626) ) ;
    buf_clk new_AGEMA_reg_buffer_2178 ( .C (CLK), .D (new_AGEMA_signal_3629), .Q (new_AGEMA_signal_3630) ) ;
    buf_clk new_AGEMA_reg_buffer_2182 ( .C (CLK), .D (new_AGEMA_signal_3633), .Q (new_AGEMA_signal_3634) ) ;
    buf_clk new_AGEMA_reg_buffer_2186 ( .C (CLK), .D (new_AGEMA_signal_3637), .Q (new_AGEMA_signal_3638) ) ;
    buf_clk new_AGEMA_reg_buffer_2190 ( .C (CLK), .D (new_AGEMA_signal_3641), .Q (new_AGEMA_signal_3642) ) ;
    buf_clk new_AGEMA_reg_buffer_2194 ( .C (CLK), .D (new_AGEMA_signal_3645), .Q (new_AGEMA_signal_3646) ) ;
    buf_clk new_AGEMA_reg_buffer_2198 ( .C (CLK), .D (new_AGEMA_signal_3649), .Q (new_AGEMA_signal_3650) ) ;
    buf_clk new_AGEMA_reg_buffer_2202 ( .C (CLK), .D (new_AGEMA_signal_3653), .Q (new_AGEMA_signal_3654) ) ;
    buf_clk new_AGEMA_reg_buffer_2206 ( .C (CLK), .D (new_AGEMA_signal_3657), .Q (new_AGEMA_signal_3658) ) ;
    buf_clk new_AGEMA_reg_buffer_2210 ( .C (CLK), .D (new_AGEMA_signal_3661), .Q (new_AGEMA_signal_3662) ) ;
    buf_clk new_AGEMA_reg_buffer_2214 ( .C (CLK), .D (new_AGEMA_signal_3665), .Q (new_AGEMA_signal_3666) ) ;
    buf_clk new_AGEMA_reg_buffer_2218 ( .C (CLK), .D (new_AGEMA_signal_3669), .Q (new_AGEMA_signal_3670) ) ;
    buf_clk new_AGEMA_reg_buffer_2222 ( .C (CLK), .D (new_AGEMA_signal_3673), .Q (new_AGEMA_signal_3674) ) ;
    buf_clk new_AGEMA_reg_buffer_2226 ( .C (CLK), .D (new_AGEMA_signal_3677), .Q (new_AGEMA_signal_3678) ) ;
    buf_clk new_AGEMA_reg_buffer_2230 ( .C (CLK), .D (new_AGEMA_signal_3681), .Q (new_AGEMA_signal_3682) ) ;
    buf_clk new_AGEMA_reg_buffer_2234 ( .C (CLK), .D (new_AGEMA_signal_3685), .Q (new_AGEMA_signal_3686) ) ;
    buf_clk new_AGEMA_reg_buffer_2238 ( .C (CLK), .D (new_AGEMA_signal_3689), .Q (new_AGEMA_signal_3690) ) ;
    buf_clk new_AGEMA_reg_buffer_2242 ( .C (CLK), .D (new_AGEMA_signal_3693), .Q (new_AGEMA_signal_3694) ) ;
    buf_clk new_AGEMA_reg_buffer_2246 ( .C (CLK), .D (new_AGEMA_signal_3697), .Q (new_AGEMA_signal_3698) ) ;
    buf_clk new_AGEMA_reg_buffer_2250 ( .C (CLK), .D (new_AGEMA_signal_3701), .Q (new_AGEMA_signal_3702) ) ;
    buf_clk new_AGEMA_reg_buffer_2254 ( .C (CLK), .D (new_AGEMA_signal_3705), .Q (new_AGEMA_signal_3706) ) ;
    buf_clk new_AGEMA_reg_buffer_2258 ( .C (CLK), .D (new_AGEMA_signal_3709), .Q (new_AGEMA_signal_3710) ) ;
    buf_clk new_AGEMA_reg_buffer_2262 ( .C (CLK), .D (new_AGEMA_signal_3713), .Q (new_AGEMA_signal_3714) ) ;
    buf_clk new_AGEMA_reg_buffer_2266 ( .C (CLK), .D (new_AGEMA_signal_3717), .Q (new_AGEMA_signal_3718) ) ;
    buf_clk new_AGEMA_reg_buffer_2270 ( .C (CLK), .D (new_AGEMA_signal_3721), .Q (new_AGEMA_signal_3722) ) ;
    buf_clk new_AGEMA_reg_buffer_2274 ( .C (CLK), .D (new_AGEMA_signal_3725), .Q (new_AGEMA_signal_3726) ) ;
    buf_clk new_AGEMA_reg_buffer_2278 ( .C (CLK), .D (new_AGEMA_signal_3729), .Q (new_AGEMA_signal_3730) ) ;
    buf_clk new_AGEMA_reg_buffer_2282 ( .C (CLK), .D (new_AGEMA_signal_3733), .Q (new_AGEMA_signal_3734) ) ;
    buf_clk new_AGEMA_reg_buffer_2286 ( .C (CLK), .D (new_AGEMA_signal_3737), .Q (new_AGEMA_signal_3738) ) ;
    buf_clk new_AGEMA_reg_buffer_2290 ( .C (CLK), .D (new_AGEMA_signal_3741), .Q (new_AGEMA_signal_3742) ) ;
    buf_clk new_AGEMA_reg_buffer_2294 ( .C (CLK), .D (new_AGEMA_signal_3745), .Q (new_AGEMA_signal_3746) ) ;
    buf_clk new_AGEMA_reg_buffer_2298 ( .C (CLK), .D (new_AGEMA_signal_3749), .Q (new_AGEMA_signal_3750) ) ;
    buf_clk new_AGEMA_reg_buffer_2302 ( .C (CLK), .D (new_AGEMA_signal_3753), .Q (new_AGEMA_signal_3754) ) ;
    buf_clk new_AGEMA_reg_buffer_2306 ( .C (CLK), .D (new_AGEMA_signal_3757), .Q (new_AGEMA_signal_3758) ) ;
    buf_clk new_AGEMA_reg_buffer_2310 ( .C (CLK), .D (new_AGEMA_signal_3761), .Q (new_AGEMA_signal_3762) ) ;
    buf_clk new_AGEMA_reg_buffer_2314 ( .C (CLK), .D (new_AGEMA_signal_3765), .Q (new_AGEMA_signal_3766) ) ;
    buf_clk new_AGEMA_reg_buffer_2318 ( .C (CLK), .D (new_AGEMA_signal_3769), .Q (new_AGEMA_signal_3770) ) ;
    buf_clk new_AGEMA_reg_buffer_2322 ( .C (CLK), .D (new_AGEMA_signal_3773), .Q (new_AGEMA_signal_3774) ) ;
    buf_clk new_AGEMA_reg_buffer_2326 ( .C (CLK), .D (new_AGEMA_signal_3777), .Q (new_AGEMA_signal_3778) ) ;
    buf_clk new_AGEMA_reg_buffer_2330 ( .C (CLK), .D (new_AGEMA_signal_3781), .Q (new_AGEMA_signal_3782) ) ;
    buf_clk new_AGEMA_reg_buffer_2334 ( .C (CLK), .D (new_AGEMA_signal_3785), .Q (new_AGEMA_signal_3786) ) ;
    buf_clk new_AGEMA_reg_buffer_2338 ( .C (CLK), .D (new_AGEMA_signal_3789), .Q (new_AGEMA_signal_3790) ) ;
    buf_clk new_AGEMA_reg_buffer_2342 ( .C (CLK), .D (new_AGEMA_signal_3793), .Q (new_AGEMA_signal_3794) ) ;
    buf_clk new_AGEMA_reg_buffer_2346 ( .C (CLK), .D (new_AGEMA_signal_3797), .Q (new_AGEMA_signal_3798) ) ;
    buf_clk new_AGEMA_reg_buffer_2350 ( .C (CLK), .D (new_AGEMA_signal_3801), .Q (new_AGEMA_signal_3802) ) ;
    buf_clk new_AGEMA_reg_buffer_2354 ( .C (CLK), .D (new_AGEMA_signal_3805), .Q (new_AGEMA_signal_3806) ) ;
    buf_clk new_AGEMA_reg_buffer_2358 ( .C (CLK), .D (new_AGEMA_signal_3809), .Q (new_AGEMA_signal_3810) ) ;
    buf_clk new_AGEMA_reg_buffer_2362 ( .C (CLK), .D (new_AGEMA_signal_3813), .Q (new_AGEMA_signal_3814) ) ;
    buf_clk new_AGEMA_reg_buffer_2372 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_0_L5), .Q (new_AGEMA_signal_3824) ) ;
    buf_clk new_AGEMA_reg_buffer_2374 ( .C (CLK), .D (new_AGEMA_signal_1965), .Q (new_AGEMA_signal_3826) ) ;
    buf_clk new_AGEMA_reg_buffer_2378 ( .C (CLK), .D (new_AGEMA_signal_3829), .Q (new_AGEMA_signal_3830) ) ;
    buf_clk new_AGEMA_reg_buffer_2382 ( .C (CLK), .D (new_AGEMA_signal_3833), .Q (new_AGEMA_signal_3834) ) ;
    buf_clk new_AGEMA_reg_buffer_2386 ( .C (CLK), .D (new_AGEMA_signal_3837), .Q (new_AGEMA_signal_3838) ) ;
    buf_clk new_AGEMA_reg_buffer_2390 ( .C (CLK), .D (new_AGEMA_signal_3841), .Q (new_AGEMA_signal_3842) ) ;
    buf_clk new_AGEMA_reg_buffer_2392 ( .C (CLK), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_3844) ) ;
    buf_clk new_AGEMA_reg_buffer_2394 ( .C (CLK), .D (new_AGEMA_signal_2587), .Q (new_AGEMA_signal_3846) ) ;
    buf_clk new_AGEMA_reg_buffer_2404 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_1_L5), .Q (new_AGEMA_signal_3856) ) ;
    buf_clk new_AGEMA_reg_buffer_2406 ( .C (CLK), .D (new_AGEMA_signal_1967), .Q (new_AGEMA_signal_3858) ) ;
    buf_clk new_AGEMA_reg_buffer_2410 ( .C (CLK), .D (new_AGEMA_signal_3861), .Q (new_AGEMA_signal_3862) ) ;
    buf_clk new_AGEMA_reg_buffer_2414 ( .C (CLK), .D (new_AGEMA_signal_3865), .Q (new_AGEMA_signal_3866) ) ;
    buf_clk new_AGEMA_reg_buffer_2418 ( .C (CLK), .D (new_AGEMA_signal_3869), .Q (new_AGEMA_signal_3870) ) ;
    buf_clk new_AGEMA_reg_buffer_2422 ( .C (CLK), .D (new_AGEMA_signal_3873), .Q (new_AGEMA_signal_3874) ) ;
    buf_clk new_AGEMA_reg_buffer_2424 ( .C (CLK), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_3876) ) ;
    buf_clk new_AGEMA_reg_buffer_2426 ( .C (CLK), .D (new_AGEMA_signal_2599), .Q (new_AGEMA_signal_3878) ) ;
    buf_clk new_AGEMA_reg_buffer_2436 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_2_L5), .Q (new_AGEMA_signal_3888) ) ;
    buf_clk new_AGEMA_reg_buffer_2438 ( .C (CLK), .D (new_AGEMA_signal_1937), .Q (new_AGEMA_signal_3890) ) ;
    buf_clk new_AGEMA_reg_buffer_2442 ( .C (CLK), .D (new_AGEMA_signal_3893), .Q (new_AGEMA_signal_3894) ) ;
    buf_clk new_AGEMA_reg_buffer_2446 ( .C (CLK), .D (new_AGEMA_signal_3897), .Q (new_AGEMA_signal_3898) ) ;
    buf_clk new_AGEMA_reg_buffer_2448 ( .C (CLK), .D (new_AGEMA_signal_2609), .Q (new_AGEMA_signal_3900) ) ;
    buf_clk new_AGEMA_reg_buffer_2450 ( .C (CLK), .D (new_AGEMA_signal_2611), .Q (new_AGEMA_signal_3902) ) ;
    buf_clk new_AGEMA_reg_buffer_2460 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_3_L5), .Q (new_AGEMA_signal_3912) ) ;
    buf_clk new_AGEMA_reg_buffer_2462 ( .C (CLK), .D (new_AGEMA_signal_1939), .Q (new_AGEMA_signal_3914) ) ;
    buf_clk new_AGEMA_reg_buffer_2466 ( .C (CLK), .D (new_AGEMA_signal_3917), .Q (new_AGEMA_signal_3918) ) ;
    buf_clk new_AGEMA_reg_buffer_2470 ( .C (CLK), .D (new_AGEMA_signal_3921), .Q (new_AGEMA_signal_3922) ) ;
    buf_clk new_AGEMA_reg_buffer_2472 ( .C (CLK), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_3924) ) ;
    buf_clk new_AGEMA_reg_buffer_2474 ( .C (CLK), .D (new_AGEMA_signal_2623), .Q (new_AGEMA_signal_3926) ) ;
    buf_clk new_AGEMA_reg_buffer_2484 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_4_L5), .Q (new_AGEMA_signal_3936) ) ;
    buf_clk new_AGEMA_reg_buffer_2486 ( .C (CLK), .D (new_AGEMA_signal_1973), .Q (new_AGEMA_signal_3938) ) ;
    buf_clk new_AGEMA_reg_buffer_2490 ( .C (CLK), .D (new_AGEMA_signal_3941), .Q (new_AGEMA_signal_3942) ) ;
    buf_clk new_AGEMA_reg_buffer_2494 ( .C (CLK), .D (new_AGEMA_signal_3945), .Q (new_AGEMA_signal_3946) ) ;
    buf_clk new_AGEMA_reg_buffer_2498 ( .C (CLK), .D (new_AGEMA_signal_3949), .Q (new_AGEMA_signal_3950) ) ;
    buf_clk new_AGEMA_reg_buffer_2502 ( .C (CLK), .D (new_AGEMA_signal_3953), .Q (new_AGEMA_signal_3954) ) ;
    buf_clk new_AGEMA_reg_buffer_2504 ( .C (CLK), .D (new_AGEMA_signal_2633), .Q (new_AGEMA_signal_3956) ) ;
    buf_clk new_AGEMA_reg_buffer_2506 ( .C (CLK), .D (new_AGEMA_signal_2635), .Q (new_AGEMA_signal_3958) ) ;
    buf_clk new_AGEMA_reg_buffer_2516 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_5_L5), .Q (new_AGEMA_signal_3968) ) ;
    buf_clk new_AGEMA_reg_buffer_2518 ( .C (CLK), .D (new_AGEMA_signal_1975), .Q (new_AGEMA_signal_3970) ) ;
    buf_clk new_AGEMA_reg_buffer_2522 ( .C (CLK), .D (new_AGEMA_signal_3973), .Q (new_AGEMA_signal_3974) ) ;
    buf_clk new_AGEMA_reg_buffer_2526 ( .C (CLK), .D (new_AGEMA_signal_3977), .Q (new_AGEMA_signal_3978) ) ;
    buf_clk new_AGEMA_reg_buffer_2530 ( .C (CLK), .D (new_AGEMA_signal_3981), .Q (new_AGEMA_signal_3982) ) ;
    buf_clk new_AGEMA_reg_buffer_2534 ( .C (CLK), .D (new_AGEMA_signal_3985), .Q (new_AGEMA_signal_3986) ) ;
    buf_clk new_AGEMA_reg_buffer_2536 ( .C (CLK), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_3988) ) ;
    buf_clk new_AGEMA_reg_buffer_2538 ( .C (CLK), .D (new_AGEMA_signal_2647), .Q (new_AGEMA_signal_3990) ) ;
    buf_clk new_AGEMA_reg_buffer_2548 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_6_L5), .Q (new_AGEMA_signal_4000) ) ;
    buf_clk new_AGEMA_reg_buffer_2550 ( .C (CLK), .D (new_AGEMA_signal_1945), .Q (new_AGEMA_signal_4002) ) ;
    buf_clk new_AGEMA_reg_buffer_2554 ( .C (CLK), .D (new_AGEMA_signal_4005), .Q (new_AGEMA_signal_4006) ) ;
    buf_clk new_AGEMA_reg_buffer_2558 ( .C (CLK), .D (new_AGEMA_signal_4009), .Q (new_AGEMA_signal_4010) ) ;
    buf_clk new_AGEMA_reg_buffer_2560 ( .C (CLK), .D (new_AGEMA_signal_2657), .Q (new_AGEMA_signal_4012) ) ;
    buf_clk new_AGEMA_reg_buffer_2562 ( .C (CLK), .D (new_AGEMA_signal_2659), .Q (new_AGEMA_signal_4014) ) ;
    buf_clk new_AGEMA_reg_buffer_2572 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_7_L5), .Q (new_AGEMA_signal_4024) ) ;
    buf_clk new_AGEMA_reg_buffer_2574 ( .C (CLK), .D (new_AGEMA_signal_1947), .Q (new_AGEMA_signal_4026) ) ;
    buf_clk new_AGEMA_reg_buffer_2578 ( .C (CLK), .D (new_AGEMA_signal_4029), .Q (new_AGEMA_signal_4030) ) ;
    buf_clk new_AGEMA_reg_buffer_2582 ( .C (CLK), .D (new_AGEMA_signal_4033), .Q (new_AGEMA_signal_4034) ) ;
    buf_clk new_AGEMA_reg_buffer_2584 ( .C (CLK), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_4036) ) ;
    buf_clk new_AGEMA_reg_buffer_2586 ( .C (CLK), .D (new_AGEMA_signal_2671), .Q (new_AGEMA_signal_4038) ) ;
    buf_clk new_AGEMA_reg_buffer_2596 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_8_L5), .Q (new_AGEMA_signal_4048) ) ;
    buf_clk new_AGEMA_reg_buffer_2598 ( .C (CLK), .D (new_AGEMA_signal_1981), .Q (new_AGEMA_signal_4050) ) ;
    buf_clk new_AGEMA_reg_buffer_2602 ( .C (CLK), .D (new_AGEMA_signal_4053), .Q (new_AGEMA_signal_4054) ) ;
    buf_clk new_AGEMA_reg_buffer_2606 ( .C (CLK), .D (new_AGEMA_signal_4057), .Q (new_AGEMA_signal_4058) ) ;
    buf_clk new_AGEMA_reg_buffer_2610 ( .C (CLK), .D (new_AGEMA_signal_4061), .Q (new_AGEMA_signal_4062) ) ;
    buf_clk new_AGEMA_reg_buffer_2614 ( .C (CLK), .D (new_AGEMA_signal_4065), .Q (new_AGEMA_signal_4066) ) ;
    buf_clk new_AGEMA_reg_buffer_2616 ( .C (CLK), .D (new_AGEMA_signal_2681), .Q (new_AGEMA_signal_4068) ) ;
    buf_clk new_AGEMA_reg_buffer_2618 ( .C (CLK), .D (new_AGEMA_signal_2683), .Q (new_AGEMA_signal_4070) ) ;
    buf_clk new_AGEMA_reg_buffer_2628 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_9_L5), .Q (new_AGEMA_signal_4080) ) ;
    buf_clk new_AGEMA_reg_buffer_2630 ( .C (CLK), .D (new_AGEMA_signal_1983), .Q (new_AGEMA_signal_4082) ) ;
    buf_clk new_AGEMA_reg_buffer_2634 ( .C (CLK), .D (new_AGEMA_signal_4085), .Q (new_AGEMA_signal_4086) ) ;
    buf_clk new_AGEMA_reg_buffer_2638 ( .C (CLK), .D (new_AGEMA_signal_4089), .Q (new_AGEMA_signal_4090) ) ;
    buf_clk new_AGEMA_reg_buffer_2642 ( .C (CLK), .D (new_AGEMA_signal_4093), .Q (new_AGEMA_signal_4094) ) ;
    buf_clk new_AGEMA_reg_buffer_2646 ( .C (CLK), .D (new_AGEMA_signal_4097), .Q (new_AGEMA_signal_4098) ) ;
    buf_clk new_AGEMA_reg_buffer_2648 ( .C (CLK), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_4100) ) ;
    buf_clk new_AGEMA_reg_buffer_2650 ( .C (CLK), .D (new_AGEMA_signal_2695), .Q (new_AGEMA_signal_4102) ) ;
    buf_clk new_AGEMA_reg_buffer_2660 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_10_L5), .Q (new_AGEMA_signal_4112) ) ;
    buf_clk new_AGEMA_reg_buffer_2662 ( .C (CLK), .D (new_AGEMA_signal_1953), .Q (new_AGEMA_signal_4114) ) ;
    buf_clk new_AGEMA_reg_buffer_2666 ( .C (CLK), .D (new_AGEMA_signal_4117), .Q (new_AGEMA_signal_4118) ) ;
    buf_clk new_AGEMA_reg_buffer_2670 ( .C (CLK), .D (new_AGEMA_signal_4121), .Q (new_AGEMA_signal_4122) ) ;
    buf_clk new_AGEMA_reg_buffer_2672 ( .C (CLK), .D (new_AGEMA_signal_2705), .Q (new_AGEMA_signal_4124) ) ;
    buf_clk new_AGEMA_reg_buffer_2674 ( .C (CLK), .D (new_AGEMA_signal_2707), .Q (new_AGEMA_signal_4126) ) ;
    buf_clk new_AGEMA_reg_buffer_2684 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_11_L5), .Q (new_AGEMA_signal_4136) ) ;
    buf_clk new_AGEMA_reg_buffer_2686 ( .C (CLK), .D (new_AGEMA_signal_1955), .Q (new_AGEMA_signal_4138) ) ;
    buf_clk new_AGEMA_reg_buffer_2690 ( .C (CLK), .D (new_AGEMA_signal_4141), .Q (new_AGEMA_signal_4142) ) ;
    buf_clk new_AGEMA_reg_buffer_2694 ( .C (CLK), .D (new_AGEMA_signal_4145), .Q (new_AGEMA_signal_4146) ) ;
    buf_clk new_AGEMA_reg_buffer_2696 ( .C (CLK), .D (new_AGEMA_signal_2717), .Q (new_AGEMA_signal_4148) ) ;
    buf_clk new_AGEMA_reg_buffer_2698 ( .C (CLK), .D (new_AGEMA_signal_2719), .Q (new_AGEMA_signal_4150) ) ;
    buf_clk new_AGEMA_reg_buffer_2708 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_12_L5), .Q (new_AGEMA_signal_4160) ) ;
    buf_clk new_AGEMA_reg_buffer_2710 ( .C (CLK), .D (new_AGEMA_signal_1989), .Q (new_AGEMA_signal_4162) ) ;
    buf_clk new_AGEMA_reg_buffer_2714 ( .C (CLK), .D (new_AGEMA_signal_4165), .Q (new_AGEMA_signal_4166) ) ;
    buf_clk new_AGEMA_reg_buffer_2718 ( .C (CLK), .D (new_AGEMA_signal_4169), .Q (new_AGEMA_signal_4170) ) ;
    buf_clk new_AGEMA_reg_buffer_2722 ( .C (CLK), .D (new_AGEMA_signal_4173), .Q (new_AGEMA_signal_4174) ) ;
    buf_clk new_AGEMA_reg_buffer_2726 ( .C (CLK), .D (new_AGEMA_signal_4177), .Q (new_AGEMA_signal_4178) ) ;
    buf_clk new_AGEMA_reg_buffer_2728 ( .C (CLK), .D (new_AGEMA_signal_2729), .Q (new_AGEMA_signal_4180) ) ;
    buf_clk new_AGEMA_reg_buffer_2730 ( .C (CLK), .D (new_AGEMA_signal_2731), .Q (new_AGEMA_signal_4182) ) ;
    buf_clk new_AGEMA_reg_buffer_2740 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_13_L5), .Q (new_AGEMA_signal_4192) ) ;
    buf_clk new_AGEMA_reg_buffer_2742 ( .C (CLK), .D (new_AGEMA_signal_1991), .Q (new_AGEMA_signal_4194) ) ;
    buf_clk new_AGEMA_reg_buffer_2746 ( .C (CLK), .D (new_AGEMA_signal_4197), .Q (new_AGEMA_signal_4198) ) ;
    buf_clk new_AGEMA_reg_buffer_2750 ( .C (CLK), .D (new_AGEMA_signal_4201), .Q (new_AGEMA_signal_4202) ) ;
    buf_clk new_AGEMA_reg_buffer_2754 ( .C (CLK), .D (new_AGEMA_signal_4205), .Q (new_AGEMA_signal_4206) ) ;
    buf_clk new_AGEMA_reg_buffer_2758 ( .C (CLK), .D (new_AGEMA_signal_4209), .Q (new_AGEMA_signal_4210) ) ;
    buf_clk new_AGEMA_reg_buffer_2760 ( .C (CLK), .D (new_AGEMA_signal_2741), .Q (new_AGEMA_signal_4212) ) ;
    buf_clk new_AGEMA_reg_buffer_2762 ( .C (CLK), .D (new_AGEMA_signal_2743), .Q (new_AGEMA_signal_4214) ) ;
    buf_clk new_AGEMA_reg_buffer_2772 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_14_L5), .Q (new_AGEMA_signal_4224) ) ;
    buf_clk new_AGEMA_reg_buffer_2774 ( .C (CLK), .D (new_AGEMA_signal_1961), .Q (new_AGEMA_signal_4226) ) ;
    buf_clk new_AGEMA_reg_buffer_2778 ( .C (CLK), .D (new_AGEMA_signal_4229), .Q (new_AGEMA_signal_4230) ) ;
    buf_clk new_AGEMA_reg_buffer_2782 ( .C (CLK), .D (new_AGEMA_signal_4233), .Q (new_AGEMA_signal_4234) ) ;
    buf_clk new_AGEMA_reg_buffer_2784 ( .C (CLK), .D (new_AGEMA_signal_2753), .Q (new_AGEMA_signal_4236) ) ;
    buf_clk new_AGEMA_reg_buffer_2786 ( .C (CLK), .D (new_AGEMA_signal_2755), .Q (new_AGEMA_signal_4238) ) ;
    buf_clk new_AGEMA_reg_buffer_2796 ( .C (CLK), .D (LED_128_Instance_SBox_Instance_15_L5), .Q (new_AGEMA_signal_4248) ) ;
    buf_clk new_AGEMA_reg_buffer_2798 ( .C (CLK), .D (new_AGEMA_signal_1963), .Q (new_AGEMA_signal_4250) ) ;
    buf_clk new_AGEMA_reg_buffer_2802 ( .C (CLK), .D (new_AGEMA_signal_4253), .Q (new_AGEMA_signal_4254) ) ;
    buf_clk new_AGEMA_reg_buffer_2806 ( .C (CLK), .D (new_AGEMA_signal_4257), .Q (new_AGEMA_signal_4258) ) ;
    buf_clk new_AGEMA_reg_buffer_2808 ( .C (CLK), .D (new_AGEMA_signal_2765), .Q (new_AGEMA_signal_4260) ) ;
    buf_clk new_AGEMA_reg_buffer_2810 ( .C (CLK), .D (new_AGEMA_signal_2767), .Q (new_AGEMA_signal_4262) ) ;
    buf_clk new_AGEMA_reg_buffer_2812 ( .C (CLK), .D (LED_128_Instance_subcells_out[60]), .Q (new_AGEMA_signal_4264) ) ;
    buf_clk new_AGEMA_reg_buffer_2814 ( .C (CLK), .D (new_AGEMA_signal_1931), .Q (new_AGEMA_signal_4266) ) ;
    buf_clk new_AGEMA_reg_buffer_2816 ( .C (CLK), .D (LED_128_Instance_subcells_out[20]), .Q (new_AGEMA_signal_4268) ) ;
    buf_clk new_AGEMA_reg_buffer_2818 ( .C (CLK), .D (new_AGEMA_signal_1943), .Q (new_AGEMA_signal_4270) ) ;
    buf_clk new_AGEMA_reg_buffer_2820 ( .C (CLK), .D (LED_128_Instance_subcells_out[40]), .Q (new_AGEMA_signal_4272) ) ;
    buf_clk new_AGEMA_reg_buffer_2822 ( .C (CLK), .D (new_AGEMA_signal_1915), .Q (new_AGEMA_signal_4274) ) ;
    buf_clk new_AGEMA_reg_buffer_2824 ( .C (CLK), .D (LED_128_Instance_subcells_out[0]), .Q (new_AGEMA_signal_4276) ) ;
    buf_clk new_AGEMA_reg_buffer_2826 ( .C (CLK), .D (new_AGEMA_signal_1933), .Q (new_AGEMA_signal_4278) ) ;
    buf_clk new_AGEMA_reg_buffer_2828 ( .C (CLK), .D (LED_128_Instance_subcells_out[48]), .Q (new_AGEMA_signal_4280) ) ;
    buf_clk new_AGEMA_reg_buffer_2830 ( .C (CLK), .D (new_AGEMA_signal_1957), .Q (new_AGEMA_signal_4282) ) ;
    buf_clk new_AGEMA_reg_buffer_2832 ( .C (CLK), .D (LED_128_Instance_subcells_out[24]), .Q (new_AGEMA_signal_4284) ) ;
    buf_clk new_AGEMA_reg_buffer_2834 ( .C (CLK), .D (new_AGEMA_signal_1901), .Q (new_AGEMA_signal_4286) ) ;
    buf_clk new_AGEMA_reg_buffer_2836 ( .C (CLK), .D (LED_128_Instance_subcells_out[44]), .Q (new_AGEMA_signal_4288) ) ;
    buf_clk new_AGEMA_reg_buffer_2838 ( .C (CLK), .D (new_AGEMA_signal_1917), .Q (new_AGEMA_signal_4290) ) ;
    buf_clk new_AGEMA_reg_buffer_2840 ( .C (CLK), .D (LED_128_Instance_subcells_out[4]), .Q (new_AGEMA_signal_4292) ) ;
    buf_clk new_AGEMA_reg_buffer_2842 ( .C (CLK), .D (new_AGEMA_signal_1935), .Q (new_AGEMA_signal_4294) ) ;
    buf_clk new_AGEMA_reg_buffer_2844 ( .C (CLK), .D (LED_128_Instance_subcells_out[52]), .Q (new_AGEMA_signal_4296) ) ;
    buf_clk new_AGEMA_reg_buffer_2846 ( .C (CLK), .D (new_AGEMA_signal_1959), .Q (new_AGEMA_signal_4298) ) ;
    buf_clk new_AGEMA_reg_buffer_2848 ( .C (CLK), .D (LED_128_Instance_subcells_out[28]), .Q (new_AGEMA_signal_4300) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (CLK), .D (new_AGEMA_signal_1903), .Q (new_AGEMA_signal_4302) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (CLK), .D (LED_128_Instance_subcells_out[32]), .Q (new_AGEMA_signal_4304) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (CLK), .D (new_AGEMA_signal_1949), .Q (new_AGEMA_signal_4306) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (CLK), .D (LED_128_Instance_subcells_out[8]), .Q (new_AGEMA_signal_4308) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (CLK), .D (new_AGEMA_signal_1887), .Q (new_AGEMA_signal_4310) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (CLK), .D (LED_128_Instance_subcells_out[56]), .Q (new_AGEMA_signal_4312) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (CLK), .D (new_AGEMA_signal_1929), .Q (new_AGEMA_signal_4314) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (CLK), .D (LED_128_Instance_subcells_out[16]), .Q (new_AGEMA_signal_4316) ) ;
    buf_clk new_AGEMA_reg_buffer_2866 ( .C (CLK), .D (new_AGEMA_signal_1941), .Q (new_AGEMA_signal_4318) ) ;
    buf_clk new_AGEMA_reg_buffer_2868 ( .C (CLK), .D (LED_128_Instance_subcells_out[36]), .Q (new_AGEMA_signal_4320) ) ;
    buf_clk new_AGEMA_reg_buffer_2870 ( .C (CLK), .D (new_AGEMA_signal_1951), .Q (new_AGEMA_signal_4322) ) ;
    buf_clk new_AGEMA_reg_buffer_2872 ( .C (CLK), .D (LED_128_Instance_subcells_out[12]), .Q (new_AGEMA_signal_4324) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (CLK), .D (new_AGEMA_signal_1889), .Q (new_AGEMA_signal_4326) ) ;
    buf_clk new_AGEMA_reg_buffer_2878 ( .C (CLK), .D (new_AGEMA_signal_4329), .Q (new_AGEMA_signal_4330) ) ;
    buf_clk new_AGEMA_reg_buffer_2882 ( .C (CLK), .D (new_AGEMA_signal_4333), .Q (new_AGEMA_signal_4334) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (CLK), .D (new_AGEMA_signal_4337), .Q (new_AGEMA_signal_4338) ) ;
    buf_clk new_AGEMA_reg_buffer_2890 ( .C (CLK), .D (new_AGEMA_signal_4341), .Q (new_AGEMA_signal_4342) ) ;
    buf_clk new_AGEMA_reg_buffer_2894 ( .C (CLK), .D (new_AGEMA_signal_4345), .Q (new_AGEMA_signal_4346) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (CLK), .D (new_AGEMA_signal_4349), .Q (new_AGEMA_signal_4350) ) ;
    buf_clk new_AGEMA_reg_buffer_2902 ( .C (CLK), .D (new_AGEMA_signal_4353), .Q (new_AGEMA_signal_4354) ) ;
    buf_clk new_AGEMA_reg_buffer_2906 ( .C (CLK), .D (new_AGEMA_signal_4357), .Q (new_AGEMA_signal_4358) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (CLK), .D (new_AGEMA_signal_4361), .Q (new_AGEMA_signal_4362) ) ;
    buf_clk new_AGEMA_reg_buffer_2914 ( .C (CLK), .D (new_AGEMA_signal_4365), .Q (new_AGEMA_signal_4366) ) ;
    buf_clk new_AGEMA_reg_buffer_2918 ( .C (CLK), .D (new_AGEMA_signal_4369), .Q (new_AGEMA_signal_4370) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_0_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}), .a ({new_AGEMA_signal_2783, new_AGEMA_signal_2779}), .c ({new_AGEMA_signal_2171, LED_128_Instance_state0[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_1_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}), .a ({new_AGEMA_signal_2791, new_AGEMA_signal_2787}), .c ({new_AGEMA_signal_2268, LED_128_Instance_state0[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_2_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .a ({new_AGEMA_signal_2803, new_AGEMA_signal_2799}), .c ({new_AGEMA_signal_2191, LED_128_Instance_state0[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_3_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .a ({new_AGEMA_signal_2815, new_AGEMA_signal_2811}), .c ({new_AGEMA_signal_2222, LED_128_Instance_state0[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_4_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}), .a ({new_AGEMA_signal_2823, new_AGEMA_signal_2819}), .c ({new_AGEMA_signal_2192, LED_128_Instance_state0[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_5_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}), .a ({new_AGEMA_signal_2831, new_AGEMA_signal_2827}), .c ({new_AGEMA_signal_2269, LED_128_Instance_state0[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_6_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .a ({new_AGEMA_signal_2839, new_AGEMA_signal_2835}), .c ({new_AGEMA_signal_2193, LED_128_Instance_state0[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_7_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .a ({new_AGEMA_signal_2847, new_AGEMA_signal_2843}), .c ({new_AGEMA_signal_2194, LED_128_Instance_state0[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_8_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}), .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2851}), .c ({new_AGEMA_signal_2195, LED_128_Instance_state0[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_9_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}), .a ({new_AGEMA_signal_2863, new_AGEMA_signal_2859}), .c ({new_AGEMA_signal_2223, LED_128_Instance_state0[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_10_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .a ({new_AGEMA_signal_2871, new_AGEMA_signal_2867}), .c ({new_AGEMA_signal_2196, LED_128_Instance_state0[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_11_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2875}), .c ({new_AGEMA_signal_2197, LED_128_Instance_state0[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_12_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}), .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2883}), .c ({new_AGEMA_signal_2198, LED_128_Instance_state0[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_13_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}), .a ({new_AGEMA_signal_2895, new_AGEMA_signal_2891}), .c ({new_AGEMA_signal_2224, LED_128_Instance_state0[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_14_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2899}), .c ({new_AGEMA_signal_2199, LED_128_Instance_state0[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_15_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .a ({new_AGEMA_signal_2911, new_AGEMA_signal_2907}), .c ({new_AGEMA_signal_2225, LED_128_Instance_state0[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_16_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2288, LED_128_Instance_mixcolumns_out[16]}), .a ({new_AGEMA_signal_2919, new_AGEMA_signal_2915}), .c ({new_AGEMA_signal_2310, LED_128_Instance_state0[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_17_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2340, LED_128_Instance_mixcolumns_out[17]}), .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2923}), .c ({new_AGEMA_signal_2355, LED_128_Instance_state0[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_18_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}), .a ({new_AGEMA_signal_2935, new_AGEMA_signal_2931}), .c ({new_AGEMA_signal_2356, LED_128_Instance_state0[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_19_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .a ({new_AGEMA_signal_2943, new_AGEMA_signal_2939}), .c ({new_AGEMA_signal_2270, LED_128_Instance_state0[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_20_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2252, LED_128_Instance_mixcolumns_out[20]}), .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2947}), .c ({new_AGEMA_signal_2271, LED_128_Instance_state0[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_21_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2297, LED_128_Instance_mixcolumns_out[21]}), .a ({new_AGEMA_signal_2959, new_AGEMA_signal_2955}), .c ({new_AGEMA_signal_2311, LED_128_Instance_state0[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_22_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}), .a ({new_AGEMA_signal_2967, new_AGEMA_signal_2963}), .c ({new_AGEMA_signal_2357, LED_128_Instance_state0[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_23_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .a ({new_AGEMA_signal_2975, new_AGEMA_signal_2971}), .c ({new_AGEMA_signal_2272, LED_128_Instance_state0[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_24_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2258, LED_128_Instance_mixcolumns_out[24]}), .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2979}), .c ({new_AGEMA_signal_2273, LED_128_Instance_state0[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_25_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2304, LED_128_Instance_mixcolumns_out[25]}), .a ({new_AGEMA_signal_2991, new_AGEMA_signal_2987}), .c ({new_AGEMA_signal_2312, LED_128_Instance_state0[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_26_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}), .a ({new_AGEMA_signal_2999, new_AGEMA_signal_2995}), .c ({new_AGEMA_signal_2313, LED_128_Instance_state0[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_27_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .a ({new_AGEMA_signal_3007, new_AGEMA_signal_3003}), .c ({new_AGEMA_signal_2274, LED_128_Instance_state0[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_28_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2308, LED_128_Instance_mixcolumns_out[28]}), .a ({new_AGEMA_signal_3015, new_AGEMA_signal_3011}), .c ({new_AGEMA_signal_2314, LED_128_Instance_state0[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_29_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2354, LED_128_Instance_mixcolumns_out[29]}), .a ({new_AGEMA_signal_3023, new_AGEMA_signal_3019}), .c ({new_AGEMA_signal_2358, LED_128_Instance_state0[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_30_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}), .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3027}), .c ({new_AGEMA_signal_2315, LED_128_Instance_state0[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_31_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .a ({new_AGEMA_signal_3039, new_AGEMA_signal_3035}), .c ({new_AGEMA_signal_2275, LED_128_Instance_state0[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_32_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2336, LED_128_Instance_mixcolumns_out[32]}), .a ({new_AGEMA_signal_3047, new_AGEMA_signal_3043}), .c ({new_AGEMA_signal_2359, LED_128_Instance_state0[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_33_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2385, LED_128_Instance_mixcolumns_out[33]}), .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3051}), .c ({new_AGEMA_signal_2395, LED_128_Instance_state0[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_34_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2334, LED_128_Instance_mixcolumns_out[34]}), .a ({new_AGEMA_signal_3063, new_AGEMA_signal_3059}), .c ({new_AGEMA_signal_2360, LED_128_Instance_state0[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_35_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2428, LED_128_Instance_mixcolumns_out[35]}), .a ({new_AGEMA_signal_3071, new_AGEMA_signal_3067}), .c ({new_AGEMA_signal_2435, LED_128_Instance_state0[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_36_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2341, LED_128_Instance_mixcolumns_out[36]}), .a ({new_AGEMA_signal_3079, new_AGEMA_signal_3075}), .c ({new_AGEMA_signal_2361, LED_128_Instance_state0[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_37_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2343, LED_128_Instance_mixcolumns_out[37]}), .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3083}), .c ({new_AGEMA_signal_2362, LED_128_Instance_state0[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_38_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2290, LED_128_Instance_mixcolumns_out[38]}), .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3091}), .c ({new_AGEMA_signal_2316, LED_128_Instance_state0[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_39_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2430, LED_128_Instance_mixcolumns_out[39]}), .a ({new_AGEMA_signal_3103, new_AGEMA_signal_3099}), .c ({new_AGEMA_signal_2436, LED_128_Instance_state0[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_40_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2345, LED_128_Instance_mixcolumns_out[40]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3107}), .c ({new_AGEMA_signal_2363, LED_128_Instance_state0[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_41_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2347, LED_128_Instance_mixcolumns_out[41]}), .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3115}), .c ({new_AGEMA_signal_2364, LED_128_Instance_state0[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_42_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2298, LED_128_Instance_mixcolumns_out[42]}), .a ({new_AGEMA_signal_3127, new_AGEMA_signal_3123}), .c ({new_AGEMA_signal_2317, LED_128_Instance_state0[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_43_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2391, LED_128_Instance_mixcolumns_out[43]}), .a ({new_AGEMA_signal_3139, new_AGEMA_signal_3135}), .c ({new_AGEMA_signal_2396, LED_128_Instance_state0[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_44_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2350, LED_128_Instance_mixcolumns_out[44]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3143}), .c ({new_AGEMA_signal_2365, LED_128_Instance_state0[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_45_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2394, LED_128_Instance_mixcolumns_out[45]}), .a ({new_AGEMA_signal_3155, new_AGEMA_signal_3151}), .c ({new_AGEMA_signal_2397, LED_128_Instance_state0[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_46_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2348, LED_128_Instance_mixcolumns_out[46]}), .a ({new_AGEMA_signal_3163, new_AGEMA_signal_3159}), .c ({new_AGEMA_signal_2366, LED_128_Instance_state0[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_47_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2393, LED_128_Instance_mixcolumns_out[47]}), .a ({new_AGEMA_signal_3171, new_AGEMA_signal_3167}), .c ({new_AGEMA_signal_2398, LED_128_Instance_state0[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_48_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2487, LED_128_Instance_mixcolumns_out[48]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3175}), .c ({new_AGEMA_signal_2492, LED_128_Instance_state0[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_49_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2500, LED_128_Instance_mixcolumns_out[49]}), .a ({new_AGEMA_signal_3187, new_AGEMA_signal_3183}), .c ({new_AGEMA_signal_2502, LED_128_Instance_state0[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_50_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2427, LED_128_Instance_mixcolumns_out[50]}), .a ({new_AGEMA_signal_3195, new_AGEMA_signal_3191}), .c ({new_AGEMA_signal_2437, LED_128_Instance_state0[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_51_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2426, LED_128_Instance_mixcolumns_out[51]}), .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3199}), .c ({new_AGEMA_signal_2438, LED_128_Instance_state0[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_52_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2489, LED_128_Instance_mixcolumns_out[52]}), .a ({new_AGEMA_signal_3211, new_AGEMA_signal_3207}), .c ({new_AGEMA_signal_2493, LED_128_Instance_state0[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_53_U1 ( .s (new_AGEMA_signal_3131), .b ({new_AGEMA_signal_2501, LED_128_Instance_mixcolumns_out[53]}), .a ({new_AGEMA_signal_3219, new_AGEMA_signal_3215}), .c ({new_AGEMA_signal_2503, LED_128_Instance_state0[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_54_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2387, LED_128_Instance_mixcolumns_out[54]}), .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3223}), .c ({new_AGEMA_signal_2399, LED_128_Instance_state0[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_55_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2429, LED_128_Instance_mixcolumns_out[55]}), .a ({new_AGEMA_signal_3235, new_AGEMA_signal_3231}), .c ({new_AGEMA_signal_2439, LED_128_Instance_state0[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_56_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2481, LED_128_Instance_mixcolumns_out[56]}), .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3239}), .c ({new_AGEMA_signal_2484, LED_128_Instance_state0[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_57_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2490, LED_128_Instance_mixcolumns_out[57]}), .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3247}), .c ({new_AGEMA_signal_2494, LED_128_Instance_state0[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_58_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2390, LED_128_Instance_mixcolumns_out[58]}), .a ({new_AGEMA_signal_3259, new_AGEMA_signal_3255}), .c ({new_AGEMA_signal_2400, LED_128_Instance_state0[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_59_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2389, LED_128_Instance_mixcolumns_out[59]}), .a ({new_AGEMA_signal_3267, new_AGEMA_signal_3263}), .c ({new_AGEMA_signal_2401, LED_128_Instance_state0[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_60_U1 ( .s (new_AGEMA_signal_2775), .b ({new_AGEMA_signal_2483, LED_128_Instance_mixcolumns_out[60]}), .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3271}), .c ({new_AGEMA_signal_2485, LED_128_Instance_state0[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_61_U1 ( .s (new_AGEMA_signal_2807), .b ({new_AGEMA_signal_2491, LED_128_Instance_mixcolumns_out[61]}), .a ({new_AGEMA_signal_3283, new_AGEMA_signal_3279}), .c ({new_AGEMA_signal_2495, LED_128_Instance_state0[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_62_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2433, LED_128_Instance_mixcolumns_out[62]}), .a ({new_AGEMA_signal_3291, new_AGEMA_signal_3287}), .c ({new_AGEMA_signal_2440, LED_128_Instance_state0[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state0_mux_inst_63_U1 ( .s (new_AGEMA_signal_2795), .b ({new_AGEMA_signal_2432, LED_128_Instance_mixcolumns_out[63]}), .a ({new_AGEMA_signal_3299, new_AGEMA_signal_3295}), .c ({new_AGEMA_signal_2441, LED_128_Instance_state0[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_0_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2171, LED_128_Instance_state0[0]}), .a ({new_AGEMA_signal_3311, new_AGEMA_signal_3307}), .c ({new_AGEMA_signal_2201, LED_128_Instance_state1[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_1_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2268, LED_128_Instance_state0[1]}), .a ({new_AGEMA_signal_3319, new_AGEMA_signal_3315}), .c ({new_AGEMA_signal_2319, LED_128_Instance_state1[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_2_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2191, LED_128_Instance_state0[2]}), .a ({new_AGEMA_signal_3327, new_AGEMA_signal_3323}), .c ({new_AGEMA_signal_2227, LED_128_Instance_state1[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_3_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2222, LED_128_Instance_state0[3]}), .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3331}), .c ({new_AGEMA_signal_2277, LED_128_Instance_state1[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_4_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2192, LED_128_Instance_state0[4]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3339}), .c ({new_AGEMA_signal_2229, LED_128_Instance_state1[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_5_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2269, LED_128_Instance_state0[5]}), .a ({new_AGEMA_signal_3351, new_AGEMA_signal_3347}), .c ({new_AGEMA_signal_2321, LED_128_Instance_state1[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_6_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2193, LED_128_Instance_state0[6]}), .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3355}), .c ({new_AGEMA_signal_2231, LED_128_Instance_state1[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_7_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2194, LED_128_Instance_state0[7]}), .a ({new_AGEMA_signal_3367, new_AGEMA_signal_3363}), .c ({new_AGEMA_signal_2233, LED_128_Instance_state1[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_8_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2195, LED_128_Instance_state0[8]}), .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3371}), .c ({new_AGEMA_signal_2235, LED_128_Instance_state1[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_9_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2223, LED_128_Instance_state0[9]}), .a ({new_AGEMA_signal_3383, new_AGEMA_signal_3379}), .c ({new_AGEMA_signal_2279, LED_128_Instance_state1[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_10_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2196, LED_128_Instance_state0[10]}), .a ({new_AGEMA_signal_3391, new_AGEMA_signal_3387}), .c ({new_AGEMA_signal_2237, LED_128_Instance_state1[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_11_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2197, LED_128_Instance_state0[11]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3395}), .c ({new_AGEMA_signal_2239, LED_128_Instance_state1[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_12_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2198, LED_128_Instance_state0[12]}), .a ({new_AGEMA_signal_3407, new_AGEMA_signal_3403}), .c ({new_AGEMA_signal_2241, LED_128_Instance_state1[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_13_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2224, LED_128_Instance_state0[13]}), .a ({new_AGEMA_signal_3415, new_AGEMA_signal_3411}), .c ({new_AGEMA_signal_2281, LED_128_Instance_state1[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_14_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2199, LED_128_Instance_state0[14]}), .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3419}), .c ({new_AGEMA_signal_2243, LED_128_Instance_state1[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_15_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2225, LED_128_Instance_state0[15]}), .a ({new_AGEMA_signal_3431, new_AGEMA_signal_3427}), .c ({new_AGEMA_signal_2283, LED_128_Instance_state1[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_16_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2310, LED_128_Instance_state0[16]}), .a ({new_AGEMA_signal_3439, new_AGEMA_signal_3435}), .c ({new_AGEMA_signal_2368, LED_128_Instance_state1[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_17_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2355, LED_128_Instance_state0[17]}), .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3443}), .c ({new_AGEMA_signal_2403, LED_128_Instance_state1[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_18_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2356, LED_128_Instance_state0[18]}), .a ({new_AGEMA_signal_3455, new_AGEMA_signal_3451}), .c ({new_AGEMA_signal_2405, LED_128_Instance_state1[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_19_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2270, LED_128_Instance_state0[19]}), .a ({new_AGEMA_signal_3463, new_AGEMA_signal_3459}), .c ({new_AGEMA_signal_2323, LED_128_Instance_state1[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_20_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2271, LED_128_Instance_state0[20]}), .a ({new_AGEMA_signal_3471, new_AGEMA_signal_3467}), .c ({new_AGEMA_signal_2325, LED_128_Instance_state1[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_21_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2311, LED_128_Instance_state0[21]}), .a ({new_AGEMA_signal_3479, new_AGEMA_signal_3475}), .c ({new_AGEMA_signal_2370, LED_128_Instance_state1[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_22_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2357, LED_128_Instance_state0[22]}), .a ({new_AGEMA_signal_3487, new_AGEMA_signal_3483}), .c ({new_AGEMA_signal_2407, LED_128_Instance_state1[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_23_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2272, LED_128_Instance_state0[23]}), .a ({new_AGEMA_signal_3495, new_AGEMA_signal_3491}), .c ({new_AGEMA_signal_2327, LED_128_Instance_state1[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_24_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2273, LED_128_Instance_state0[24]}), .a ({new_AGEMA_signal_3503, new_AGEMA_signal_3499}), .c ({new_AGEMA_signal_2329, LED_128_Instance_state1[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_25_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2312, LED_128_Instance_state0[25]}), .a ({new_AGEMA_signal_3511, new_AGEMA_signal_3507}), .c ({new_AGEMA_signal_2372, LED_128_Instance_state1[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_26_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2313, LED_128_Instance_state0[26]}), .a ({new_AGEMA_signal_3519, new_AGEMA_signal_3515}), .c ({new_AGEMA_signal_2374, LED_128_Instance_state1[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_27_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2274, LED_128_Instance_state0[27]}), .a ({new_AGEMA_signal_3527, new_AGEMA_signal_3523}), .c ({new_AGEMA_signal_2331, LED_128_Instance_state1[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_28_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2314, LED_128_Instance_state0[28]}), .a ({new_AGEMA_signal_3535, new_AGEMA_signal_3531}), .c ({new_AGEMA_signal_2376, LED_128_Instance_state1[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_29_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2358, LED_128_Instance_state0[29]}), .a ({new_AGEMA_signal_3543, new_AGEMA_signal_3539}), .c ({new_AGEMA_signal_2409, LED_128_Instance_state1[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_30_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2315, LED_128_Instance_state0[30]}), .a ({new_AGEMA_signal_3551, new_AGEMA_signal_3547}), .c ({new_AGEMA_signal_2378, LED_128_Instance_state1[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_31_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2275, LED_128_Instance_state0[31]}), .a ({new_AGEMA_signal_3559, new_AGEMA_signal_3555}), .c ({new_AGEMA_signal_2333, LED_128_Instance_state1[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_32_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2359, LED_128_Instance_state0[32]}), .a ({new_AGEMA_signal_3567, new_AGEMA_signal_3563}), .c ({new_AGEMA_signal_2411, LED_128_Instance_state1[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_33_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2395, LED_128_Instance_state0[33]}), .a ({new_AGEMA_signal_3575, new_AGEMA_signal_3571}), .c ({new_AGEMA_signal_2443, LED_128_Instance_state1[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_34_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2360, LED_128_Instance_state0[34]}), .a ({new_AGEMA_signal_3583, new_AGEMA_signal_3579}), .c ({new_AGEMA_signal_2413, LED_128_Instance_state1[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_35_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2435, LED_128_Instance_state0[35]}), .a ({new_AGEMA_signal_3591, new_AGEMA_signal_3587}), .c ({new_AGEMA_signal_2463, LED_128_Instance_state1[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_36_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2361, LED_128_Instance_state0[36]}), .a ({new_AGEMA_signal_3599, new_AGEMA_signal_3595}), .c ({new_AGEMA_signal_2415, LED_128_Instance_state1[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_37_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2362, LED_128_Instance_state0[37]}), .a ({new_AGEMA_signal_3607, new_AGEMA_signal_3603}), .c ({new_AGEMA_signal_2417, LED_128_Instance_state1[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_38_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2316, LED_128_Instance_state0[38]}), .a ({new_AGEMA_signal_3615, new_AGEMA_signal_3611}), .c ({new_AGEMA_signal_2380, LED_128_Instance_state1[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_39_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2436, LED_128_Instance_state0[39]}), .a ({new_AGEMA_signal_3623, new_AGEMA_signal_3619}), .c ({new_AGEMA_signal_2465, LED_128_Instance_state1[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_40_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2363, LED_128_Instance_state0[40]}), .a ({new_AGEMA_signal_3631, new_AGEMA_signal_3627}), .c ({new_AGEMA_signal_2419, LED_128_Instance_state1[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_41_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2364, LED_128_Instance_state0[41]}), .a ({new_AGEMA_signal_3639, new_AGEMA_signal_3635}), .c ({new_AGEMA_signal_2421, LED_128_Instance_state1[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_42_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2317, LED_128_Instance_state0[42]}), .a ({new_AGEMA_signal_3647, new_AGEMA_signal_3643}), .c ({new_AGEMA_signal_2382, LED_128_Instance_state1[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_43_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2396, LED_128_Instance_state0[43]}), .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3651}), .c ({new_AGEMA_signal_2445, LED_128_Instance_state1[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_44_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2365, LED_128_Instance_state0[44]}), .a ({new_AGEMA_signal_3663, new_AGEMA_signal_3659}), .c ({new_AGEMA_signal_2423, LED_128_Instance_state1[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_45_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2397, LED_128_Instance_state0[45]}), .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3667}), .c ({new_AGEMA_signal_2447, LED_128_Instance_state1[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_46_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2366, LED_128_Instance_state0[46]}), .a ({new_AGEMA_signal_3679, new_AGEMA_signal_3675}), .c ({new_AGEMA_signal_2425, LED_128_Instance_state1[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_47_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2398, LED_128_Instance_state0[47]}), .a ({new_AGEMA_signal_3687, new_AGEMA_signal_3683}), .c ({new_AGEMA_signal_2449, LED_128_Instance_state1[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_48_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2492, LED_128_Instance_state0[48]}), .a ({new_AGEMA_signal_3695, new_AGEMA_signal_3691}), .c ({new_AGEMA_signal_2505, LED_128_Instance_state1[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_49_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2502, LED_128_Instance_state0[49]}), .a ({new_AGEMA_signal_3703, new_AGEMA_signal_3699}), .c ({new_AGEMA_signal_2513, LED_128_Instance_state1[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_50_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2437, LED_128_Instance_state0[50]}), .a ({new_AGEMA_signal_3711, new_AGEMA_signal_3707}), .c ({new_AGEMA_signal_2467, LED_128_Instance_state1[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_51_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2438, LED_128_Instance_state0[51]}), .a ({new_AGEMA_signal_3719, new_AGEMA_signal_3715}), .c ({new_AGEMA_signal_2469, LED_128_Instance_state1[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_52_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2493, LED_128_Instance_state0[52]}), .a ({new_AGEMA_signal_3727, new_AGEMA_signal_3723}), .c ({new_AGEMA_signal_2507, LED_128_Instance_state1[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_53_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2503, LED_128_Instance_state0[53]}), .a ({new_AGEMA_signal_3735, new_AGEMA_signal_3731}), .c ({new_AGEMA_signal_2515, LED_128_Instance_state1[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_54_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2399, LED_128_Instance_state0[54]}), .a ({new_AGEMA_signal_3743, new_AGEMA_signal_3739}), .c ({new_AGEMA_signal_2451, LED_128_Instance_state1[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_55_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2439, LED_128_Instance_state0[55]}), .a ({new_AGEMA_signal_3751, new_AGEMA_signal_3747}), .c ({new_AGEMA_signal_2471, LED_128_Instance_state1[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_56_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2484, LED_128_Instance_state0[56]}), .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3755}), .c ({new_AGEMA_signal_2497, LED_128_Instance_state1[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_57_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2494, LED_128_Instance_state0[57]}), .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3763}), .c ({new_AGEMA_signal_2509, LED_128_Instance_state1[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_58_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2400, LED_128_Instance_state0[58]}), .a ({new_AGEMA_signal_3775, new_AGEMA_signal_3771}), .c ({new_AGEMA_signal_2453, LED_128_Instance_state1[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_59_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2401, LED_128_Instance_state0[59]}), .a ({new_AGEMA_signal_3783, new_AGEMA_signal_3779}), .c ({new_AGEMA_signal_2455, LED_128_Instance_state1[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_60_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2485, LED_128_Instance_state0[60]}), .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3787}), .c ({new_AGEMA_signal_2499, LED_128_Instance_state1[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_61_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2495, LED_128_Instance_state0[61]}), .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3795}), .c ({new_AGEMA_signal_2511, LED_128_Instance_state1[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_62_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2440, LED_128_Instance_state0[62]}), .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3803}), .c ({new_AGEMA_signal_2473, LED_128_Instance_state1[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_MUX_state1_mux_inst_63_U1 ( .s (new_AGEMA_signal_3303), .b ({new_AGEMA_signal_2441, LED_128_Instance_state0[63]}), .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3811}), .c ({new_AGEMA_signal_2475, LED_128_Instance_state1[63]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND2_U1 ( .a ({new_AGEMA_signal_1964, LED_128_Instance_SBox_Instance_0_Q2}), .b ({new_AGEMA_signal_3819, new_AGEMA_signal_3817}), .clk (CLK), .r (Fresh[32]), .c ({new_AGEMA_signal_1997, LED_128_Instance_SBox_Instance_0_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_AND4_U1 ( .a ({new_AGEMA_signal_1996, LED_128_Instance_SBox_Instance_0_Q6}), .b ({new_AGEMA_signal_3823, new_AGEMA_signal_3821}), .clk (CLK), .r (Fresh[33]), .c ({new_AGEMA_signal_2028, LED_128_Instance_SBox_Instance_0_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR10_U1 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3825}), .b ({new_AGEMA_signal_2028, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2068, LED_128_Instance_SBox_Instance_0_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR11_U1 ( .a ({new_AGEMA_signal_3835, new_AGEMA_signal_3831}), .b ({new_AGEMA_signal_2068, LED_128_Instance_SBox_Instance_0_L7}), .c ({new_AGEMA_signal_2107, LED_128_Instance_subcells_out[3]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR12_U1 ( .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3825}), .b ({new_AGEMA_signal_1997, LED_128_Instance_SBox_Instance_0_T1}), .c ({new_AGEMA_signal_2029, LED_128_Instance_SBox_Instance_0_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR13_U1 ( .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3839}), .b ({new_AGEMA_signal_2029, LED_128_Instance_SBox_Instance_0_L8}), .c ({new_AGEMA_signal_2069, LED_128_Instance_subcells_out[2]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_0_XOR14_U1 ( .a ({new_AGEMA_signal_3847, new_AGEMA_signal_3845}), .b ({new_AGEMA_signal_2028, LED_128_Instance_SBox_Instance_0_T3}), .c ({new_AGEMA_signal_2070, LED_128_Instance_subcells_out[1]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND2_U1 ( .a ({new_AGEMA_signal_1966, LED_128_Instance_SBox_Instance_1_Q2}), .b ({new_AGEMA_signal_3851, new_AGEMA_signal_3849}), .clk (CLK), .r (Fresh[34]), .c ({new_AGEMA_signal_1999, LED_128_Instance_SBox_Instance_1_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_AND4_U1 ( .a ({new_AGEMA_signal_1998, LED_128_Instance_SBox_Instance_1_Q6}), .b ({new_AGEMA_signal_3855, new_AGEMA_signal_3853}), .clk (CLK), .r (Fresh[35]), .c ({new_AGEMA_signal_2030, LED_128_Instance_SBox_Instance_1_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR10_U1 ( .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3857}), .b ({new_AGEMA_signal_2030, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2071, LED_128_Instance_SBox_Instance_1_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR11_U1 ( .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3863}), .b ({new_AGEMA_signal_2071, LED_128_Instance_SBox_Instance_1_L7}), .c ({new_AGEMA_signal_2108, LED_128_Instance_subcells_out[7]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR12_U1 ( .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3857}), .b ({new_AGEMA_signal_1999, LED_128_Instance_SBox_Instance_1_T1}), .c ({new_AGEMA_signal_2031, LED_128_Instance_SBox_Instance_1_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR13_U1 ( .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3871}), .b ({new_AGEMA_signal_2031, LED_128_Instance_SBox_Instance_1_L8}), .c ({new_AGEMA_signal_2072, LED_128_Instance_subcells_out[6]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_1_XOR14_U1 ( .a ({new_AGEMA_signal_3879, new_AGEMA_signal_3877}), .b ({new_AGEMA_signal_2030, LED_128_Instance_SBox_Instance_1_T3}), .c ({new_AGEMA_signal_2073, LED_128_Instance_subcells_out[5]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND2_U1 ( .a ({new_AGEMA_signal_1936, LED_128_Instance_SBox_Instance_2_Q2}), .b ({new_AGEMA_signal_3883, new_AGEMA_signal_3881}), .clk (CLK), .r (Fresh[36]), .c ({new_AGEMA_signal_1969, LED_128_Instance_SBox_Instance_2_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_AND4_U1 ( .a ({new_AGEMA_signal_1968, LED_128_Instance_SBox_Instance_2_Q6}), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3885}), .clk (CLK), .r (Fresh[37]), .c ({new_AGEMA_signal_2000, LED_128_Instance_SBox_Instance_2_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR10_U1 ( .a ({new_AGEMA_signal_3891, new_AGEMA_signal_3889}), .b ({new_AGEMA_signal_2000, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2032, LED_128_Instance_SBox_Instance_2_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR11_U1 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2851}), .b ({new_AGEMA_signal_2032, LED_128_Instance_SBox_Instance_2_L7}), .c ({new_AGEMA_signal_2074, LED_128_Instance_subcells_out[11]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR12_U1 ( .a ({new_AGEMA_signal_3891, new_AGEMA_signal_3889}), .b ({new_AGEMA_signal_1969, LED_128_Instance_SBox_Instance_2_T1}), .c ({new_AGEMA_signal_2001, LED_128_Instance_SBox_Instance_2_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR13_U1 ( .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3895}), .b ({new_AGEMA_signal_2001, LED_128_Instance_SBox_Instance_2_L8}), .c ({new_AGEMA_signal_2033, LED_128_Instance_subcells_out[10]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_2_XOR14_U1 ( .a ({new_AGEMA_signal_3903, new_AGEMA_signal_3901}), .b ({new_AGEMA_signal_2000, LED_128_Instance_SBox_Instance_2_T3}), .c ({new_AGEMA_signal_2034, LED_128_Instance_subcells_out[9]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND2_U1 ( .a ({new_AGEMA_signal_1938, LED_128_Instance_SBox_Instance_3_Q2}), .b ({new_AGEMA_signal_3907, new_AGEMA_signal_3905}), .clk (CLK), .r (Fresh[38]), .c ({new_AGEMA_signal_1971, LED_128_Instance_SBox_Instance_3_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_AND4_U1 ( .a ({new_AGEMA_signal_1970, LED_128_Instance_SBox_Instance_3_Q6}), .b ({new_AGEMA_signal_3911, new_AGEMA_signal_3909}), .clk (CLK), .r (Fresh[39]), .c ({new_AGEMA_signal_2002, LED_128_Instance_SBox_Instance_3_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR10_U1 ( .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3913}), .b ({new_AGEMA_signal_2002, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2035, LED_128_Instance_SBox_Instance_3_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR11_U1 ( .a ({new_AGEMA_signal_2887, new_AGEMA_signal_2883}), .b ({new_AGEMA_signal_2035, LED_128_Instance_SBox_Instance_3_L7}), .c ({new_AGEMA_signal_2075, LED_128_Instance_subcells_out[15]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR12_U1 ( .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3913}), .b ({new_AGEMA_signal_1971, LED_128_Instance_SBox_Instance_3_T1}), .c ({new_AGEMA_signal_2003, LED_128_Instance_SBox_Instance_3_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR13_U1 ( .a ({new_AGEMA_signal_3923, new_AGEMA_signal_3919}), .b ({new_AGEMA_signal_2003, LED_128_Instance_SBox_Instance_3_L8}), .c ({new_AGEMA_signal_2036, LED_128_Instance_subcells_out[14]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_3_XOR14_U1 ( .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3925}), .b ({new_AGEMA_signal_2002, LED_128_Instance_SBox_Instance_3_T3}), .c ({new_AGEMA_signal_2037, LED_128_Instance_subcells_out[13]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND2_U1 ( .a ({new_AGEMA_signal_1972, LED_128_Instance_SBox_Instance_4_Q2}), .b ({new_AGEMA_signal_3931, new_AGEMA_signal_3929}), .clk (CLK), .r (Fresh[40]), .c ({new_AGEMA_signal_2005, LED_128_Instance_SBox_Instance_4_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_AND4_U1 ( .a ({new_AGEMA_signal_2004, LED_128_Instance_SBox_Instance_4_Q6}), .b ({new_AGEMA_signal_3935, new_AGEMA_signal_3933}), .clk (CLK), .r (Fresh[41]), .c ({new_AGEMA_signal_2038, LED_128_Instance_SBox_Instance_4_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR10_U1 ( .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3937}), .b ({new_AGEMA_signal_2038, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2076, LED_128_Instance_SBox_Instance_4_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR11_U1 ( .a ({new_AGEMA_signal_3947, new_AGEMA_signal_3943}), .b ({new_AGEMA_signal_2076, LED_128_Instance_SBox_Instance_4_L7}), .c ({new_AGEMA_signal_2109, LED_128_Instance_subcells_out[19]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR12_U1 ( .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3937}), .b ({new_AGEMA_signal_2005, LED_128_Instance_SBox_Instance_4_T1}), .c ({new_AGEMA_signal_2039, LED_128_Instance_SBox_Instance_4_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR13_U1 ( .a ({new_AGEMA_signal_3955, new_AGEMA_signal_3951}), .b ({new_AGEMA_signal_2039, LED_128_Instance_SBox_Instance_4_L8}), .c ({new_AGEMA_signal_2077, LED_128_Instance_subcells_out[18]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_4_XOR14_U1 ( .a ({new_AGEMA_signal_3959, new_AGEMA_signal_3957}), .b ({new_AGEMA_signal_2038, LED_128_Instance_SBox_Instance_4_T3}), .c ({new_AGEMA_signal_2078, LED_128_Instance_subcells_out[17]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND2_U1 ( .a ({new_AGEMA_signal_1974, LED_128_Instance_SBox_Instance_5_Q2}), .b ({new_AGEMA_signal_3963, new_AGEMA_signal_3961}), .clk (CLK), .r (Fresh[42]), .c ({new_AGEMA_signal_2007, LED_128_Instance_SBox_Instance_5_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_AND4_U1 ( .a ({new_AGEMA_signal_2006, LED_128_Instance_SBox_Instance_5_Q6}), .b ({new_AGEMA_signal_3967, new_AGEMA_signal_3965}), .clk (CLK), .r (Fresh[43]), .c ({new_AGEMA_signal_2040, LED_128_Instance_SBox_Instance_5_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR10_U1 ( .a ({new_AGEMA_signal_3971, new_AGEMA_signal_3969}), .b ({new_AGEMA_signal_2040, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2079, LED_128_Instance_SBox_Instance_5_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR11_U1 ( .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3975}), .b ({new_AGEMA_signal_2079, LED_128_Instance_SBox_Instance_5_L7}), .c ({new_AGEMA_signal_2110, LED_128_Instance_subcells_out[23]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR12_U1 ( .a ({new_AGEMA_signal_3971, new_AGEMA_signal_3969}), .b ({new_AGEMA_signal_2007, LED_128_Instance_SBox_Instance_5_T1}), .c ({new_AGEMA_signal_2041, LED_128_Instance_SBox_Instance_5_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR13_U1 ( .a ({new_AGEMA_signal_3987, new_AGEMA_signal_3983}), .b ({new_AGEMA_signal_2041, LED_128_Instance_SBox_Instance_5_L8}), .c ({new_AGEMA_signal_2080, LED_128_Instance_subcells_out[22]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_5_XOR14_U1 ( .a ({new_AGEMA_signal_3991, new_AGEMA_signal_3989}), .b ({new_AGEMA_signal_2040, LED_128_Instance_SBox_Instance_5_T3}), .c ({new_AGEMA_signal_2081, LED_128_Instance_subcells_out[21]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND2_U1 ( .a ({new_AGEMA_signal_1944, LED_128_Instance_SBox_Instance_6_Q2}), .b ({new_AGEMA_signal_3995, new_AGEMA_signal_3993}), .clk (CLK), .r (Fresh[44]), .c ({new_AGEMA_signal_1977, LED_128_Instance_SBox_Instance_6_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_AND4_U1 ( .a ({new_AGEMA_signal_1976, LED_128_Instance_SBox_Instance_6_Q6}), .b ({new_AGEMA_signal_3999, new_AGEMA_signal_3997}), .clk (CLK), .r (Fresh[45]), .c ({new_AGEMA_signal_2008, LED_128_Instance_SBox_Instance_6_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR10_U1 ( .a ({new_AGEMA_signal_4003, new_AGEMA_signal_4001}), .b ({new_AGEMA_signal_2008, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2042, LED_128_Instance_SBox_Instance_6_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR11_U1 ( .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2979}), .b ({new_AGEMA_signal_2042, LED_128_Instance_SBox_Instance_6_L7}), .c ({new_AGEMA_signal_2082, LED_128_Instance_subcells_out[27]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR12_U1 ( .a ({new_AGEMA_signal_4003, new_AGEMA_signal_4001}), .b ({new_AGEMA_signal_1977, LED_128_Instance_SBox_Instance_6_T1}), .c ({new_AGEMA_signal_2009, LED_128_Instance_SBox_Instance_6_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR13_U1 ( .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4007}), .b ({new_AGEMA_signal_2009, LED_128_Instance_SBox_Instance_6_L8}), .c ({new_AGEMA_signal_2043, LED_128_Instance_subcells_out[26]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_6_XOR14_U1 ( .a ({new_AGEMA_signal_4015, new_AGEMA_signal_4013}), .b ({new_AGEMA_signal_2008, LED_128_Instance_SBox_Instance_6_T3}), .c ({new_AGEMA_signal_2044, LED_128_Instance_subcells_out[25]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND2_U1 ( .a ({new_AGEMA_signal_1946, LED_128_Instance_SBox_Instance_7_Q2}), .b ({new_AGEMA_signal_4019, new_AGEMA_signal_4017}), .clk (CLK), .r (Fresh[46]), .c ({new_AGEMA_signal_1979, LED_128_Instance_SBox_Instance_7_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_AND4_U1 ( .a ({new_AGEMA_signal_1978, LED_128_Instance_SBox_Instance_7_Q6}), .b ({new_AGEMA_signal_4023, new_AGEMA_signal_4021}), .clk (CLK), .r (Fresh[47]), .c ({new_AGEMA_signal_2010, LED_128_Instance_SBox_Instance_7_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR10_U1 ( .a ({new_AGEMA_signal_4027, new_AGEMA_signal_4025}), .b ({new_AGEMA_signal_2010, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2045, LED_128_Instance_SBox_Instance_7_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR11_U1 ( .a ({new_AGEMA_signal_3015, new_AGEMA_signal_3011}), .b ({new_AGEMA_signal_2045, LED_128_Instance_SBox_Instance_7_L7}), .c ({new_AGEMA_signal_2083, LED_128_Instance_subcells_out[31]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR12_U1 ( .a ({new_AGEMA_signal_4027, new_AGEMA_signal_4025}), .b ({new_AGEMA_signal_1979, LED_128_Instance_SBox_Instance_7_T1}), .c ({new_AGEMA_signal_2011, LED_128_Instance_SBox_Instance_7_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR13_U1 ( .a ({new_AGEMA_signal_4035, new_AGEMA_signal_4031}), .b ({new_AGEMA_signal_2011, LED_128_Instance_SBox_Instance_7_L8}), .c ({new_AGEMA_signal_2046, LED_128_Instance_subcells_out[30]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_7_XOR14_U1 ( .a ({new_AGEMA_signal_4039, new_AGEMA_signal_4037}), .b ({new_AGEMA_signal_2010, LED_128_Instance_SBox_Instance_7_T3}), .c ({new_AGEMA_signal_2047, LED_128_Instance_subcells_out[29]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND2_U1 ( .a ({new_AGEMA_signal_1980, LED_128_Instance_SBox_Instance_8_Q2}), .b ({new_AGEMA_signal_4043, new_AGEMA_signal_4041}), .clk (CLK), .r (Fresh[48]), .c ({new_AGEMA_signal_2013, LED_128_Instance_SBox_Instance_8_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_AND4_U1 ( .a ({new_AGEMA_signal_2012, LED_128_Instance_SBox_Instance_8_Q6}), .b ({new_AGEMA_signal_4047, new_AGEMA_signal_4045}), .clk (CLK), .r (Fresh[49]), .c ({new_AGEMA_signal_2048, LED_128_Instance_SBox_Instance_8_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR10_U1 ( .a ({new_AGEMA_signal_4051, new_AGEMA_signal_4049}), .b ({new_AGEMA_signal_2048, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2084, LED_128_Instance_SBox_Instance_8_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR11_U1 ( .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4055}), .b ({new_AGEMA_signal_2084, LED_128_Instance_SBox_Instance_8_L7}), .c ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR12_U1 ( .a ({new_AGEMA_signal_4051, new_AGEMA_signal_4049}), .b ({new_AGEMA_signal_2013, LED_128_Instance_SBox_Instance_8_T1}), .c ({new_AGEMA_signal_2049, LED_128_Instance_SBox_Instance_8_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR13_U1 ( .a ({new_AGEMA_signal_4067, new_AGEMA_signal_4063}), .b ({new_AGEMA_signal_2049, LED_128_Instance_SBox_Instance_8_L8}), .c ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_8_XOR14_U1 ( .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4069}), .b ({new_AGEMA_signal_2048, LED_128_Instance_SBox_Instance_8_T3}), .c ({new_AGEMA_signal_2086, LED_128_Instance_subcells_out[33]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND2_U1 ( .a ({new_AGEMA_signal_1982, LED_128_Instance_SBox_Instance_9_Q2}), .b ({new_AGEMA_signal_4075, new_AGEMA_signal_4073}), .clk (CLK), .r (Fresh[50]), .c ({new_AGEMA_signal_2015, LED_128_Instance_SBox_Instance_9_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_AND4_U1 ( .a ({new_AGEMA_signal_2014, LED_128_Instance_SBox_Instance_9_Q6}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4077}), .clk (CLK), .r (Fresh[51]), .c ({new_AGEMA_signal_2050, LED_128_Instance_SBox_Instance_9_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR10_U1 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4081}), .b ({new_AGEMA_signal_2050, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2087, LED_128_Instance_SBox_Instance_9_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR11_U1 ( .a ({new_AGEMA_signal_4091, new_AGEMA_signal_4087}), .b ({new_AGEMA_signal_2087, LED_128_Instance_SBox_Instance_9_L7}), .c ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR12_U1 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4081}), .b ({new_AGEMA_signal_2015, LED_128_Instance_SBox_Instance_9_T1}), .c ({new_AGEMA_signal_2051, LED_128_Instance_SBox_Instance_9_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR13_U1 ( .a ({new_AGEMA_signal_4099, new_AGEMA_signal_4095}), .b ({new_AGEMA_signal_2051, LED_128_Instance_SBox_Instance_9_L8}), .c ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_9_XOR14_U1 ( .a ({new_AGEMA_signal_4103, new_AGEMA_signal_4101}), .b ({new_AGEMA_signal_2050, LED_128_Instance_SBox_Instance_9_T3}), .c ({new_AGEMA_signal_2089, LED_128_Instance_subcells_out[37]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND2_U1 ( .a ({new_AGEMA_signal_1952, LED_128_Instance_SBox_Instance_10_Q2}), .b ({new_AGEMA_signal_4107, new_AGEMA_signal_4105}), .clk (CLK), .r (Fresh[52]), .c ({new_AGEMA_signal_1985, LED_128_Instance_SBox_Instance_10_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_AND4_U1 ( .a ({new_AGEMA_signal_1984, LED_128_Instance_SBox_Instance_10_Q6}), .b ({new_AGEMA_signal_4111, new_AGEMA_signal_4109}), .clk (CLK), .r (Fresh[53]), .c ({new_AGEMA_signal_2016, LED_128_Instance_SBox_Instance_10_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR10_U1 ( .a ({new_AGEMA_signal_4115, new_AGEMA_signal_4113}), .b ({new_AGEMA_signal_2016, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2052, LED_128_Instance_SBox_Instance_10_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR11_U1 ( .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3107}), .b ({new_AGEMA_signal_2052, LED_128_Instance_SBox_Instance_10_L7}), .c ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR12_U1 ( .a ({new_AGEMA_signal_4115, new_AGEMA_signal_4113}), .b ({new_AGEMA_signal_1985, LED_128_Instance_SBox_Instance_10_T1}), .c ({new_AGEMA_signal_2017, LED_128_Instance_SBox_Instance_10_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR13_U1 ( .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4119}), .b ({new_AGEMA_signal_2017, LED_128_Instance_SBox_Instance_10_L8}), .c ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_10_XOR14_U1 ( .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4125}), .b ({new_AGEMA_signal_2016, LED_128_Instance_SBox_Instance_10_T3}), .c ({new_AGEMA_signal_2054, LED_128_Instance_subcells_out[41]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND2_U1 ( .a ({new_AGEMA_signal_1954, LED_128_Instance_SBox_Instance_11_Q2}), .b ({new_AGEMA_signal_4131, new_AGEMA_signal_4129}), .clk (CLK), .r (Fresh[54]), .c ({new_AGEMA_signal_1987, LED_128_Instance_SBox_Instance_11_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_AND4_U1 ( .a ({new_AGEMA_signal_1986, LED_128_Instance_SBox_Instance_11_Q6}), .b ({new_AGEMA_signal_4135, new_AGEMA_signal_4133}), .clk (CLK), .r (Fresh[55]), .c ({new_AGEMA_signal_2018, LED_128_Instance_SBox_Instance_11_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR10_U1 ( .a ({new_AGEMA_signal_4139, new_AGEMA_signal_4137}), .b ({new_AGEMA_signal_2018, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2055, LED_128_Instance_SBox_Instance_11_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR11_U1 ( .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3143}), .b ({new_AGEMA_signal_2055, LED_128_Instance_SBox_Instance_11_L7}), .c ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR12_U1 ( .a ({new_AGEMA_signal_4139, new_AGEMA_signal_4137}), .b ({new_AGEMA_signal_1987, LED_128_Instance_SBox_Instance_11_T1}), .c ({new_AGEMA_signal_2019, LED_128_Instance_SBox_Instance_11_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR13_U1 ( .a ({new_AGEMA_signal_4147, new_AGEMA_signal_4143}), .b ({new_AGEMA_signal_2019, LED_128_Instance_SBox_Instance_11_L8}), .c ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_11_XOR14_U1 ( .a ({new_AGEMA_signal_4151, new_AGEMA_signal_4149}), .b ({new_AGEMA_signal_2018, LED_128_Instance_SBox_Instance_11_T3}), .c ({new_AGEMA_signal_2057, LED_128_Instance_subcells_out[45]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND2_U1 ( .a ({new_AGEMA_signal_1988, LED_128_Instance_SBox_Instance_12_Q2}), .b ({new_AGEMA_signal_4155, new_AGEMA_signal_4153}), .clk (CLK), .r (Fresh[56]), .c ({new_AGEMA_signal_2021, LED_128_Instance_SBox_Instance_12_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_AND4_U1 ( .a ({new_AGEMA_signal_2020, LED_128_Instance_SBox_Instance_12_Q6}), .b ({new_AGEMA_signal_4159, new_AGEMA_signal_4157}), .clk (CLK), .r (Fresh[57]), .c ({new_AGEMA_signal_2058, LED_128_Instance_SBox_Instance_12_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR10_U1 ( .a ({new_AGEMA_signal_4163, new_AGEMA_signal_4161}), .b ({new_AGEMA_signal_2058, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2092, LED_128_Instance_SBox_Instance_12_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR11_U1 ( .a ({new_AGEMA_signal_4171, new_AGEMA_signal_4167}), .b ({new_AGEMA_signal_2092, LED_128_Instance_SBox_Instance_12_L7}), .c ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR12_U1 ( .a ({new_AGEMA_signal_4163, new_AGEMA_signal_4161}), .b ({new_AGEMA_signal_2021, LED_128_Instance_SBox_Instance_12_T1}), .c ({new_AGEMA_signal_2059, LED_128_Instance_SBox_Instance_12_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR13_U1 ( .a ({new_AGEMA_signal_4179, new_AGEMA_signal_4175}), .b ({new_AGEMA_signal_2059, LED_128_Instance_SBox_Instance_12_L8}), .c ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_12_XOR14_U1 ( .a ({new_AGEMA_signal_4183, new_AGEMA_signal_4181}), .b ({new_AGEMA_signal_2058, LED_128_Instance_SBox_Instance_12_T3}), .c ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND2_U1 ( .a ({new_AGEMA_signal_1990, LED_128_Instance_SBox_Instance_13_Q2}), .b ({new_AGEMA_signal_4187, new_AGEMA_signal_4185}), .clk (CLK), .r (Fresh[58]), .c ({new_AGEMA_signal_2023, LED_128_Instance_SBox_Instance_13_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_AND4_U1 ( .a ({new_AGEMA_signal_2022, LED_128_Instance_SBox_Instance_13_Q6}), .b ({new_AGEMA_signal_4191, new_AGEMA_signal_4189}), .clk (CLK), .r (Fresh[59]), .c ({new_AGEMA_signal_2060, LED_128_Instance_SBox_Instance_13_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR10_U1 ( .a ({new_AGEMA_signal_4195, new_AGEMA_signal_4193}), .b ({new_AGEMA_signal_2060, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2095, LED_128_Instance_SBox_Instance_13_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR11_U1 ( .a ({new_AGEMA_signal_4203, new_AGEMA_signal_4199}), .b ({new_AGEMA_signal_2095, LED_128_Instance_SBox_Instance_13_L7}), .c ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR12_U1 ( .a ({new_AGEMA_signal_4195, new_AGEMA_signal_4193}), .b ({new_AGEMA_signal_2023, LED_128_Instance_SBox_Instance_13_T1}), .c ({new_AGEMA_signal_2061, LED_128_Instance_SBox_Instance_13_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR13_U1 ( .a ({new_AGEMA_signal_4211, new_AGEMA_signal_4207}), .b ({new_AGEMA_signal_2061, LED_128_Instance_SBox_Instance_13_L8}), .c ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_13_XOR14_U1 ( .a ({new_AGEMA_signal_4215, new_AGEMA_signal_4213}), .b ({new_AGEMA_signal_2060, LED_128_Instance_SBox_Instance_13_T3}), .c ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND2_U1 ( .a ({new_AGEMA_signal_1960, LED_128_Instance_SBox_Instance_14_Q2}), .b ({new_AGEMA_signal_4219, new_AGEMA_signal_4217}), .clk (CLK), .r (Fresh[60]), .c ({new_AGEMA_signal_1993, LED_128_Instance_SBox_Instance_14_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_AND4_U1 ( .a ({new_AGEMA_signal_1992, LED_128_Instance_SBox_Instance_14_Q6}), .b ({new_AGEMA_signal_4223, new_AGEMA_signal_4221}), .clk (CLK), .r (Fresh[61]), .c ({new_AGEMA_signal_2024, LED_128_Instance_SBox_Instance_14_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR10_U1 ( .a ({new_AGEMA_signal_4227, new_AGEMA_signal_4225}), .b ({new_AGEMA_signal_2024, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2062, LED_128_Instance_SBox_Instance_14_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR11_U1 ( .a ({new_AGEMA_signal_3243, new_AGEMA_signal_3239}), .b ({new_AGEMA_signal_2062, LED_128_Instance_SBox_Instance_14_L7}), .c ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR12_U1 ( .a ({new_AGEMA_signal_4227, new_AGEMA_signal_4225}), .b ({new_AGEMA_signal_1993, LED_128_Instance_SBox_Instance_14_T1}), .c ({new_AGEMA_signal_2025, LED_128_Instance_SBox_Instance_14_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR13_U1 ( .a ({new_AGEMA_signal_4235, new_AGEMA_signal_4231}), .b ({new_AGEMA_signal_2025, LED_128_Instance_SBox_Instance_14_L8}), .c ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_14_XOR14_U1 ( .a ({new_AGEMA_signal_4239, new_AGEMA_signal_4237}), .b ({new_AGEMA_signal_2024, LED_128_Instance_SBox_Instance_14_T3}), .c ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND2_U1 ( .a ({new_AGEMA_signal_1962, LED_128_Instance_SBox_Instance_15_Q2}), .b ({new_AGEMA_signal_4243, new_AGEMA_signal_4241}), .clk (CLK), .r (Fresh[62]), .c ({new_AGEMA_signal_1995, LED_128_Instance_SBox_Instance_15_T1}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_AND4_U1 ( .a ({new_AGEMA_signal_1994, LED_128_Instance_SBox_Instance_15_Q6}), .b ({new_AGEMA_signal_4247, new_AGEMA_signal_4245}), .clk (CLK), .r (Fresh[63]), .c ({new_AGEMA_signal_2026, LED_128_Instance_SBox_Instance_15_T3}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR10_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4249}), .b ({new_AGEMA_signal_2026, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2065, LED_128_Instance_SBox_Instance_15_L7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR11_U1 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3271}), .b ({new_AGEMA_signal_2065, LED_128_Instance_SBox_Instance_15_L7}), .c ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR12_U1 ( .a ({new_AGEMA_signal_4251, new_AGEMA_signal_4249}), .b ({new_AGEMA_signal_1995, LED_128_Instance_SBox_Instance_15_T1}), .c ({new_AGEMA_signal_2027, LED_128_Instance_SBox_Instance_15_L8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR13_U1 ( .a ({new_AGEMA_signal_4259, new_AGEMA_signal_4255}), .b ({new_AGEMA_signal_2027, LED_128_Instance_SBox_Instance_15_L8}), .c ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_SBox_Instance_15_XOR14_U1 ( .a ({new_AGEMA_signal_4263, new_AGEMA_signal_4261}), .b ({new_AGEMA_signal_2026, LED_128_Instance_SBox_Instance_15_T3}), .c ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U54 ( .a ({new_AGEMA_signal_2383, LED_128_Instance_MCS_Instance_0_n38}), .b ({new_AGEMA_signal_2244, LED_128_Instance_MCS_Instance_0_n37}), .c ({new_AGEMA_signal_2426, LED_128_Instance_mixcolumns_out[51]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U53 ( .a ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2244, LED_128_Instance_MCS_Instance_0_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U52 ( .a ({new_AGEMA_signal_2334, LED_128_Instance_mixcolumns_out[34]}), .b ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}), .c ({new_AGEMA_signal_2383, LED_128_Instance_MCS_Instance_0_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U51 ( .a ({new_AGEMA_signal_2202, LED_128_Instance_MCS_Instance_0_n36}), .b ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_2334, LED_128_Instance_mixcolumns_out[34]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U50 ( .a ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2173, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_2202, LED_128_Instance_MCS_Instance_0_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U49 ( .a ({new_AGEMA_signal_2335, LED_128_Instance_MCS_Instance_0_n33}), .b ({new_AGEMA_signal_2385, LED_128_Instance_mixcolumns_out[33]}), .c ({new_AGEMA_signal_2427, LED_128_Instance_mixcolumns_out[50]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U48 ( .a ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_2335, LED_128_Instance_MCS_Instance_0_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U47 ( .a ({new_AGEMA_signal_2486, LED_128_Instance_MCS_Instance_0_n32}), .b ({new_AGEMA_signal_2338, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_2500, LED_128_Instance_mixcolumns_out[49]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U46 ( .a ({new_AGEMA_signal_2476, LED_128_Instance_MCS_Instance_0_n30}), .b ({new_AGEMA_signal_2284, LED_128_Instance_MCS_Instance_0_n29}), .c ({new_AGEMA_signal_2486, LED_128_Instance_MCS_Instance_0_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U45 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}), .c ({new_AGEMA_signal_2284, LED_128_Instance_MCS_Instance_0_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U44 ( .a ({new_AGEMA_signal_2336, LED_128_Instance_mixcolumns_out[32]}), .b ({new_AGEMA_signal_2456, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_2476, LED_128_Instance_MCS_Instance_0_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U43 ( .a ({new_AGEMA_signal_2285, LED_128_Instance_MCS_Instance_0_n27}), .b ({new_AGEMA_signal_2245, LED_128_Instance_MCS_Instance_0_n26}), .c ({new_AGEMA_signal_2336, LED_128_Instance_mixcolumns_out[32]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U42 ( .a ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .c ({new_AGEMA_signal_2245, LED_128_Instance_MCS_Instance_0_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U41 ( .a ({new_AGEMA_signal_4267, new_AGEMA_signal_4265}), .b ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_2285, LED_128_Instance_MCS_Instance_0_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U40 ( .a ({new_AGEMA_signal_2477, LED_128_Instance_MCS_Instance_0_n25}), .b ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_2487, LED_128_Instance_mixcolumns_out[48]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U39 ( .a ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .b ({new_AGEMA_signal_2456, LED_128_Instance_MCS_Instance_0_n28}), .c ({new_AGEMA_signal_2477, LED_128_Instance_MCS_Instance_0_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U38 ( .a ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2428, LED_128_Instance_mixcolumns_out[35]}), .c ({new_AGEMA_signal_2456, LED_128_Instance_MCS_Instance_0_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U37 ( .a ({new_AGEMA_signal_2384, LED_128_Instance_MCS_Instance_0_n24}), .b ({new_AGEMA_signal_2115, LED_128_Instance_MCS_Instance_0_n23}), .c ({new_AGEMA_signal_2428, LED_128_Instance_mixcolumns_out[35]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U36 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2054, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2115, LED_128_Instance_MCS_Instance_0_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U35 ( .a ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}), .b ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .c ({new_AGEMA_signal_2384, LED_128_Instance_MCS_Instance_0_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U34 ( .a ({new_AGEMA_signal_2286, LED_128_Instance_MCS_Instance_0_n22}), .b ({new_AGEMA_signal_2172, LED_128_Instance_MCS_Instance_0_n21}), .c ({new_AGEMA_signal_2337, LED_128_Instance_mixcolumns_out[18]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U33 ( .a ({new_AGEMA_signal_2144, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2172, LED_128_Instance_MCS_Instance_0_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U32 ( .a ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}), .b ({new_AGEMA_signal_4271, new_AGEMA_signal_4269}), .c ({new_AGEMA_signal_2286, LED_128_Instance_MCS_Instance_0_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U31 ( .a ({new_AGEMA_signal_2203, LED_128_Instance_MCS_Instance_0_n19}), .b ({new_AGEMA_signal_2116, LED_128_Instance_MCS_Instance_0_n18}), .c ({new_AGEMA_signal_2246, LED_128_Instance_mixcolumns_out[1]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U30 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4273}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2116, LED_128_Instance_MCS_Instance_0_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U29 ( .a ({new_AGEMA_signal_2121, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_2173, LED_128_Instance_MCS_Instance_0_n34}), .c ({new_AGEMA_signal_2203, LED_128_Instance_MCS_Instance_0_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U28 ( .a ({new_AGEMA_signal_2140, LED_128_Instance_MCS_Instance_0_n16}), .b ({new_AGEMA_signal_2069, LED_128_Instance_subcells_out[2]}), .c ({new_AGEMA_signal_2173, LED_128_Instance_MCS_Instance_0_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U27 ( .a ({new_AGEMA_signal_2081, LED_128_Instance_subcells_out[21]}), .b ({new_AGEMA_signal_2107, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2140, LED_128_Instance_MCS_Instance_0_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U26 ( .a ({new_AGEMA_signal_2339, LED_128_Instance_MCS_Instance_0_n15}), .b ({new_AGEMA_signal_2338, LED_128_Instance_MCS_Instance_0_n31}), .c ({new_AGEMA_signal_2385, LED_128_Instance_mixcolumns_out[33]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U25 ( .a ({new_AGEMA_signal_2288, LED_128_Instance_mixcolumns_out[16]}), .b ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}), .c ({new_AGEMA_signal_2338, LED_128_Instance_MCS_Instance_0_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U24 ( .a ({new_AGEMA_signal_2287, LED_128_Instance_MCS_Instance_0_n14}), .b ({new_AGEMA_signal_2117, LED_128_Instance_MCS_Instance_0_n13}), .c ({new_AGEMA_signal_2339, LED_128_Instance_MCS_Instance_0_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U23 ( .a ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2117, LED_128_Instance_MCS_Instance_0_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U22 ( .a ({new_AGEMA_signal_2249, LED_128_Instance_MCS_Instance_0_n12}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2287, LED_128_Instance_MCS_Instance_0_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U21 ( .a ({new_AGEMA_signal_2118, LED_128_Instance_MCS_Instance_0_n11}), .b ({new_AGEMA_signal_2247, LED_128_Instance_MCS_Instance_0_n10}), .c ({new_AGEMA_signal_2288, LED_128_Instance_mixcolumns_out[16]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U20 ( .a ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .c ({new_AGEMA_signal_2247, LED_128_Instance_MCS_Instance_0_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U19 ( .a ({new_AGEMA_signal_4275, new_AGEMA_signal_4273}), .b ({new_AGEMA_signal_2080, LED_128_Instance_subcells_out[22]}), .c ({new_AGEMA_signal_2118, LED_128_Instance_MCS_Instance_0_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U18 ( .a ({new_AGEMA_signal_2204, LED_128_Instance_MCS_Instance_0_n9}), .b ({new_AGEMA_signal_2119, LED_128_Instance_MCS_Instance_0_n8}), .c ({new_AGEMA_signal_2248, LED_128_Instance_mixcolumns_out[19]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U17 ( .a ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2119, LED_128_Instance_MCS_Instance_0_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U16 ( .a ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}), .b ({new_AGEMA_signal_2081, LED_128_Instance_subcells_out[21]}), .c ({new_AGEMA_signal_2204, LED_128_Instance_MCS_Instance_0_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U15 ( .a ({new_AGEMA_signal_2100, LED_128_Instance_MCS_Instance_0_n7}), .b ({new_AGEMA_signal_2141, LED_128_Instance_MCS_Instance_0_n6}), .c ({new_AGEMA_signal_2174, LED_128_Instance_mixcolumns_out[2]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U14 ( .a ({new_AGEMA_signal_2120, LED_128_Instance_MCS_Instance_0_n5}), .b ({new_AGEMA_signal_2107, LED_128_Instance_subcells_out[3]}), .c ({new_AGEMA_signal_2141, LED_128_Instance_MCS_Instance_0_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U13 ( .a ({new_AGEMA_signal_4279, new_AGEMA_signal_4277}), .b ({new_AGEMA_signal_2067, LED_128_Instance_subcells_out[61]}), .c ({new_AGEMA_signal_2100, LED_128_Instance_MCS_Instance_0_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U12 ( .a ({new_AGEMA_signal_2121, LED_128_Instance_MCS_Instance_0_n17}), .b ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}), .c ({new_AGEMA_signal_2340, LED_128_Instance_mixcolumns_out[17]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U11 ( .a ({new_AGEMA_signal_2142, LED_128_Instance_MCS_Instance_0_n4}), .b ({new_AGEMA_signal_2249, LED_128_Instance_MCS_Instance_0_n12}), .c ({new_AGEMA_signal_2289, LED_128_Instance_MCS_Instance_0_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U10 ( .a ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}), .b ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}), .c ({new_AGEMA_signal_2249, LED_128_Instance_MCS_Instance_0_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U9 ( .a ({new_AGEMA_signal_2110, LED_128_Instance_subcells_out[23]}), .b ({new_AGEMA_signal_2120, LED_128_Instance_MCS_Instance_0_n5}), .c ({new_AGEMA_signal_2142, LED_128_Instance_MCS_Instance_0_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U8 ( .a ({new_AGEMA_signal_2080, LED_128_Instance_subcells_out[22]}), .b ({new_AGEMA_signal_2054, LED_128_Instance_subcells_out[41]}), .c ({new_AGEMA_signal_2120, LED_128_Instance_MCS_Instance_0_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U7 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_4267, new_AGEMA_signal_4265}), .c ({new_AGEMA_signal_2121, LED_128_Instance_MCS_Instance_0_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U6 ( .a ({new_AGEMA_signal_2123, LED_128_Instance_MCS_Instance_0_n3}), .b ({new_AGEMA_signal_2122, LED_128_Instance_MCS_Instance_0_n2}), .c ({new_AGEMA_signal_2143, LED_128_Instance_mixcolumns_out[0]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U5 ( .a ({new_AGEMA_signal_2099, LED_128_Instance_subcells_out[63]}), .b ({new_AGEMA_signal_2090, LED_128_Instance_subcells_out[43]}), .c ({new_AGEMA_signal_2122, LED_128_Instance_MCS_Instance_0_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U4 ( .a ({new_AGEMA_signal_2069, LED_128_Instance_subcells_out[2]}), .b ({new_AGEMA_signal_4271, new_AGEMA_signal_4269}), .c ({new_AGEMA_signal_2123, LED_128_Instance_MCS_Instance_0_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U3 ( .a ({new_AGEMA_signal_2175, LED_128_Instance_MCS_Instance_0_n1}), .b ({new_AGEMA_signal_2066, LED_128_Instance_subcells_out[62]}), .c ({new_AGEMA_signal_2205, LED_128_Instance_mixcolumns_out[3]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U2 ( .a ({new_AGEMA_signal_2144, LED_128_Instance_MCS_Instance_0_n20}), .b ({new_AGEMA_signal_2070, LED_128_Instance_subcells_out[1]}), .c ({new_AGEMA_signal_2175, LED_128_Instance_MCS_Instance_0_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_0_U1 ( .a ({new_AGEMA_signal_2053, LED_128_Instance_subcells_out[42]}), .b ({new_AGEMA_signal_2110, LED_128_Instance_subcells_out[23]}), .c ({new_AGEMA_signal_2144, LED_128_Instance_MCS_Instance_0_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U54 ( .a ({new_AGEMA_signal_2386, LED_128_Instance_MCS_Instance_1_n38}), .b ({new_AGEMA_signal_2206, LED_128_Instance_MCS_Instance_1_n37}), .c ({new_AGEMA_signal_2429, LED_128_Instance_mixcolumns_out[55]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U53 ( .a ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2206, LED_128_Instance_MCS_Instance_1_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U52 ( .a ({new_AGEMA_signal_2290, LED_128_Instance_mixcolumns_out[38]}), .b ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}), .c ({new_AGEMA_signal_2386, LED_128_Instance_MCS_Instance_1_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U51 ( .a ({new_AGEMA_signal_2207, LED_128_Instance_MCS_Instance_1_n36}), .b ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_2290, LED_128_Instance_mixcolumns_out[38]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U50 ( .a ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2176, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_2207, LED_128_Instance_MCS_Instance_1_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U49 ( .a ({new_AGEMA_signal_2291, LED_128_Instance_MCS_Instance_1_n33}), .b ({new_AGEMA_signal_2343, LED_128_Instance_mixcolumns_out[37]}), .c ({new_AGEMA_signal_2387, LED_128_Instance_mixcolumns_out[54]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U48 ( .a ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_2291, LED_128_Instance_MCS_Instance_1_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U47 ( .a ({new_AGEMA_signal_2488, LED_128_Instance_MCS_Instance_1_n32}), .b ({new_AGEMA_signal_2295, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_2501, LED_128_Instance_mixcolumns_out[53]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U46 ( .a ({new_AGEMA_signal_2478, LED_128_Instance_MCS_Instance_1_n30}), .b ({new_AGEMA_signal_2292, LED_128_Instance_MCS_Instance_1_n29}), .c ({new_AGEMA_signal_2488, LED_128_Instance_MCS_Instance_1_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U45 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}), .c ({new_AGEMA_signal_2292, LED_128_Instance_MCS_Instance_1_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U44 ( .a ({new_AGEMA_signal_2341, LED_128_Instance_mixcolumns_out[36]}), .b ({new_AGEMA_signal_2457, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_2478, LED_128_Instance_MCS_Instance_1_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U43 ( .a ({new_AGEMA_signal_2293, LED_128_Instance_MCS_Instance_1_n27}), .b ({new_AGEMA_signal_2208, LED_128_Instance_MCS_Instance_1_n26}), .c ({new_AGEMA_signal_2341, LED_128_Instance_mixcolumns_out[36]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U42 ( .a ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .c ({new_AGEMA_signal_2208, LED_128_Instance_MCS_Instance_1_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U41 ( .a ({new_AGEMA_signal_4283, new_AGEMA_signal_4281}), .b ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_2293, LED_128_Instance_MCS_Instance_1_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U40 ( .a ({new_AGEMA_signal_2479, LED_128_Instance_MCS_Instance_1_n25}), .b ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_2489, LED_128_Instance_mixcolumns_out[52]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U39 ( .a ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .b ({new_AGEMA_signal_2457, LED_128_Instance_MCS_Instance_1_n28}), .c ({new_AGEMA_signal_2479, LED_128_Instance_MCS_Instance_1_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U38 ( .a ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2430, LED_128_Instance_mixcolumns_out[39]}), .c ({new_AGEMA_signal_2457, LED_128_Instance_MCS_Instance_1_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U37 ( .a ({new_AGEMA_signal_2388, LED_128_Instance_MCS_Instance_1_n24}), .b ({new_AGEMA_signal_2145, LED_128_Instance_MCS_Instance_1_n23}), .c ({new_AGEMA_signal_2430, LED_128_Instance_mixcolumns_out[39]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U36 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2057, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2145, LED_128_Instance_MCS_Instance_1_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U35 ( .a ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}), .b ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .c ({new_AGEMA_signal_2388, LED_128_Instance_MCS_Instance_1_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U34 ( .a ({new_AGEMA_signal_2294, LED_128_Instance_MCS_Instance_1_n22}), .b ({new_AGEMA_signal_2146, LED_128_Instance_MCS_Instance_1_n21}), .c ({new_AGEMA_signal_2342, LED_128_Instance_mixcolumns_out[22]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U33 ( .a ({new_AGEMA_signal_2130, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2146, LED_128_Instance_MCS_Instance_1_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U32 ( .a ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}), .b ({new_AGEMA_signal_4287, new_AGEMA_signal_4285}), .c ({new_AGEMA_signal_2294, LED_128_Instance_MCS_Instance_1_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U31 ( .a ({new_AGEMA_signal_2209, LED_128_Instance_MCS_Instance_1_n19}), .b ({new_AGEMA_signal_2124, LED_128_Instance_MCS_Instance_1_n18}), .c ({new_AGEMA_signal_2250, LED_128_Instance_mixcolumns_out[5]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U30 ( .a ({new_AGEMA_signal_4291, new_AGEMA_signal_4289}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2124, LED_128_Instance_MCS_Instance_1_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U29 ( .a ({new_AGEMA_signal_2149, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_2176, LED_128_Instance_MCS_Instance_1_n34}), .c ({new_AGEMA_signal_2209, LED_128_Instance_MCS_Instance_1_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U28 ( .a ({new_AGEMA_signal_2147, LED_128_Instance_MCS_Instance_1_n16}), .b ({new_AGEMA_signal_2072, LED_128_Instance_subcells_out[6]}), .c ({new_AGEMA_signal_2176, LED_128_Instance_MCS_Instance_1_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U27 ( .a ({new_AGEMA_signal_2044, LED_128_Instance_subcells_out[25]}), .b ({new_AGEMA_signal_2108, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2147, LED_128_Instance_MCS_Instance_1_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U26 ( .a ({new_AGEMA_signal_2296, LED_128_Instance_MCS_Instance_1_n15}), .b ({new_AGEMA_signal_2295, LED_128_Instance_MCS_Instance_1_n31}), .c ({new_AGEMA_signal_2343, LED_128_Instance_mixcolumns_out[37]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U25 ( .a ({new_AGEMA_signal_2252, LED_128_Instance_mixcolumns_out[20]}), .b ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}), .c ({new_AGEMA_signal_2295, LED_128_Instance_MCS_Instance_1_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U24 ( .a ({new_AGEMA_signal_2251, LED_128_Instance_MCS_Instance_1_n14}), .b ({new_AGEMA_signal_2125, LED_128_Instance_MCS_Instance_1_n13}), .c ({new_AGEMA_signal_2296, LED_128_Instance_MCS_Instance_1_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U23 ( .a ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2125, LED_128_Instance_MCS_Instance_1_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U22 ( .a ({new_AGEMA_signal_2212, LED_128_Instance_MCS_Instance_1_n12}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2251, LED_128_Instance_MCS_Instance_1_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U21 ( .a ({new_AGEMA_signal_2101, LED_128_Instance_MCS_Instance_1_n11}), .b ({new_AGEMA_signal_2210, LED_128_Instance_MCS_Instance_1_n10}), .c ({new_AGEMA_signal_2252, LED_128_Instance_mixcolumns_out[20]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U20 ( .a ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .c ({new_AGEMA_signal_2210, LED_128_Instance_MCS_Instance_1_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U19 ( .a ({new_AGEMA_signal_4291, new_AGEMA_signal_4289}), .b ({new_AGEMA_signal_2043, LED_128_Instance_subcells_out[26]}), .c ({new_AGEMA_signal_2101, LED_128_Instance_MCS_Instance_1_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U18 ( .a ({new_AGEMA_signal_2211, LED_128_Instance_MCS_Instance_1_n9}), .b ({new_AGEMA_signal_2126, LED_128_Instance_MCS_Instance_1_n8}), .c ({new_AGEMA_signal_2253, LED_128_Instance_mixcolumns_out[23]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U17 ( .a ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2126, LED_128_Instance_MCS_Instance_1_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U16 ( .a ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}), .b ({new_AGEMA_signal_2044, LED_128_Instance_subcells_out[25]}), .c ({new_AGEMA_signal_2211, LED_128_Instance_MCS_Instance_1_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U15 ( .a ({new_AGEMA_signal_2127, LED_128_Instance_MCS_Instance_1_n7}), .b ({new_AGEMA_signal_2148, LED_128_Instance_MCS_Instance_1_n6}), .c ({new_AGEMA_signal_2177, LED_128_Instance_mixcolumns_out[6]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U14 ( .a ({new_AGEMA_signal_2102, LED_128_Instance_MCS_Instance_1_n5}), .b ({new_AGEMA_signal_2108, LED_128_Instance_subcells_out[7]}), .c ({new_AGEMA_signal_2148, LED_128_Instance_MCS_Instance_1_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U13 ( .a ({new_AGEMA_signal_4295, new_AGEMA_signal_4293}), .b ({new_AGEMA_signal_2094, LED_128_Instance_subcells_out[49]}), .c ({new_AGEMA_signal_2127, LED_128_Instance_MCS_Instance_1_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U12 ( .a ({new_AGEMA_signal_2149, LED_128_Instance_MCS_Instance_1_n17}), .b ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}), .c ({new_AGEMA_signal_2297, LED_128_Instance_mixcolumns_out[21]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U11 ( .a ({new_AGEMA_signal_2128, LED_128_Instance_MCS_Instance_1_n4}), .b ({new_AGEMA_signal_2212, LED_128_Instance_MCS_Instance_1_n12}), .c ({new_AGEMA_signal_2254, LED_128_Instance_MCS_Instance_1_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U10 ( .a ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}), .b ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}), .c ({new_AGEMA_signal_2212, LED_128_Instance_MCS_Instance_1_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U9 ( .a ({new_AGEMA_signal_2082, LED_128_Instance_subcells_out[27]}), .b ({new_AGEMA_signal_2102, LED_128_Instance_MCS_Instance_1_n5}), .c ({new_AGEMA_signal_2128, LED_128_Instance_MCS_Instance_1_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U8 ( .a ({new_AGEMA_signal_2043, LED_128_Instance_subcells_out[26]}), .b ({new_AGEMA_signal_2057, LED_128_Instance_subcells_out[45]}), .c ({new_AGEMA_signal_2102, LED_128_Instance_MCS_Instance_1_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U7 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_4283, new_AGEMA_signal_4281}), .c ({new_AGEMA_signal_2149, LED_128_Instance_MCS_Instance_1_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U6 ( .a ({new_AGEMA_signal_2129, LED_128_Instance_MCS_Instance_1_n3}), .b ({new_AGEMA_signal_2150, LED_128_Instance_MCS_Instance_1_n2}), .c ({new_AGEMA_signal_2178, LED_128_Instance_mixcolumns_out[4]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U5 ( .a ({new_AGEMA_signal_2113, LED_128_Instance_subcells_out[51]}), .b ({new_AGEMA_signal_2091, LED_128_Instance_subcells_out[47]}), .c ({new_AGEMA_signal_2150, LED_128_Instance_MCS_Instance_1_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U4 ( .a ({new_AGEMA_signal_2072, LED_128_Instance_subcells_out[6]}), .b ({new_AGEMA_signal_4287, new_AGEMA_signal_4285}), .c ({new_AGEMA_signal_2129, LED_128_Instance_MCS_Instance_1_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U3 ( .a ({new_AGEMA_signal_2151, LED_128_Instance_MCS_Instance_1_n1}), .b ({new_AGEMA_signal_2093, LED_128_Instance_subcells_out[50]}), .c ({new_AGEMA_signal_2179, LED_128_Instance_mixcolumns_out[7]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U2 ( .a ({new_AGEMA_signal_2130, LED_128_Instance_MCS_Instance_1_n20}), .b ({new_AGEMA_signal_2073, LED_128_Instance_subcells_out[5]}), .c ({new_AGEMA_signal_2151, LED_128_Instance_MCS_Instance_1_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_1_U1 ( .a ({new_AGEMA_signal_2056, LED_128_Instance_subcells_out[46]}), .b ({new_AGEMA_signal_2082, LED_128_Instance_subcells_out[27]}), .c ({new_AGEMA_signal_2130, LED_128_Instance_MCS_Instance_1_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U54 ( .a ({new_AGEMA_signal_2344, LED_128_Instance_MCS_Instance_2_n38}), .b ({new_AGEMA_signal_2213, LED_128_Instance_MCS_Instance_2_n37}), .c ({new_AGEMA_signal_2389, LED_128_Instance_mixcolumns_out[59]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U53 ( .a ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2213, LED_128_Instance_MCS_Instance_2_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U52 ( .a ({new_AGEMA_signal_2298, LED_128_Instance_mixcolumns_out[42]}), .b ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}), .c ({new_AGEMA_signal_2344, LED_128_Instance_MCS_Instance_2_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U51 ( .a ({new_AGEMA_signal_2180, LED_128_Instance_MCS_Instance_2_n36}), .b ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_2298, LED_128_Instance_mixcolumns_out[42]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U50 ( .a ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2155, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_2180, LED_128_Instance_MCS_Instance_2_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U49 ( .a ({new_AGEMA_signal_2299, LED_128_Instance_MCS_Instance_2_n33}), .b ({new_AGEMA_signal_2347, LED_128_Instance_mixcolumns_out[41]}), .c ({new_AGEMA_signal_2390, LED_128_Instance_mixcolumns_out[58]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U48 ( .a ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_2299, LED_128_Instance_MCS_Instance_2_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U47 ( .a ({new_AGEMA_signal_2480, LED_128_Instance_MCS_Instance_2_n32}), .b ({new_AGEMA_signal_2302, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_2490, LED_128_Instance_mixcolumns_out[57]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U46 ( .a ({new_AGEMA_signal_2458, LED_128_Instance_MCS_Instance_2_n30}), .b ({new_AGEMA_signal_2255, LED_128_Instance_MCS_Instance_2_n29}), .c ({new_AGEMA_signal_2480, LED_128_Instance_MCS_Instance_2_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U45 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}), .c ({new_AGEMA_signal_2255, LED_128_Instance_MCS_Instance_2_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U44 ( .a ({new_AGEMA_signal_2345, LED_128_Instance_mixcolumns_out[40]}), .b ({new_AGEMA_signal_2431, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_2458, LED_128_Instance_MCS_Instance_2_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U43 ( .a ({new_AGEMA_signal_2300, LED_128_Instance_MCS_Instance_2_n27}), .b ({new_AGEMA_signal_2214, LED_128_Instance_MCS_Instance_2_n26}), .c ({new_AGEMA_signal_2345, LED_128_Instance_mixcolumns_out[40]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U42 ( .a ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .c ({new_AGEMA_signal_2214, LED_128_Instance_MCS_Instance_2_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U41 ( .a ({new_AGEMA_signal_4299, new_AGEMA_signal_4297}), .b ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_2300, LED_128_Instance_MCS_Instance_2_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U40 ( .a ({new_AGEMA_signal_2459, LED_128_Instance_MCS_Instance_2_n25}), .b ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_2481, LED_128_Instance_mixcolumns_out[56]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U39 ( .a ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .b ({new_AGEMA_signal_2431, LED_128_Instance_MCS_Instance_2_n28}), .c ({new_AGEMA_signal_2459, LED_128_Instance_MCS_Instance_2_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U38 ( .a ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2391, LED_128_Instance_mixcolumns_out[43]}), .c ({new_AGEMA_signal_2431, LED_128_Instance_MCS_Instance_2_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U37 ( .a ({new_AGEMA_signal_2346, LED_128_Instance_MCS_Instance_2_n24}), .b ({new_AGEMA_signal_2152, LED_128_Instance_MCS_Instance_2_n23}), .c ({new_AGEMA_signal_2391, LED_128_Instance_mixcolumns_out[43]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U36 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2086, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2152, LED_128_Instance_MCS_Instance_2_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U35 ( .a ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}), .b ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .c ({new_AGEMA_signal_2346, LED_128_Instance_MCS_Instance_2_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U34 ( .a ({new_AGEMA_signal_2256, LED_128_Instance_MCS_Instance_2_n22}), .b ({new_AGEMA_signal_2153, LED_128_Instance_MCS_Instance_2_n21}), .c ({new_AGEMA_signal_2301, LED_128_Instance_mixcolumns_out[26]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U33 ( .a ({new_AGEMA_signal_2134, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2153, LED_128_Instance_MCS_Instance_2_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U32 ( .a ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}), .b ({new_AGEMA_signal_4303, new_AGEMA_signal_4301}), .c ({new_AGEMA_signal_2256, LED_128_Instance_MCS_Instance_2_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U31 ( .a ({new_AGEMA_signal_2181, LED_128_Instance_MCS_Instance_2_n19}), .b ({new_AGEMA_signal_2154, LED_128_Instance_MCS_Instance_2_n18}), .c ({new_AGEMA_signal_2215, LED_128_Instance_mixcolumns_out[9]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U30 ( .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4305}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2154, LED_128_Instance_MCS_Instance_2_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U29 ( .a ({new_AGEMA_signal_2160, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_2155, LED_128_Instance_MCS_Instance_2_n34}), .c ({new_AGEMA_signal_2181, LED_128_Instance_MCS_Instance_2_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U28 ( .a ({new_AGEMA_signal_2131, LED_128_Instance_MCS_Instance_2_n16}), .b ({new_AGEMA_signal_2033, LED_128_Instance_subcells_out[10]}), .c ({new_AGEMA_signal_2155, LED_128_Instance_MCS_Instance_2_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U27 ( .a ({new_AGEMA_signal_2047, LED_128_Instance_subcells_out[29]}), .b ({new_AGEMA_signal_2074, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2131, LED_128_Instance_MCS_Instance_2_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U26 ( .a ({new_AGEMA_signal_2303, LED_128_Instance_MCS_Instance_2_n15}), .b ({new_AGEMA_signal_2302, LED_128_Instance_MCS_Instance_2_n31}), .c ({new_AGEMA_signal_2347, LED_128_Instance_mixcolumns_out[41]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U25 ( .a ({new_AGEMA_signal_2258, LED_128_Instance_mixcolumns_out[24]}), .b ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}), .c ({new_AGEMA_signal_2302, LED_128_Instance_MCS_Instance_2_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U24 ( .a ({new_AGEMA_signal_2257, LED_128_Instance_MCS_Instance_2_n14}), .b ({new_AGEMA_signal_2156, LED_128_Instance_MCS_Instance_2_n13}), .c ({new_AGEMA_signal_2303, LED_128_Instance_MCS_Instance_2_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U23 ( .a ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2156, LED_128_Instance_MCS_Instance_2_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U22 ( .a ({new_AGEMA_signal_2218, LED_128_Instance_MCS_Instance_2_n12}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2257, LED_128_Instance_MCS_Instance_2_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U21 ( .a ({new_AGEMA_signal_2103, LED_128_Instance_MCS_Instance_2_n11}), .b ({new_AGEMA_signal_2216, LED_128_Instance_MCS_Instance_2_n10}), .c ({new_AGEMA_signal_2258, LED_128_Instance_mixcolumns_out[24]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U20 ( .a ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .c ({new_AGEMA_signal_2216, LED_128_Instance_MCS_Instance_2_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U19 ( .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4305}), .b ({new_AGEMA_signal_2046, LED_128_Instance_subcells_out[30]}), .c ({new_AGEMA_signal_2103, LED_128_Instance_MCS_Instance_2_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U18 ( .a ({new_AGEMA_signal_2217, LED_128_Instance_MCS_Instance_2_n9}), .b ({new_AGEMA_signal_2157, LED_128_Instance_MCS_Instance_2_n8}), .c ({new_AGEMA_signal_2259, LED_128_Instance_mixcolumns_out[27]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U17 ( .a ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2157, LED_128_Instance_MCS_Instance_2_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U16 ( .a ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}), .b ({new_AGEMA_signal_2047, LED_128_Instance_subcells_out[29]}), .c ({new_AGEMA_signal_2217, LED_128_Instance_MCS_Instance_2_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U15 ( .a ({new_AGEMA_signal_2132, LED_128_Instance_MCS_Instance_2_n7}), .b ({new_AGEMA_signal_2158, LED_128_Instance_MCS_Instance_2_n6}), .c ({new_AGEMA_signal_2182, LED_128_Instance_mixcolumns_out[10]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U14 ( .a ({new_AGEMA_signal_2133, LED_128_Instance_MCS_Instance_2_n5}), .b ({new_AGEMA_signal_2074, LED_128_Instance_subcells_out[11]}), .c ({new_AGEMA_signal_2158, LED_128_Instance_MCS_Instance_2_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U13 ( .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4309}), .b ({new_AGEMA_signal_2097, LED_128_Instance_subcells_out[53]}), .c ({new_AGEMA_signal_2132, LED_128_Instance_MCS_Instance_2_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U12 ( .a ({new_AGEMA_signal_2160, LED_128_Instance_MCS_Instance_2_n17}), .b ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}), .c ({new_AGEMA_signal_2304, LED_128_Instance_mixcolumns_out[25]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U11 ( .a ({new_AGEMA_signal_2159, LED_128_Instance_MCS_Instance_2_n4}), .b ({new_AGEMA_signal_2218, LED_128_Instance_MCS_Instance_2_n12}), .c ({new_AGEMA_signal_2260, LED_128_Instance_MCS_Instance_2_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U10 ( .a ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}), .b ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}), .c ({new_AGEMA_signal_2218, LED_128_Instance_MCS_Instance_2_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U9 ( .a ({new_AGEMA_signal_2083, LED_128_Instance_subcells_out[31]}), .b ({new_AGEMA_signal_2133, LED_128_Instance_MCS_Instance_2_n5}), .c ({new_AGEMA_signal_2159, LED_128_Instance_MCS_Instance_2_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U8 ( .a ({new_AGEMA_signal_2046, LED_128_Instance_subcells_out[30]}), .b ({new_AGEMA_signal_2086, LED_128_Instance_subcells_out[33]}), .c ({new_AGEMA_signal_2133, LED_128_Instance_MCS_Instance_2_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U7 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_4299, new_AGEMA_signal_4297}), .c ({new_AGEMA_signal_2160, LED_128_Instance_MCS_Instance_2_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U6 ( .a ({new_AGEMA_signal_2104, LED_128_Instance_MCS_Instance_2_n3}), .b ({new_AGEMA_signal_2161, LED_128_Instance_MCS_Instance_2_n2}), .c ({new_AGEMA_signal_2183, LED_128_Instance_mixcolumns_out[8]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U5 ( .a ({new_AGEMA_signal_2114, LED_128_Instance_subcells_out[55]}), .b ({new_AGEMA_signal_2111, LED_128_Instance_subcells_out[35]}), .c ({new_AGEMA_signal_2161, LED_128_Instance_MCS_Instance_2_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U4 ( .a ({new_AGEMA_signal_2033, LED_128_Instance_subcells_out[10]}), .b ({new_AGEMA_signal_4303, new_AGEMA_signal_4301}), .c ({new_AGEMA_signal_2104, LED_128_Instance_MCS_Instance_2_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U3 ( .a ({new_AGEMA_signal_2162, LED_128_Instance_MCS_Instance_2_n1}), .b ({new_AGEMA_signal_2096, LED_128_Instance_subcells_out[54]}), .c ({new_AGEMA_signal_2184, LED_128_Instance_mixcolumns_out[11]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U2 ( .a ({new_AGEMA_signal_2134, LED_128_Instance_MCS_Instance_2_n20}), .b ({new_AGEMA_signal_2034, LED_128_Instance_subcells_out[9]}), .c ({new_AGEMA_signal_2162, LED_128_Instance_MCS_Instance_2_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_2_U1 ( .a ({new_AGEMA_signal_2085, LED_128_Instance_subcells_out[34]}), .b ({new_AGEMA_signal_2083, LED_128_Instance_subcells_out[31]}), .c ({new_AGEMA_signal_2134, LED_128_Instance_MCS_Instance_2_n20}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U54 ( .a ({new_AGEMA_signal_2392, LED_128_Instance_MCS_Instance_3_n38}), .b ({new_AGEMA_signal_2261, LED_128_Instance_MCS_Instance_3_n37}), .c ({new_AGEMA_signal_2432, LED_128_Instance_mixcolumns_out[63]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U53 ( .a ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2261, LED_128_Instance_MCS_Instance_3_n37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U52 ( .a ({new_AGEMA_signal_2348, LED_128_Instance_mixcolumns_out[46]}), .b ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}), .c ({new_AGEMA_signal_2392, LED_128_Instance_MCS_Instance_3_n38}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U51 ( .a ({new_AGEMA_signal_2185, LED_128_Instance_MCS_Instance_3_n36}), .b ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_2348, LED_128_Instance_mixcolumns_out[46]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U50 ( .a ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2164, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_2185, LED_128_Instance_MCS_Instance_3_n36}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U49 ( .a ({new_AGEMA_signal_2349, LED_128_Instance_MCS_Instance_3_n33}), .b ({new_AGEMA_signal_2394, LED_128_Instance_mixcolumns_out[45]}), .c ({new_AGEMA_signal_2433, LED_128_Instance_mixcolumns_out[62]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U48 ( .a ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_2349, LED_128_Instance_MCS_Instance_3_n33}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U47 ( .a ({new_AGEMA_signal_2482, LED_128_Instance_MCS_Instance_3_n32}), .b ({new_AGEMA_signal_2352, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_2491, LED_128_Instance_mixcolumns_out[61]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U46 ( .a ({new_AGEMA_signal_2460, LED_128_Instance_MCS_Instance_3_n30}), .b ({new_AGEMA_signal_2262, LED_128_Instance_MCS_Instance_3_n29}), .c ({new_AGEMA_signal_2482, LED_128_Instance_MCS_Instance_3_n32}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U45 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}), .c ({new_AGEMA_signal_2262, LED_128_Instance_MCS_Instance_3_n29}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U44 ( .a ({new_AGEMA_signal_2350, LED_128_Instance_mixcolumns_out[44]}), .b ({new_AGEMA_signal_2434, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_2460, LED_128_Instance_MCS_Instance_3_n30}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U43 ( .a ({new_AGEMA_signal_2305, LED_128_Instance_MCS_Instance_3_n27}), .b ({new_AGEMA_signal_2263, LED_128_Instance_MCS_Instance_3_n26}), .c ({new_AGEMA_signal_2350, LED_128_Instance_mixcolumns_out[44]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U42 ( .a ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .c ({new_AGEMA_signal_2263, LED_128_Instance_MCS_Instance_3_n26}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U41 ( .a ({new_AGEMA_signal_4315, new_AGEMA_signal_4313}), .b ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_2305, LED_128_Instance_MCS_Instance_3_n27}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U40 ( .a ({new_AGEMA_signal_2461, LED_128_Instance_MCS_Instance_3_n25}), .b ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_2483, LED_128_Instance_mixcolumns_out[60]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U39 ( .a ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .b ({new_AGEMA_signal_2434, LED_128_Instance_MCS_Instance_3_n28}), .c ({new_AGEMA_signal_2461, LED_128_Instance_MCS_Instance_3_n25}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U38 ( .a ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2393, LED_128_Instance_mixcolumns_out[47]}), .c ({new_AGEMA_signal_2434, LED_128_Instance_MCS_Instance_3_n28}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U37 ( .a ({new_AGEMA_signal_2351, LED_128_Instance_MCS_Instance_3_n24}), .b ({new_AGEMA_signal_2135, LED_128_Instance_MCS_Instance_3_n23}), .c ({new_AGEMA_signal_2393, LED_128_Instance_mixcolumns_out[47]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U36 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2089, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2135, LED_128_Instance_MCS_Instance_3_n23}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U35 ( .a ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}), .b ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .c ({new_AGEMA_signal_2351, LED_128_Instance_MCS_Instance_3_n24}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U34 ( .a ({new_AGEMA_signal_2264, LED_128_Instance_MCS_Instance_3_n22}), .b ({new_AGEMA_signal_2186, LED_128_Instance_MCS_Instance_3_n21}), .c ({new_AGEMA_signal_2306, LED_128_Instance_mixcolumns_out[30]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U33 ( .a ({new_AGEMA_signal_2170, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2186, LED_128_Instance_MCS_Instance_3_n21}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U32 ( .a ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}), .b ({new_AGEMA_signal_4319, new_AGEMA_signal_4317}), .c ({new_AGEMA_signal_2264, LED_128_Instance_MCS_Instance_3_n22}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U31 ( .a ({new_AGEMA_signal_2187, LED_128_Instance_MCS_Instance_3_n19}), .b ({new_AGEMA_signal_2163, LED_128_Instance_MCS_Instance_3_n18}), .c ({new_AGEMA_signal_2219, LED_128_Instance_mixcolumns_out[13]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U30 ( .a ({new_AGEMA_signal_4323, new_AGEMA_signal_4321}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2163, LED_128_Instance_MCS_Instance_3_n18}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U29 ( .a ({new_AGEMA_signal_2139, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_2164, LED_128_Instance_MCS_Instance_3_n34}), .c ({new_AGEMA_signal_2187, LED_128_Instance_MCS_Instance_3_n19}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U28 ( .a ({new_AGEMA_signal_2136, LED_128_Instance_MCS_Instance_3_n16}), .b ({new_AGEMA_signal_2036, LED_128_Instance_subcells_out[14]}), .c ({new_AGEMA_signal_2164, LED_128_Instance_MCS_Instance_3_n34}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U27 ( .a ({new_AGEMA_signal_2078, LED_128_Instance_subcells_out[17]}), .b ({new_AGEMA_signal_2075, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_2136, LED_128_Instance_MCS_Instance_3_n16}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U26 ( .a ({new_AGEMA_signal_2353, LED_128_Instance_MCS_Instance_3_n15}), .b ({new_AGEMA_signal_2352, LED_128_Instance_MCS_Instance_3_n31}), .c ({new_AGEMA_signal_2394, LED_128_Instance_mixcolumns_out[45]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U25 ( .a ({new_AGEMA_signal_2308, LED_128_Instance_mixcolumns_out[28]}), .b ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}), .c ({new_AGEMA_signal_2352, LED_128_Instance_MCS_Instance_3_n31}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U24 ( .a ({new_AGEMA_signal_2307, LED_128_Instance_MCS_Instance_3_n14}), .b ({new_AGEMA_signal_2165, LED_128_Instance_MCS_Instance_3_n13}), .c ({new_AGEMA_signal_2353, LED_128_Instance_MCS_Instance_3_n15}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U23 ( .a ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2165, LED_128_Instance_MCS_Instance_3_n13}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U22 ( .a ({new_AGEMA_signal_2267, LED_128_Instance_MCS_Instance_3_n12}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2307, LED_128_Instance_MCS_Instance_3_n14}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U21 ( .a ({new_AGEMA_signal_2137, LED_128_Instance_MCS_Instance_3_n11}), .b ({new_AGEMA_signal_2265, LED_128_Instance_MCS_Instance_3_n10}), .c ({new_AGEMA_signal_2308, LED_128_Instance_mixcolumns_out[28]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U20 ( .a ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .c ({new_AGEMA_signal_2265, LED_128_Instance_MCS_Instance_3_n10}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U19 ( .a ({new_AGEMA_signal_4323, new_AGEMA_signal_4321}), .b ({new_AGEMA_signal_2077, LED_128_Instance_subcells_out[18]}), .c ({new_AGEMA_signal_2137, LED_128_Instance_MCS_Instance_3_n11}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U18 ( .a ({new_AGEMA_signal_2220, LED_128_Instance_MCS_Instance_3_n9}), .b ({new_AGEMA_signal_2166, LED_128_Instance_MCS_Instance_3_n8}), .c ({new_AGEMA_signal_2266, LED_128_Instance_mixcolumns_out[31]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U17 ( .a ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2166, LED_128_Instance_MCS_Instance_3_n8}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U16 ( .a ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}), .b ({new_AGEMA_signal_2078, LED_128_Instance_subcells_out[17]}), .c ({new_AGEMA_signal_2220, LED_128_Instance_MCS_Instance_3_n9}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U15 ( .a ({new_AGEMA_signal_2105, LED_128_Instance_MCS_Instance_3_n7}), .b ({new_AGEMA_signal_2167, LED_128_Instance_MCS_Instance_3_n6}), .c ({new_AGEMA_signal_2188, LED_128_Instance_mixcolumns_out[14]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U14 ( .a ({new_AGEMA_signal_2138, LED_128_Instance_MCS_Instance_3_n5}), .b ({new_AGEMA_signal_2075, LED_128_Instance_subcells_out[15]}), .c ({new_AGEMA_signal_2167, LED_128_Instance_MCS_Instance_3_n6}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U13 ( .a ({new_AGEMA_signal_4327, new_AGEMA_signal_4325}), .b ({new_AGEMA_signal_2064, LED_128_Instance_subcells_out[57]}), .c ({new_AGEMA_signal_2105, LED_128_Instance_MCS_Instance_3_n7}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U12 ( .a ({new_AGEMA_signal_2139, LED_128_Instance_MCS_Instance_3_n17}), .b ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}), .c ({new_AGEMA_signal_2354, LED_128_Instance_mixcolumns_out[29]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U11 ( .a ({new_AGEMA_signal_2168, LED_128_Instance_MCS_Instance_3_n4}), .b ({new_AGEMA_signal_2267, LED_128_Instance_MCS_Instance_3_n12}), .c ({new_AGEMA_signal_2309, LED_128_Instance_MCS_Instance_3_n35}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U10 ( .a ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}), .b ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}), .c ({new_AGEMA_signal_2267, LED_128_Instance_MCS_Instance_3_n12}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U9 ( .a ({new_AGEMA_signal_2109, LED_128_Instance_subcells_out[19]}), .b ({new_AGEMA_signal_2138, LED_128_Instance_MCS_Instance_3_n5}), .c ({new_AGEMA_signal_2168, LED_128_Instance_MCS_Instance_3_n4}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U8 ( .a ({new_AGEMA_signal_2077, LED_128_Instance_subcells_out[18]}), .b ({new_AGEMA_signal_2089, LED_128_Instance_subcells_out[37]}), .c ({new_AGEMA_signal_2138, LED_128_Instance_MCS_Instance_3_n5}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U7 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_4315, new_AGEMA_signal_4313}), .c ({new_AGEMA_signal_2139, LED_128_Instance_MCS_Instance_3_n17}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U6 ( .a ({new_AGEMA_signal_2106, LED_128_Instance_MCS_Instance_3_n3}), .b ({new_AGEMA_signal_2169, LED_128_Instance_MCS_Instance_3_n2}), .c ({new_AGEMA_signal_2189, LED_128_Instance_mixcolumns_out[12]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U5 ( .a ({new_AGEMA_signal_2098, LED_128_Instance_subcells_out[59]}), .b ({new_AGEMA_signal_2112, LED_128_Instance_subcells_out[39]}), .c ({new_AGEMA_signal_2169, LED_128_Instance_MCS_Instance_3_n2}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U4 ( .a ({new_AGEMA_signal_2036, LED_128_Instance_subcells_out[14]}), .b ({new_AGEMA_signal_4319, new_AGEMA_signal_4317}), .c ({new_AGEMA_signal_2106, LED_128_Instance_MCS_Instance_3_n3}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U3 ( .a ({new_AGEMA_signal_2190, LED_128_Instance_MCS_Instance_3_n1}), .b ({new_AGEMA_signal_2063, LED_128_Instance_subcells_out[58]}), .c ({new_AGEMA_signal_2221, LED_128_Instance_mixcolumns_out[15]}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U2 ( .a ({new_AGEMA_signal_2170, LED_128_Instance_MCS_Instance_3_n20}), .b ({new_AGEMA_signal_2037, LED_128_Instance_subcells_out[13]}), .c ({new_AGEMA_signal_2190, LED_128_Instance_MCS_Instance_3_n1}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) LED_128_Instance_MCS_Instance_3_U1 ( .a ({new_AGEMA_signal_2088, LED_128_Instance_subcells_out[38]}), .b ({new_AGEMA_signal_2109, LED_128_Instance_subcells_out[19]}), .c ({new_AGEMA_signal_2170, LED_128_Instance_MCS_Instance_3_n20}) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (CLK), .D (new_AGEMA_signal_2774), .Q (new_AGEMA_signal_2775) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (CLK), .D (new_AGEMA_signal_2778), .Q (new_AGEMA_signal_2779) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (CLK), .D (new_AGEMA_signal_2782), .Q (new_AGEMA_signal_2783) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (CLK), .D (new_AGEMA_signal_2786), .Q (new_AGEMA_signal_2787) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (CLK), .D (new_AGEMA_signal_2790), .Q (new_AGEMA_signal_2791) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (CLK), .D (new_AGEMA_signal_2794), .Q (new_AGEMA_signal_2795) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (CLK), .D (new_AGEMA_signal_2798), .Q (new_AGEMA_signal_2799) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (CLK), .D (new_AGEMA_signal_2802), .Q (new_AGEMA_signal_2803) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (CLK), .D (new_AGEMA_signal_2806), .Q (new_AGEMA_signal_2807) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (CLK), .D (new_AGEMA_signal_2810), .Q (new_AGEMA_signal_2811) ) ;
    buf_clk new_AGEMA_reg_buffer_1363 ( .C (CLK), .D (new_AGEMA_signal_2814), .Q (new_AGEMA_signal_2815) ) ;
    buf_clk new_AGEMA_reg_buffer_1367 ( .C (CLK), .D (new_AGEMA_signal_2818), .Q (new_AGEMA_signal_2819) ) ;
    buf_clk new_AGEMA_reg_buffer_1371 ( .C (CLK), .D (new_AGEMA_signal_2822), .Q (new_AGEMA_signal_2823) ) ;
    buf_clk new_AGEMA_reg_buffer_1375 ( .C (CLK), .D (new_AGEMA_signal_2826), .Q (new_AGEMA_signal_2827) ) ;
    buf_clk new_AGEMA_reg_buffer_1379 ( .C (CLK), .D (new_AGEMA_signal_2830), .Q (new_AGEMA_signal_2831) ) ;
    buf_clk new_AGEMA_reg_buffer_1383 ( .C (CLK), .D (new_AGEMA_signal_2834), .Q (new_AGEMA_signal_2835) ) ;
    buf_clk new_AGEMA_reg_buffer_1387 ( .C (CLK), .D (new_AGEMA_signal_2838), .Q (new_AGEMA_signal_2839) ) ;
    buf_clk new_AGEMA_reg_buffer_1391 ( .C (CLK), .D (new_AGEMA_signal_2842), .Q (new_AGEMA_signal_2843) ) ;
    buf_clk new_AGEMA_reg_buffer_1395 ( .C (CLK), .D (new_AGEMA_signal_2846), .Q (new_AGEMA_signal_2847) ) ;
    buf_clk new_AGEMA_reg_buffer_1399 ( .C (CLK), .D (new_AGEMA_signal_2850), .Q (new_AGEMA_signal_2851) ) ;
    buf_clk new_AGEMA_reg_buffer_1403 ( .C (CLK), .D (new_AGEMA_signal_2854), .Q (new_AGEMA_signal_2855) ) ;
    buf_clk new_AGEMA_reg_buffer_1407 ( .C (CLK), .D (new_AGEMA_signal_2858), .Q (new_AGEMA_signal_2859) ) ;
    buf_clk new_AGEMA_reg_buffer_1411 ( .C (CLK), .D (new_AGEMA_signal_2862), .Q (new_AGEMA_signal_2863) ) ;
    buf_clk new_AGEMA_reg_buffer_1415 ( .C (CLK), .D (new_AGEMA_signal_2866), .Q (new_AGEMA_signal_2867) ) ;
    buf_clk new_AGEMA_reg_buffer_1419 ( .C (CLK), .D (new_AGEMA_signal_2870), .Q (new_AGEMA_signal_2871) ) ;
    buf_clk new_AGEMA_reg_buffer_1423 ( .C (CLK), .D (new_AGEMA_signal_2874), .Q (new_AGEMA_signal_2875) ) ;
    buf_clk new_AGEMA_reg_buffer_1427 ( .C (CLK), .D (new_AGEMA_signal_2878), .Q (new_AGEMA_signal_2879) ) ;
    buf_clk new_AGEMA_reg_buffer_1431 ( .C (CLK), .D (new_AGEMA_signal_2882), .Q (new_AGEMA_signal_2883) ) ;
    buf_clk new_AGEMA_reg_buffer_1435 ( .C (CLK), .D (new_AGEMA_signal_2886), .Q (new_AGEMA_signal_2887) ) ;
    buf_clk new_AGEMA_reg_buffer_1439 ( .C (CLK), .D (new_AGEMA_signal_2890), .Q (new_AGEMA_signal_2891) ) ;
    buf_clk new_AGEMA_reg_buffer_1443 ( .C (CLK), .D (new_AGEMA_signal_2894), .Q (new_AGEMA_signal_2895) ) ;
    buf_clk new_AGEMA_reg_buffer_1447 ( .C (CLK), .D (new_AGEMA_signal_2898), .Q (new_AGEMA_signal_2899) ) ;
    buf_clk new_AGEMA_reg_buffer_1451 ( .C (CLK), .D (new_AGEMA_signal_2902), .Q (new_AGEMA_signal_2903) ) ;
    buf_clk new_AGEMA_reg_buffer_1455 ( .C (CLK), .D (new_AGEMA_signal_2906), .Q (new_AGEMA_signal_2907) ) ;
    buf_clk new_AGEMA_reg_buffer_1459 ( .C (CLK), .D (new_AGEMA_signal_2910), .Q (new_AGEMA_signal_2911) ) ;
    buf_clk new_AGEMA_reg_buffer_1463 ( .C (CLK), .D (new_AGEMA_signal_2914), .Q (new_AGEMA_signal_2915) ) ;
    buf_clk new_AGEMA_reg_buffer_1467 ( .C (CLK), .D (new_AGEMA_signal_2918), .Q (new_AGEMA_signal_2919) ) ;
    buf_clk new_AGEMA_reg_buffer_1471 ( .C (CLK), .D (new_AGEMA_signal_2922), .Q (new_AGEMA_signal_2923) ) ;
    buf_clk new_AGEMA_reg_buffer_1475 ( .C (CLK), .D (new_AGEMA_signal_2926), .Q (new_AGEMA_signal_2927) ) ;
    buf_clk new_AGEMA_reg_buffer_1479 ( .C (CLK), .D (new_AGEMA_signal_2930), .Q (new_AGEMA_signal_2931) ) ;
    buf_clk new_AGEMA_reg_buffer_1483 ( .C (CLK), .D (new_AGEMA_signal_2934), .Q (new_AGEMA_signal_2935) ) ;
    buf_clk new_AGEMA_reg_buffer_1487 ( .C (CLK), .D (new_AGEMA_signal_2938), .Q (new_AGEMA_signal_2939) ) ;
    buf_clk new_AGEMA_reg_buffer_1491 ( .C (CLK), .D (new_AGEMA_signal_2942), .Q (new_AGEMA_signal_2943) ) ;
    buf_clk new_AGEMA_reg_buffer_1495 ( .C (CLK), .D (new_AGEMA_signal_2946), .Q (new_AGEMA_signal_2947) ) ;
    buf_clk new_AGEMA_reg_buffer_1499 ( .C (CLK), .D (new_AGEMA_signal_2950), .Q (new_AGEMA_signal_2951) ) ;
    buf_clk new_AGEMA_reg_buffer_1503 ( .C (CLK), .D (new_AGEMA_signal_2954), .Q (new_AGEMA_signal_2955) ) ;
    buf_clk new_AGEMA_reg_buffer_1507 ( .C (CLK), .D (new_AGEMA_signal_2958), .Q (new_AGEMA_signal_2959) ) ;
    buf_clk new_AGEMA_reg_buffer_1511 ( .C (CLK), .D (new_AGEMA_signal_2962), .Q (new_AGEMA_signal_2963) ) ;
    buf_clk new_AGEMA_reg_buffer_1515 ( .C (CLK), .D (new_AGEMA_signal_2966), .Q (new_AGEMA_signal_2967) ) ;
    buf_clk new_AGEMA_reg_buffer_1519 ( .C (CLK), .D (new_AGEMA_signal_2970), .Q (new_AGEMA_signal_2971) ) ;
    buf_clk new_AGEMA_reg_buffer_1523 ( .C (CLK), .D (new_AGEMA_signal_2974), .Q (new_AGEMA_signal_2975) ) ;
    buf_clk new_AGEMA_reg_buffer_1527 ( .C (CLK), .D (new_AGEMA_signal_2978), .Q (new_AGEMA_signal_2979) ) ;
    buf_clk new_AGEMA_reg_buffer_1531 ( .C (CLK), .D (new_AGEMA_signal_2982), .Q (new_AGEMA_signal_2983) ) ;
    buf_clk new_AGEMA_reg_buffer_1535 ( .C (CLK), .D (new_AGEMA_signal_2986), .Q (new_AGEMA_signal_2987) ) ;
    buf_clk new_AGEMA_reg_buffer_1539 ( .C (CLK), .D (new_AGEMA_signal_2990), .Q (new_AGEMA_signal_2991) ) ;
    buf_clk new_AGEMA_reg_buffer_1543 ( .C (CLK), .D (new_AGEMA_signal_2994), .Q (new_AGEMA_signal_2995) ) ;
    buf_clk new_AGEMA_reg_buffer_1547 ( .C (CLK), .D (new_AGEMA_signal_2998), .Q (new_AGEMA_signal_2999) ) ;
    buf_clk new_AGEMA_reg_buffer_1551 ( .C (CLK), .D (new_AGEMA_signal_3002), .Q (new_AGEMA_signal_3003) ) ;
    buf_clk new_AGEMA_reg_buffer_1555 ( .C (CLK), .D (new_AGEMA_signal_3006), .Q (new_AGEMA_signal_3007) ) ;
    buf_clk new_AGEMA_reg_buffer_1559 ( .C (CLK), .D (new_AGEMA_signal_3010), .Q (new_AGEMA_signal_3011) ) ;
    buf_clk new_AGEMA_reg_buffer_1563 ( .C (CLK), .D (new_AGEMA_signal_3014), .Q (new_AGEMA_signal_3015) ) ;
    buf_clk new_AGEMA_reg_buffer_1567 ( .C (CLK), .D (new_AGEMA_signal_3018), .Q (new_AGEMA_signal_3019) ) ;
    buf_clk new_AGEMA_reg_buffer_1571 ( .C (CLK), .D (new_AGEMA_signal_3022), .Q (new_AGEMA_signal_3023) ) ;
    buf_clk new_AGEMA_reg_buffer_1575 ( .C (CLK), .D (new_AGEMA_signal_3026), .Q (new_AGEMA_signal_3027) ) ;
    buf_clk new_AGEMA_reg_buffer_1579 ( .C (CLK), .D (new_AGEMA_signal_3030), .Q (new_AGEMA_signal_3031) ) ;
    buf_clk new_AGEMA_reg_buffer_1583 ( .C (CLK), .D (new_AGEMA_signal_3034), .Q (new_AGEMA_signal_3035) ) ;
    buf_clk new_AGEMA_reg_buffer_1587 ( .C (CLK), .D (new_AGEMA_signal_3038), .Q (new_AGEMA_signal_3039) ) ;
    buf_clk new_AGEMA_reg_buffer_1591 ( .C (CLK), .D (new_AGEMA_signal_3042), .Q (new_AGEMA_signal_3043) ) ;
    buf_clk new_AGEMA_reg_buffer_1595 ( .C (CLK), .D (new_AGEMA_signal_3046), .Q (new_AGEMA_signal_3047) ) ;
    buf_clk new_AGEMA_reg_buffer_1599 ( .C (CLK), .D (new_AGEMA_signal_3050), .Q (new_AGEMA_signal_3051) ) ;
    buf_clk new_AGEMA_reg_buffer_1603 ( .C (CLK), .D (new_AGEMA_signal_3054), .Q (new_AGEMA_signal_3055) ) ;
    buf_clk new_AGEMA_reg_buffer_1607 ( .C (CLK), .D (new_AGEMA_signal_3058), .Q (new_AGEMA_signal_3059) ) ;
    buf_clk new_AGEMA_reg_buffer_1611 ( .C (CLK), .D (new_AGEMA_signal_3062), .Q (new_AGEMA_signal_3063) ) ;
    buf_clk new_AGEMA_reg_buffer_1615 ( .C (CLK), .D (new_AGEMA_signal_3066), .Q (new_AGEMA_signal_3067) ) ;
    buf_clk new_AGEMA_reg_buffer_1619 ( .C (CLK), .D (new_AGEMA_signal_3070), .Q (new_AGEMA_signal_3071) ) ;
    buf_clk new_AGEMA_reg_buffer_1623 ( .C (CLK), .D (new_AGEMA_signal_3074), .Q (new_AGEMA_signal_3075) ) ;
    buf_clk new_AGEMA_reg_buffer_1627 ( .C (CLK), .D (new_AGEMA_signal_3078), .Q (new_AGEMA_signal_3079) ) ;
    buf_clk new_AGEMA_reg_buffer_1631 ( .C (CLK), .D (new_AGEMA_signal_3082), .Q (new_AGEMA_signal_3083) ) ;
    buf_clk new_AGEMA_reg_buffer_1635 ( .C (CLK), .D (new_AGEMA_signal_3086), .Q (new_AGEMA_signal_3087) ) ;
    buf_clk new_AGEMA_reg_buffer_1639 ( .C (CLK), .D (new_AGEMA_signal_3090), .Q (new_AGEMA_signal_3091) ) ;
    buf_clk new_AGEMA_reg_buffer_1643 ( .C (CLK), .D (new_AGEMA_signal_3094), .Q (new_AGEMA_signal_3095) ) ;
    buf_clk new_AGEMA_reg_buffer_1647 ( .C (CLK), .D (new_AGEMA_signal_3098), .Q (new_AGEMA_signal_3099) ) ;
    buf_clk new_AGEMA_reg_buffer_1651 ( .C (CLK), .D (new_AGEMA_signal_3102), .Q (new_AGEMA_signal_3103) ) ;
    buf_clk new_AGEMA_reg_buffer_1655 ( .C (CLK), .D (new_AGEMA_signal_3106), .Q (new_AGEMA_signal_3107) ) ;
    buf_clk new_AGEMA_reg_buffer_1659 ( .C (CLK), .D (new_AGEMA_signal_3110), .Q (new_AGEMA_signal_3111) ) ;
    buf_clk new_AGEMA_reg_buffer_1663 ( .C (CLK), .D (new_AGEMA_signal_3114), .Q (new_AGEMA_signal_3115) ) ;
    buf_clk new_AGEMA_reg_buffer_1667 ( .C (CLK), .D (new_AGEMA_signal_3118), .Q (new_AGEMA_signal_3119) ) ;
    buf_clk new_AGEMA_reg_buffer_1671 ( .C (CLK), .D (new_AGEMA_signal_3122), .Q (new_AGEMA_signal_3123) ) ;
    buf_clk new_AGEMA_reg_buffer_1675 ( .C (CLK), .D (new_AGEMA_signal_3126), .Q (new_AGEMA_signal_3127) ) ;
    buf_clk new_AGEMA_reg_buffer_1679 ( .C (CLK), .D (new_AGEMA_signal_3130), .Q (new_AGEMA_signal_3131) ) ;
    buf_clk new_AGEMA_reg_buffer_1683 ( .C (CLK), .D (new_AGEMA_signal_3134), .Q (new_AGEMA_signal_3135) ) ;
    buf_clk new_AGEMA_reg_buffer_1687 ( .C (CLK), .D (new_AGEMA_signal_3138), .Q (new_AGEMA_signal_3139) ) ;
    buf_clk new_AGEMA_reg_buffer_1691 ( .C (CLK), .D (new_AGEMA_signal_3142), .Q (new_AGEMA_signal_3143) ) ;
    buf_clk new_AGEMA_reg_buffer_1695 ( .C (CLK), .D (new_AGEMA_signal_3146), .Q (new_AGEMA_signal_3147) ) ;
    buf_clk new_AGEMA_reg_buffer_1699 ( .C (CLK), .D (new_AGEMA_signal_3150), .Q (new_AGEMA_signal_3151) ) ;
    buf_clk new_AGEMA_reg_buffer_1703 ( .C (CLK), .D (new_AGEMA_signal_3154), .Q (new_AGEMA_signal_3155) ) ;
    buf_clk new_AGEMA_reg_buffer_1707 ( .C (CLK), .D (new_AGEMA_signal_3158), .Q (new_AGEMA_signal_3159) ) ;
    buf_clk new_AGEMA_reg_buffer_1711 ( .C (CLK), .D (new_AGEMA_signal_3162), .Q (new_AGEMA_signal_3163) ) ;
    buf_clk new_AGEMA_reg_buffer_1715 ( .C (CLK), .D (new_AGEMA_signal_3166), .Q (new_AGEMA_signal_3167) ) ;
    buf_clk new_AGEMA_reg_buffer_1719 ( .C (CLK), .D (new_AGEMA_signal_3170), .Q (new_AGEMA_signal_3171) ) ;
    buf_clk new_AGEMA_reg_buffer_1723 ( .C (CLK), .D (new_AGEMA_signal_3174), .Q (new_AGEMA_signal_3175) ) ;
    buf_clk new_AGEMA_reg_buffer_1727 ( .C (CLK), .D (new_AGEMA_signal_3178), .Q (new_AGEMA_signal_3179) ) ;
    buf_clk new_AGEMA_reg_buffer_1731 ( .C (CLK), .D (new_AGEMA_signal_3182), .Q (new_AGEMA_signal_3183) ) ;
    buf_clk new_AGEMA_reg_buffer_1735 ( .C (CLK), .D (new_AGEMA_signal_3186), .Q (new_AGEMA_signal_3187) ) ;
    buf_clk new_AGEMA_reg_buffer_1739 ( .C (CLK), .D (new_AGEMA_signal_3190), .Q (new_AGEMA_signal_3191) ) ;
    buf_clk new_AGEMA_reg_buffer_1743 ( .C (CLK), .D (new_AGEMA_signal_3194), .Q (new_AGEMA_signal_3195) ) ;
    buf_clk new_AGEMA_reg_buffer_1747 ( .C (CLK), .D (new_AGEMA_signal_3198), .Q (new_AGEMA_signal_3199) ) ;
    buf_clk new_AGEMA_reg_buffer_1751 ( .C (CLK), .D (new_AGEMA_signal_3202), .Q (new_AGEMA_signal_3203) ) ;
    buf_clk new_AGEMA_reg_buffer_1755 ( .C (CLK), .D (new_AGEMA_signal_3206), .Q (new_AGEMA_signal_3207) ) ;
    buf_clk new_AGEMA_reg_buffer_1759 ( .C (CLK), .D (new_AGEMA_signal_3210), .Q (new_AGEMA_signal_3211) ) ;
    buf_clk new_AGEMA_reg_buffer_1763 ( .C (CLK), .D (new_AGEMA_signal_3214), .Q (new_AGEMA_signal_3215) ) ;
    buf_clk new_AGEMA_reg_buffer_1767 ( .C (CLK), .D (new_AGEMA_signal_3218), .Q (new_AGEMA_signal_3219) ) ;
    buf_clk new_AGEMA_reg_buffer_1771 ( .C (CLK), .D (new_AGEMA_signal_3222), .Q (new_AGEMA_signal_3223) ) ;
    buf_clk new_AGEMA_reg_buffer_1775 ( .C (CLK), .D (new_AGEMA_signal_3226), .Q (new_AGEMA_signal_3227) ) ;
    buf_clk new_AGEMA_reg_buffer_1779 ( .C (CLK), .D (new_AGEMA_signal_3230), .Q (new_AGEMA_signal_3231) ) ;
    buf_clk new_AGEMA_reg_buffer_1783 ( .C (CLK), .D (new_AGEMA_signal_3234), .Q (new_AGEMA_signal_3235) ) ;
    buf_clk new_AGEMA_reg_buffer_1787 ( .C (CLK), .D (new_AGEMA_signal_3238), .Q (new_AGEMA_signal_3239) ) ;
    buf_clk new_AGEMA_reg_buffer_1791 ( .C (CLK), .D (new_AGEMA_signal_3242), .Q (new_AGEMA_signal_3243) ) ;
    buf_clk new_AGEMA_reg_buffer_1795 ( .C (CLK), .D (new_AGEMA_signal_3246), .Q (new_AGEMA_signal_3247) ) ;
    buf_clk new_AGEMA_reg_buffer_1799 ( .C (CLK), .D (new_AGEMA_signal_3250), .Q (new_AGEMA_signal_3251) ) ;
    buf_clk new_AGEMA_reg_buffer_1803 ( .C (CLK), .D (new_AGEMA_signal_3254), .Q (new_AGEMA_signal_3255) ) ;
    buf_clk new_AGEMA_reg_buffer_1807 ( .C (CLK), .D (new_AGEMA_signal_3258), .Q (new_AGEMA_signal_3259) ) ;
    buf_clk new_AGEMA_reg_buffer_1811 ( .C (CLK), .D (new_AGEMA_signal_3262), .Q (new_AGEMA_signal_3263) ) ;
    buf_clk new_AGEMA_reg_buffer_1815 ( .C (CLK), .D (new_AGEMA_signal_3266), .Q (new_AGEMA_signal_3267) ) ;
    buf_clk new_AGEMA_reg_buffer_1819 ( .C (CLK), .D (new_AGEMA_signal_3270), .Q (new_AGEMA_signal_3271) ) ;
    buf_clk new_AGEMA_reg_buffer_1823 ( .C (CLK), .D (new_AGEMA_signal_3274), .Q (new_AGEMA_signal_3275) ) ;
    buf_clk new_AGEMA_reg_buffer_1827 ( .C (CLK), .D (new_AGEMA_signal_3278), .Q (new_AGEMA_signal_3279) ) ;
    buf_clk new_AGEMA_reg_buffer_1831 ( .C (CLK), .D (new_AGEMA_signal_3282), .Q (new_AGEMA_signal_3283) ) ;
    buf_clk new_AGEMA_reg_buffer_1835 ( .C (CLK), .D (new_AGEMA_signal_3286), .Q (new_AGEMA_signal_3287) ) ;
    buf_clk new_AGEMA_reg_buffer_1839 ( .C (CLK), .D (new_AGEMA_signal_3290), .Q (new_AGEMA_signal_3291) ) ;
    buf_clk new_AGEMA_reg_buffer_1843 ( .C (CLK), .D (new_AGEMA_signal_3294), .Q (new_AGEMA_signal_3295) ) ;
    buf_clk new_AGEMA_reg_buffer_1847 ( .C (CLK), .D (new_AGEMA_signal_3298), .Q (new_AGEMA_signal_3299) ) ;
    buf_clk new_AGEMA_reg_buffer_1851 ( .C (CLK), .D (new_AGEMA_signal_3302), .Q (new_AGEMA_signal_3303) ) ;
    buf_clk new_AGEMA_reg_buffer_1855 ( .C (CLK), .D (new_AGEMA_signal_3306), .Q (new_AGEMA_signal_3307) ) ;
    buf_clk new_AGEMA_reg_buffer_1859 ( .C (CLK), .D (new_AGEMA_signal_3310), .Q (new_AGEMA_signal_3311) ) ;
    buf_clk new_AGEMA_reg_buffer_1863 ( .C (CLK), .D (new_AGEMA_signal_3314), .Q (new_AGEMA_signal_3315) ) ;
    buf_clk new_AGEMA_reg_buffer_1867 ( .C (CLK), .D (new_AGEMA_signal_3318), .Q (new_AGEMA_signal_3319) ) ;
    buf_clk new_AGEMA_reg_buffer_1871 ( .C (CLK), .D (new_AGEMA_signal_3322), .Q (new_AGEMA_signal_3323) ) ;
    buf_clk new_AGEMA_reg_buffer_1875 ( .C (CLK), .D (new_AGEMA_signal_3326), .Q (new_AGEMA_signal_3327) ) ;
    buf_clk new_AGEMA_reg_buffer_1879 ( .C (CLK), .D (new_AGEMA_signal_3330), .Q (new_AGEMA_signal_3331) ) ;
    buf_clk new_AGEMA_reg_buffer_1883 ( .C (CLK), .D (new_AGEMA_signal_3334), .Q (new_AGEMA_signal_3335) ) ;
    buf_clk new_AGEMA_reg_buffer_1887 ( .C (CLK), .D (new_AGEMA_signal_3338), .Q (new_AGEMA_signal_3339) ) ;
    buf_clk new_AGEMA_reg_buffer_1891 ( .C (CLK), .D (new_AGEMA_signal_3342), .Q (new_AGEMA_signal_3343) ) ;
    buf_clk new_AGEMA_reg_buffer_1895 ( .C (CLK), .D (new_AGEMA_signal_3346), .Q (new_AGEMA_signal_3347) ) ;
    buf_clk new_AGEMA_reg_buffer_1899 ( .C (CLK), .D (new_AGEMA_signal_3350), .Q (new_AGEMA_signal_3351) ) ;
    buf_clk new_AGEMA_reg_buffer_1903 ( .C (CLK), .D (new_AGEMA_signal_3354), .Q (new_AGEMA_signal_3355) ) ;
    buf_clk new_AGEMA_reg_buffer_1907 ( .C (CLK), .D (new_AGEMA_signal_3358), .Q (new_AGEMA_signal_3359) ) ;
    buf_clk new_AGEMA_reg_buffer_1911 ( .C (CLK), .D (new_AGEMA_signal_3362), .Q (new_AGEMA_signal_3363) ) ;
    buf_clk new_AGEMA_reg_buffer_1915 ( .C (CLK), .D (new_AGEMA_signal_3366), .Q (new_AGEMA_signal_3367) ) ;
    buf_clk new_AGEMA_reg_buffer_1919 ( .C (CLK), .D (new_AGEMA_signal_3370), .Q (new_AGEMA_signal_3371) ) ;
    buf_clk new_AGEMA_reg_buffer_1923 ( .C (CLK), .D (new_AGEMA_signal_3374), .Q (new_AGEMA_signal_3375) ) ;
    buf_clk new_AGEMA_reg_buffer_1927 ( .C (CLK), .D (new_AGEMA_signal_3378), .Q (new_AGEMA_signal_3379) ) ;
    buf_clk new_AGEMA_reg_buffer_1931 ( .C (CLK), .D (new_AGEMA_signal_3382), .Q (new_AGEMA_signal_3383) ) ;
    buf_clk new_AGEMA_reg_buffer_1935 ( .C (CLK), .D (new_AGEMA_signal_3386), .Q (new_AGEMA_signal_3387) ) ;
    buf_clk new_AGEMA_reg_buffer_1939 ( .C (CLK), .D (new_AGEMA_signal_3390), .Q (new_AGEMA_signal_3391) ) ;
    buf_clk new_AGEMA_reg_buffer_1943 ( .C (CLK), .D (new_AGEMA_signal_3394), .Q (new_AGEMA_signal_3395) ) ;
    buf_clk new_AGEMA_reg_buffer_1947 ( .C (CLK), .D (new_AGEMA_signal_3398), .Q (new_AGEMA_signal_3399) ) ;
    buf_clk new_AGEMA_reg_buffer_1951 ( .C (CLK), .D (new_AGEMA_signal_3402), .Q (new_AGEMA_signal_3403) ) ;
    buf_clk new_AGEMA_reg_buffer_1955 ( .C (CLK), .D (new_AGEMA_signal_3406), .Q (new_AGEMA_signal_3407) ) ;
    buf_clk new_AGEMA_reg_buffer_1959 ( .C (CLK), .D (new_AGEMA_signal_3410), .Q (new_AGEMA_signal_3411) ) ;
    buf_clk new_AGEMA_reg_buffer_1963 ( .C (CLK), .D (new_AGEMA_signal_3414), .Q (new_AGEMA_signal_3415) ) ;
    buf_clk new_AGEMA_reg_buffer_1967 ( .C (CLK), .D (new_AGEMA_signal_3418), .Q (new_AGEMA_signal_3419) ) ;
    buf_clk new_AGEMA_reg_buffer_1971 ( .C (CLK), .D (new_AGEMA_signal_3422), .Q (new_AGEMA_signal_3423) ) ;
    buf_clk new_AGEMA_reg_buffer_1975 ( .C (CLK), .D (new_AGEMA_signal_3426), .Q (new_AGEMA_signal_3427) ) ;
    buf_clk new_AGEMA_reg_buffer_1979 ( .C (CLK), .D (new_AGEMA_signal_3430), .Q (new_AGEMA_signal_3431) ) ;
    buf_clk new_AGEMA_reg_buffer_1983 ( .C (CLK), .D (new_AGEMA_signal_3434), .Q (new_AGEMA_signal_3435) ) ;
    buf_clk new_AGEMA_reg_buffer_1987 ( .C (CLK), .D (new_AGEMA_signal_3438), .Q (new_AGEMA_signal_3439) ) ;
    buf_clk new_AGEMA_reg_buffer_1991 ( .C (CLK), .D (new_AGEMA_signal_3442), .Q (new_AGEMA_signal_3443) ) ;
    buf_clk new_AGEMA_reg_buffer_1995 ( .C (CLK), .D (new_AGEMA_signal_3446), .Q (new_AGEMA_signal_3447) ) ;
    buf_clk new_AGEMA_reg_buffer_1999 ( .C (CLK), .D (new_AGEMA_signal_3450), .Q (new_AGEMA_signal_3451) ) ;
    buf_clk new_AGEMA_reg_buffer_2003 ( .C (CLK), .D (new_AGEMA_signal_3454), .Q (new_AGEMA_signal_3455) ) ;
    buf_clk new_AGEMA_reg_buffer_2007 ( .C (CLK), .D (new_AGEMA_signal_3458), .Q (new_AGEMA_signal_3459) ) ;
    buf_clk new_AGEMA_reg_buffer_2011 ( .C (CLK), .D (new_AGEMA_signal_3462), .Q (new_AGEMA_signal_3463) ) ;
    buf_clk new_AGEMA_reg_buffer_2015 ( .C (CLK), .D (new_AGEMA_signal_3466), .Q (new_AGEMA_signal_3467) ) ;
    buf_clk new_AGEMA_reg_buffer_2019 ( .C (CLK), .D (new_AGEMA_signal_3470), .Q (new_AGEMA_signal_3471) ) ;
    buf_clk new_AGEMA_reg_buffer_2023 ( .C (CLK), .D (new_AGEMA_signal_3474), .Q (new_AGEMA_signal_3475) ) ;
    buf_clk new_AGEMA_reg_buffer_2027 ( .C (CLK), .D (new_AGEMA_signal_3478), .Q (new_AGEMA_signal_3479) ) ;
    buf_clk new_AGEMA_reg_buffer_2031 ( .C (CLK), .D (new_AGEMA_signal_3482), .Q (new_AGEMA_signal_3483) ) ;
    buf_clk new_AGEMA_reg_buffer_2035 ( .C (CLK), .D (new_AGEMA_signal_3486), .Q (new_AGEMA_signal_3487) ) ;
    buf_clk new_AGEMA_reg_buffer_2039 ( .C (CLK), .D (new_AGEMA_signal_3490), .Q (new_AGEMA_signal_3491) ) ;
    buf_clk new_AGEMA_reg_buffer_2043 ( .C (CLK), .D (new_AGEMA_signal_3494), .Q (new_AGEMA_signal_3495) ) ;
    buf_clk new_AGEMA_reg_buffer_2047 ( .C (CLK), .D (new_AGEMA_signal_3498), .Q (new_AGEMA_signal_3499) ) ;
    buf_clk new_AGEMA_reg_buffer_2051 ( .C (CLK), .D (new_AGEMA_signal_3502), .Q (new_AGEMA_signal_3503) ) ;
    buf_clk new_AGEMA_reg_buffer_2055 ( .C (CLK), .D (new_AGEMA_signal_3506), .Q (new_AGEMA_signal_3507) ) ;
    buf_clk new_AGEMA_reg_buffer_2059 ( .C (CLK), .D (new_AGEMA_signal_3510), .Q (new_AGEMA_signal_3511) ) ;
    buf_clk new_AGEMA_reg_buffer_2063 ( .C (CLK), .D (new_AGEMA_signal_3514), .Q (new_AGEMA_signal_3515) ) ;
    buf_clk new_AGEMA_reg_buffer_2067 ( .C (CLK), .D (new_AGEMA_signal_3518), .Q (new_AGEMA_signal_3519) ) ;
    buf_clk new_AGEMA_reg_buffer_2071 ( .C (CLK), .D (new_AGEMA_signal_3522), .Q (new_AGEMA_signal_3523) ) ;
    buf_clk new_AGEMA_reg_buffer_2075 ( .C (CLK), .D (new_AGEMA_signal_3526), .Q (new_AGEMA_signal_3527) ) ;
    buf_clk new_AGEMA_reg_buffer_2079 ( .C (CLK), .D (new_AGEMA_signal_3530), .Q (new_AGEMA_signal_3531) ) ;
    buf_clk new_AGEMA_reg_buffer_2083 ( .C (CLK), .D (new_AGEMA_signal_3534), .Q (new_AGEMA_signal_3535) ) ;
    buf_clk new_AGEMA_reg_buffer_2087 ( .C (CLK), .D (new_AGEMA_signal_3538), .Q (new_AGEMA_signal_3539) ) ;
    buf_clk new_AGEMA_reg_buffer_2091 ( .C (CLK), .D (new_AGEMA_signal_3542), .Q (new_AGEMA_signal_3543) ) ;
    buf_clk new_AGEMA_reg_buffer_2095 ( .C (CLK), .D (new_AGEMA_signal_3546), .Q (new_AGEMA_signal_3547) ) ;
    buf_clk new_AGEMA_reg_buffer_2099 ( .C (CLK), .D (new_AGEMA_signal_3550), .Q (new_AGEMA_signal_3551) ) ;
    buf_clk new_AGEMA_reg_buffer_2103 ( .C (CLK), .D (new_AGEMA_signal_3554), .Q (new_AGEMA_signal_3555) ) ;
    buf_clk new_AGEMA_reg_buffer_2107 ( .C (CLK), .D (new_AGEMA_signal_3558), .Q (new_AGEMA_signal_3559) ) ;
    buf_clk new_AGEMA_reg_buffer_2111 ( .C (CLK), .D (new_AGEMA_signal_3562), .Q (new_AGEMA_signal_3563) ) ;
    buf_clk new_AGEMA_reg_buffer_2115 ( .C (CLK), .D (new_AGEMA_signal_3566), .Q (new_AGEMA_signal_3567) ) ;
    buf_clk new_AGEMA_reg_buffer_2119 ( .C (CLK), .D (new_AGEMA_signal_3570), .Q (new_AGEMA_signal_3571) ) ;
    buf_clk new_AGEMA_reg_buffer_2123 ( .C (CLK), .D (new_AGEMA_signal_3574), .Q (new_AGEMA_signal_3575) ) ;
    buf_clk new_AGEMA_reg_buffer_2127 ( .C (CLK), .D (new_AGEMA_signal_3578), .Q (new_AGEMA_signal_3579) ) ;
    buf_clk new_AGEMA_reg_buffer_2131 ( .C (CLK), .D (new_AGEMA_signal_3582), .Q (new_AGEMA_signal_3583) ) ;
    buf_clk new_AGEMA_reg_buffer_2135 ( .C (CLK), .D (new_AGEMA_signal_3586), .Q (new_AGEMA_signal_3587) ) ;
    buf_clk new_AGEMA_reg_buffer_2139 ( .C (CLK), .D (new_AGEMA_signal_3590), .Q (new_AGEMA_signal_3591) ) ;
    buf_clk new_AGEMA_reg_buffer_2143 ( .C (CLK), .D (new_AGEMA_signal_3594), .Q (new_AGEMA_signal_3595) ) ;
    buf_clk new_AGEMA_reg_buffer_2147 ( .C (CLK), .D (new_AGEMA_signal_3598), .Q (new_AGEMA_signal_3599) ) ;
    buf_clk new_AGEMA_reg_buffer_2151 ( .C (CLK), .D (new_AGEMA_signal_3602), .Q (new_AGEMA_signal_3603) ) ;
    buf_clk new_AGEMA_reg_buffer_2155 ( .C (CLK), .D (new_AGEMA_signal_3606), .Q (new_AGEMA_signal_3607) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (CLK), .D (new_AGEMA_signal_3610), .Q (new_AGEMA_signal_3611) ) ;
    buf_clk new_AGEMA_reg_buffer_2163 ( .C (CLK), .D (new_AGEMA_signal_3614), .Q (new_AGEMA_signal_3615) ) ;
    buf_clk new_AGEMA_reg_buffer_2167 ( .C (CLK), .D (new_AGEMA_signal_3618), .Q (new_AGEMA_signal_3619) ) ;
    buf_clk new_AGEMA_reg_buffer_2171 ( .C (CLK), .D (new_AGEMA_signal_3622), .Q (new_AGEMA_signal_3623) ) ;
    buf_clk new_AGEMA_reg_buffer_2175 ( .C (CLK), .D (new_AGEMA_signal_3626), .Q (new_AGEMA_signal_3627) ) ;
    buf_clk new_AGEMA_reg_buffer_2179 ( .C (CLK), .D (new_AGEMA_signal_3630), .Q (new_AGEMA_signal_3631) ) ;
    buf_clk new_AGEMA_reg_buffer_2183 ( .C (CLK), .D (new_AGEMA_signal_3634), .Q (new_AGEMA_signal_3635) ) ;
    buf_clk new_AGEMA_reg_buffer_2187 ( .C (CLK), .D (new_AGEMA_signal_3638), .Q (new_AGEMA_signal_3639) ) ;
    buf_clk new_AGEMA_reg_buffer_2191 ( .C (CLK), .D (new_AGEMA_signal_3642), .Q (new_AGEMA_signal_3643) ) ;
    buf_clk new_AGEMA_reg_buffer_2195 ( .C (CLK), .D (new_AGEMA_signal_3646), .Q (new_AGEMA_signal_3647) ) ;
    buf_clk new_AGEMA_reg_buffer_2199 ( .C (CLK), .D (new_AGEMA_signal_3650), .Q (new_AGEMA_signal_3651) ) ;
    buf_clk new_AGEMA_reg_buffer_2203 ( .C (CLK), .D (new_AGEMA_signal_3654), .Q (new_AGEMA_signal_3655) ) ;
    buf_clk new_AGEMA_reg_buffer_2207 ( .C (CLK), .D (new_AGEMA_signal_3658), .Q (new_AGEMA_signal_3659) ) ;
    buf_clk new_AGEMA_reg_buffer_2211 ( .C (CLK), .D (new_AGEMA_signal_3662), .Q (new_AGEMA_signal_3663) ) ;
    buf_clk new_AGEMA_reg_buffer_2215 ( .C (CLK), .D (new_AGEMA_signal_3666), .Q (new_AGEMA_signal_3667) ) ;
    buf_clk new_AGEMA_reg_buffer_2219 ( .C (CLK), .D (new_AGEMA_signal_3670), .Q (new_AGEMA_signal_3671) ) ;
    buf_clk new_AGEMA_reg_buffer_2223 ( .C (CLK), .D (new_AGEMA_signal_3674), .Q (new_AGEMA_signal_3675) ) ;
    buf_clk new_AGEMA_reg_buffer_2227 ( .C (CLK), .D (new_AGEMA_signal_3678), .Q (new_AGEMA_signal_3679) ) ;
    buf_clk new_AGEMA_reg_buffer_2231 ( .C (CLK), .D (new_AGEMA_signal_3682), .Q (new_AGEMA_signal_3683) ) ;
    buf_clk new_AGEMA_reg_buffer_2235 ( .C (CLK), .D (new_AGEMA_signal_3686), .Q (new_AGEMA_signal_3687) ) ;
    buf_clk new_AGEMA_reg_buffer_2239 ( .C (CLK), .D (new_AGEMA_signal_3690), .Q (new_AGEMA_signal_3691) ) ;
    buf_clk new_AGEMA_reg_buffer_2243 ( .C (CLK), .D (new_AGEMA_signal_3694), .Q (new_AGEMA_signal_3695) ) ;
    buf_clk new_AGEMA_reg_buffer_2247 ( .C (CLK), .D (new_AGEMA_signal_3698), .Q (new_AGEMA_signal_3699) ) ;
    buf_clk new_AGEMA_reg_buffer_2251 ( .C (CLK), .D (new_AGEMA_signal_3702), .Q (new_AGEMA_signal_3703) ) ;
    buf_clk new_AGEMA_reg_buffer_2255 ( .C (CLK), .D (new_AGEMA_signal_3706), .Q (new_AGEMA_signal_3707) ) ;
    buf_clk new_AGEMA_reg_buffer_2259 ( .C (CLK), .D (new_AGEMA_signal_3710), .Q (new_AGEMA_signal_3711) ) ;
    buf_clk new_AGEMA_reg_buffer_2263 ( .C (CLK), .D (new_AGEMA_signal_3714), .Q (new_AGEMA_signal_3715) ) ;
    buf_clk new_AGEMA_reg_buffer_2267 ( .C (CLK), .D (new_AGEMA_signal_3718), .Q (new_AGEMA_signal_3719) ) ;
    buf_clk new_AGEMA_reg_buffer_2271 ( .C (CLK), .D (new_AGEMA_signal_3722), .Q (new_AGEMA_signal_3723) ) ;
    buf_clk new_AGEMA_reg_buffer_2275 ( .C (CLK), .D (new_AGEMA_signal_3726), .Q (new_AGEMA_signal_3727) ) ;
    buf_clk new_AGEMA_reg_buffer_2279 ( .C (CLK), .D (new_AGEMA_signal_3730), .Q (new_AGEMA_signal_3731) ) ;
    buf_clk new_AGEMA_reg_buffer_2283 ( .C (CLK), .D (new_AGEMA_signal_3734), .Q (new_AGEMA_signal_3735) ) ;
    buf_clk new_AGEMA_reg_buffer_2287 ( .C (CLK), .D (new_AGEMA_signal_3738), .Q (new_AGEMA_signal_3739) ) ;
    buf_clk new_AGEMA_reg_buffer_2291 ( .C (CLK), .D (new_AGEMA_signal_3742), .Q (new_AGEMA_signal_3743) ) ;
    buf_clk new_AGEMA_reg_buffer_2295 ( .C (CLK), .D (new_AGEMA_signal_3746), .Q (new_AGEMA_signal_3747) ) ;
    buf_clk new_AGEMA_reg_buffer_2299 ( .C (CLK), .D (new_AGEMA_signal_3750), .Q (new_AGEMA_signal_3751) ) ;
    buf_clk new_AGEMA_reg_buffer_2303 ( .C (CLK), .D (new_AGEMA_signal_3754), .Q (new_AGEMA_signal_3755) ) ;
    buf_clk new_AGEMA_reg_buffer_2307 ( .C (CLK), .D (new_AGEMA_signal_3758), .Q (new_AGEMA_signal_3759) ) ;
    buf_clk new_AGEMA_reg_buffer_2311 ( .C (CLK), .D (new_AGEMA_signal_3762), .Q (new_AGEMA_signal_3763) ) ;
    buf_clk new_AGEMA_reg_buffer_2315 ( .C (CLK), .D (new_AGEMA_signal_3766), .Q (new_AGEMA_signal_3767) ) ;
    buf_clk new_AGEMA_reg_buffer_2319 ( .C (CLK), .D (new_AGEMA_signal_3770), .Q (new_AGEMA_signal_3771) ) ;
    buf_clk new_AGEMA_reg_buffer_2323 ( .C (CLK), .D (new_AGEMA_signal_3774), .Q (new_AGEMA_signal_3775) ) ;
    buf_clk new_AGEMA_reg_buffer_2327 ( .C (CLK), .D (new_AGEMA_signal_3778), .Q (new_AGEMA_signal_3779) ) ;
    buf_clk new_AGEMA_reg_buffer_2331 ( .C (CLK), .D (new_AGEMA_signal_3782), .Q (new_AGEMA_signal_3783) ) ;
    buf_clk new_AGEMA_reg_buffer_2335 ( .C (CLK), .D (new_AGEMA_signal_3786), .Q (new_AGEMA_signal_3787) ) ;
    buf_clk new_AGEMA_reg_buffer_2339 ( .C (CLK), .D (new_AGEMA_signal_3790), .Q (new_AGEMA_signal_3791) ) ;
    buf_clk new_AGEMA_reg_buffer_2343 ( .C (CLK), .D (new_AGEMA_signal_3794), .Q (new_AGEMA_signal_3795) ) ;
    buf_clk new_AGEMA_reg_buffer_2347 ( .C (CLK), .D (new_AGEMA_signal_3798), .Q (new_AGEMA_signal_3799) ) ;
    buf_clk new_AGEMA_reg_buffer_2351 ( .C (CLK), .D (new_AGEMA_signal_3802), .Q (new_AGEMA_signal_3803) ) ;
    buf_clk new_AGEMA_reg_buffer_2355 ( .C (CLK), .D (new_AGEMA_signal_3806), .Q (new_AGEMA_signal_3807) ) ;
    buf_clk new_AGEMA_reg_buffer_2359 ( .C (CLK), .D (new_AGEMA_signal_3810), .Q (new_AGEMA_signal_3811) ) ;
    buf_clk new_AGEMA_reg_buffer_2363 ( .C (CLK), .D (new_AGEMA_signal_3814), .Q (new_AGEMA_signal_3815) ) ;
    buf_clk new_AGEMA_reg_buffer_2373 ( .C (CLK), .D (new_AGEMA_signal_3824), .Q (new_AGEMA_signal_3825) ) ;
    buf_clk new_AGEMA_reg_buffer_2375 ( .C (CLK), .D (new_AGEMA_signal_3826), .Q (new_AGEMA_signal_3827) ) ;
    buf_clk new_AGEMA_reg_buffer_2379 ( .C (CLK), .D (new_AGEMA_signal_3830), .Q (new_AGEMA_signal_3831) ) ;
    buf_clk new_AGEMA_reg_buffer_2383 ( .C (CLK), .D (new_AGEMA_signal_3834), .Q (new_AGEMA_signal_3835) ) ;
    buf_clk new_AGEMA_reg_buffer_2387 ( .C (CLK), .D (new_AGEMA_signal_3838), .Q (new_AGEMA_signal_3839) ) ;
    buf_clk new_AGEMA_reg_buffer_2391 ( .C (CLK), .D (new_AGEMA_signal_3842), .Q (new_AGEMA_signal_3843) ) ;
    buf_clk new_AGEMA_reg_buffer_2393 ( .C (CLK), .D (new_AGEMA_signal_3844), .Q (new_AGEMA_signal_3845) ) ;
    buf_clk new_AGEMA_reg_buffer_2395 ( .C (CLK), .D (new_AGEMA_signal_3846), .Q (new_AGEMA_signal_3847) ) ;
    buf_clk new_AGEMA_reg_buffer_2405 ( .C (CLK), .D (new_AGEMA_signal_3856), .Q (new_AGEMA_signal_3857) ) ;
    buf_clk new_AGEMA_reg_buffer_2407 ( .C (CLK), .D (new_AGEMA_signal_3858), .Q (new_AGEMA_signal_3859) ) ;
    buf_clk new_AGEMA_reg_buffer_2411 ( .C (CLK), .D (new_AGEMA_signal_3862), .Q (new_AGEMA_signal_3863) ) ;
    buf_clk new_AGEMA_reg_buffer_2415 ( .C (CLK), .D (new_AGEMA_signal_3866), .Q (new_AGEMA_signal_3867) ) ;
    buf_clk new_AGEMA_reg_buffer_2419 ( .C (CLK), .D (new_AGEMA_signal_3870), .Q (new_AGEMA_signal_3871) ) ;
    buf_clk new_AGEMA_reg_buffer_2423 ( .C (CLK), .D (new_AGEMA_signal_3874), .Q (new_AGEMA_signal_3875) ) ;
    buf_clk new_AGEMA_reg_buffer_2425 ( .C (CLK), .D (new_AGEMA_signal_3876), .Q (new_AGEMA_signal_3877) ) ;
    buf_clk new_AGEMA_reg_buffer_2427 ( .C (CLK), .D (new_AGEMA_signal_3878), .Q (new_AGEMA_signal_3879) ) ;
    buf_clk new_AGEMA_reg_buffer_2437 ( .C (CLK), .D (new_AGEMA_signal_3888), .Q (new_AGEMA_signal_3889) ) ;
    buf_clk new_AGEMA_reg_buffer_2439 ( .C (CLK), .D (new_AGEMA_signal_3890), .Q (new_AGEMA_signal_3891) ) ;
    buf_clk new_AGEMA_reg_buffer_2443 ( .C (CLK), .D (new_AGEMA_signal_3894), .Q (new_AGEMA_signal_3895) ) ;
    buf_clk new_AGEMA_reg_buffer_2447 ( .C (CLK), .D (new_AGEMA_signal_3898), .Q (new_AGEMA_signal_3899) ) ;
    buf_clk new_AGEMA_reg_buffer_2449 ( .C (CLK), .D (new_AGEMA_signal_3900), .Q (new_AGEMA_signal_3901) ) ;
    buf_clk new_AGEMA_reg_buffer_2451 ( .C (CLK), .D (new_AGEMA_signal_3902), .Q (new_AGEMA_signal_3903) ) ;
    buf_clk new_AGEMA_reg_buffer_2461 ( .C (CLK), .D (new_AGEMA_signal_3912), .Q (new_AGEMA_signal_3913) ) ;
    buf_clk new_AGEMA_reg_buffer_2463 ( .C (CLK), .D (new_AGEMA_signal_3914), .Q (new_AGEMA_signal_3915) ) ;
    buf_clk new_AGEMA_reg_buffer_2467 ( .C (CLK), .D (new_AGEMA_signal_3918), .Q (new_AGEMA_signal_3919) ) ;
    buf_clk new_AGEMA_reg_buffer_2471 ( .C (CLK), .D (new_AGEMA_signal_3922), .Q (new_AGEMA_signal_3923) ) ;
    buf_clk new_AGEMA_reg_buffer_2473 ( .C (CLK), .D (new_AGEMA_signal_3924), .Q (new_AGEMA_signal_3925) ) ;
    buf_clk new_AGEMA_reg_buffer_2475 ( .C (CLK), .D (new_AGEMA_signal_3926), .Q (new_AGEMA_signal_3927) ) ;
    buf_clk new_AGEMA_reg_buffer_2485 ( .C (CLK), .D (new_AGEMA_signal_3936), .Q (new_AGEMA_signal_3937) ) ;
    buf_clk new_AGEMA_reg_buffer_2487 ( .C (CLK), .D (new_AGEMA_signal_3938), .Q (new_AGEMA_signal_3939) ) ;
    buf_clk new_AGEMA_reg_buffer_2491 ( .C (CLK), .D (new_AGEMA_signal_3942), .Q (new_AGEMA_signal_3943) ) ;
    buf_clk new_AGEMA_reg_buffer_2495 ( .C (CLK), .D (new_AGEMA_signal_3946), .Q (new_AGEMA_signal_3947) ) ;
    buf_clk new_AGEMA_reg_buffer_2499 ( .C (CLK), .D (new_AGEMA_signal_3950), .Q (new_AGEMA_signal_3951) ) ;
    buf_clk new_AGEMA_reg_buffer_2503 ( .C (CLK), .D (new_AGEMA_signal_3954), .Q (new_AGEMA_signal_3955) ) ;
    buf_clk new_AGEMA_reg_buffer_2505 ( .C (CLK), .D (new_AGEMA_signal_3956), .Q (new_AGEMA_signal_3957) ) ;
    buf_clk new_AGEMA_reg_buffer_2507 ( .C (CLK), .D (new_AGEMA_signal_3958), .Q (new_AGEMA_signal_3959) ) ;
    buf_clk new_AGEMA_reg_buffer_2517 ( .C (CLK), .D (new_AGEMA_signal_3968), .Q (new_AGEMA_signal_3969) ) ;
    buf_clk new_AGEMA_reg_buffer_2519 ( .C (CLK), .D (new_AGEMA_signal_3970), .Q (new_AGEMA_signal_3971) ) ;
    buf_clk new_AGEMA_reg_buffer_2523 ( .C (CLK), .D (new_AGEMA_signal_3974), .Q (new_AGEMA_signal_3975) ) ;
    buf_clk new_AGEMA_reg_buffer_2527 ( .C (CLK), .D (new_AGEMA_signal_3978), .Q (new_AGEMA_signal_3979) ) ;
    buf_clk new_AGEMA_reg_buffer_2531 ( .C (CLK), .D (new_AGEMA_signal_3982), .Q (new_AGEMA_signal_3983) ) ;
    buf_clk new_AGEMA_reg_buffer_2535 ( .C (CLK), .D (new_AGEMA_signal_3986), .Q (new_AGEMA_signal_3987) ) ;
    buf_clk new_AGEMA_reg_buffer_2537 ( .C (CLK), .D (new_AGEMA_signal_3988), .Q (new_AGEMA_signal_3989) ) ;
    buf_clk new_AGEMA_reg_buffer_2539 ( .C (CLK), .D (new_AGEMA_signal_3990), .Q (new_AGEMA_signal_3991) ) ;
    buf_clk new_AGEMA_reg_buffer_2549 ( .C (CLK), .D (new_AGEMA_signal_4000), .Q (new_AGEMA_signal_4001) ) ;
    buf_clk new_AGEMA_reg_buffer_2551 ( .C (CLK), .D (new_AGEMA_signal_4002), .Q (new_AGEMA_signal_4003) ) ;
    buf_clk new_AGEMA_reg_buffer_2555 ( .C (CLK), .D (new_AGEMA_signal_4006), .Q (new_AGEMA_signal_4007) ) ;
    buf_clk new_AGEMA_reg_buffer_2559 ( .C (CLK), .D (new_AGEMA_signal_4010), .Q (new_AGEMA_signal_4011) ) ;
    buf_clk new_AGEMA_reg_buffer_2561 ( .C (CLK), .D (new_AGEMA_signal_4012), .Q (new_AGEMA_signal_4013) ) ;
    buf_clk new_AGEMA_reg_buffer_2563 ( .C (CLK), .D (new_AGEMA_signal_4014), .Q (new_AGEMA_signal_4015) ) ;
    buf_clk new_AGEMA_reg_buffer_2573 ( .C (CLK), .D (new_AGEMA_signal_4024), .Q (new_AGEMA_signal_4025) ) ;
    buf_clk new_AGEMA_reg_buffer_2575 ( .C (CLK), .D (new_AGEMA_signal_4026), .Q (new_AGEMA_signal_4027) ) ;
    buf_clk new_AGEMA_reg_buffer_2579 ( .C (CLK), .D (new_AGEMA_signal_4030), .Q (new_AGEMA_signal_4031) ) ;
    buf_clk new_AGEMA_reg_buffer_2583 ( .C (CLK), .D (new_AGEMA_signal_4034), .Q (new_AGEMA_signal_4035) ) ;
    buf_clk new_AGEMA_reg_buffer_2585 ( .C (CLK), .D (new_AGEMA_signal_4036), .Q (new_AGEMA_signal_4037) ) ;
    buf_clk new_AGEMA_reg_buffer_2587 ( .C (CLK), .D (new_AGEMA_signal_4038), .Q (new_AGEMA_signal_4039) ) ;
    buf_clk new_AGEMA_reg_buffer_2597 ( .C (CLK), .D (new_AGEMA_signal_4048), .Q (new_AGEMA_signal_4049) ) ;
    buf_clk new_AGEMA_reg_buffer_2599 ( .C (CLK), .D (new_AGEMA_signal_4050), .Q (new_AGEMA_signal_4051) ) ;
    buf_clk new_AGEMA_reg_buffer_2603 ( .C (CLK), .D (new_AGEMA_signal_4054), .Q (new_AGEMA_signal_4055) ) ;
    buf_clk new_AGEMA_reg_buffer_2607 ( .C (CLK), .D (new_AGEMA_signal_4058), .Q (new_AGEMA_signal_4059) ) ;
    buf_clk new_AGEMA_reg_buffer_2611 ( .C (CLK), .D (new_AGEMA_signal_4062), .Q (new_AGEMA_signal_4063) ) ;
    buf_clk new_AGEMA_reg_buffer_2615 ( .C (CLK), .D (new_AGEMA_signal_4066), .Q (new_AGEMA_signal_4067) ) ;
    buf_clk new_AGEMA_reg_buffer_2617 ( .C (CLK), .D (new_AGEMA_signal_4068), .Q (new_AGEMA_signal_4069) ) ;
    buf_clk new_AGEMA_reg_buffer_2619 ( .C (CLK), .D (new_AGEMA_signal_4070), .Q (new_AGEMA_signal_4071) ) ;
    buf_clk new_AGEMA_reg_buffer_2629 ( .C (CLK), .D (new_AGEMA_signal_4080), .Q (new_AGEMA_signal_4081) ) ;
    buf_clk new_AGEMA_reg_buffer_2631 ( .C (CLK), .D (new_AGEMA_signal_4082), .Q (new_AGEMA_signal_4083) ) ;
    buf_clk new_AGEMA_reg_buffer_2635 ( .C (CLK), .D (new_AGEMA_signal_4086), .Q (new_AGEMA_signal_4087) ) ;
    buf_clk new_AGEMA_reg_buffer_2639 ( .C (CLK), .D (new_AGEMA_signal_4090), .Q (new_AGEMA_signal_4091) ) ;
    buf_clk new_AGEMA_reg_buffer_2643 ( .C (CLK), .D (new_AGEMA_signal_4094), .Q (new_AGEMA_signal_4095) ) ;
    buf_clk new_AGEMA_reg_buffer_2647 ( .C (CLK), .D (new_AGEMA_signal_4098), .Q (new_AGEMA_signal_4099) ) ;
    buf_clk new_AGEMA_reg_buffer_2649 ( .C (CLK), .D (new_AGEMA_signal_4100), .Q (new_AGEMA_signal_4101) ) ;
    buf_clk new_AGEMA_reg_buffer_2651 ( .C (CLK), .D (new_AGEMA_signal_4102), .Q (new_AGEMA_signal_4103) ) ;
    buf_clk new_AGEMA_reg_buffer_2661 ( .C (CLK), .D (new_AGEMA_signal_4112), .Q (new_AGEMA_signal_4113) ) ;
    buf_clk new_AGEMA_reg_buffer_2663 ( .C (CLK), .D (new_AGEMA_signal_4114), .Q (new_AGEMA_signal_4115) ) ;
    buf_clk new_AGEMA_reg_buffer_2667 ( .C (CLK), .D (new_AGEMA_signal_4118), .Q (new_AGEMA_signal_4119) ) ;
    buf_clk new_AGEMA_reg_buffer_2671 ( .C (CLK), .D (new_AGEMA_signal_4122), .Q (new_AGEMA_signal_4123) ) ;
    buf_clk new_AGEMA_reg_buffer_2673 ( .C (CLK), .D (new_AGEMA_signal_4124), .Q (new_AGEMA_signal_4125) ) ;
    buf_clk new_AGEMA_reg_buffer_2675 ( .C (CLK), .D (new_AGEMA_signal_4126), .Q (new_AGEMA_signal_4127) ) ;
    buf_clk new_AGEMA_reg_buffer_2685 ( .C (CLK), .D (new_AGEMA_signal_4136), .Q (new_AGEMA_signal_4137) ) ;
    buf_clk new_AGEMA_reg_buffer_2687 ( .C (CLK), .D (new_AGEMA_signal_4138), .Q (new_AGEMA_signal_4139) ) ;
    buf_clk new_AGEMA_reg_buffer_2691 ( .C (CLK), .D (new_AGEMA_signal_4142), .Q (new_AGEMA_signal_4143) ) ;
    buf_clk new_AGEMA_reg_buffer_2695 ( .C (CLK), .D (new_AGEMA_signal_4146), .Q (new_AGEMA_signal_4147) ) ;
    buf_clk new_AGEMA_reg_buffer_2697 ( .C (CLK), .D (new_AGEMA_signal_4148), .Q (new_AGEMA_signal_4149) ) ;
    buf_clk new_AGEMA_reg_buffer_2699 ( .C (CLK), .D (new_AGEMA_signal_4150), .Q (new_AGEMA_signal_4151) ) ;
    buf_clk new_AGEMA_reg_buffer_2709 ( .C (CLK), .D (new_AGEMA_signal_4160), .Q (new_AGEMA_signal_4161) ) ;
    buf_clk new_AGEMA_reg_buffer_2711 ( .C (CLK), .D (new_AGEMA_signal_4162), .Q (new_AGEMA_signal_4163) ) ;
    buf_clk new_AGEMA_reg_buffer_2715 ( .C (CLK), .D (new_AGEMA_signal_4166), .Q (new_AGEMA_signal_4167) ) ;
    buf_clk new_AGEMA_reg_buffer_2719 ( .C (CLK), .D (new_AGEMA_signal_4170), .Q (new_AGEMA_signal_4171) ) ;
    buf_clk new_AGEMA_reg_buffer_2723 ( .C (CLK), .D (new_AGEMA_signal_4174), .Q (new_AGEMA_signal_4175) ) ;
    buf_clk new_AGEMA_reg_buffer_2727 ( .C (CLK), .D (new_AGEMA_signal_4178), .Q (new_AGEMA_signal_4179) ) ;
    buf_clk new_AGEMA_reg_buffer_2729 ( .C (CLK), .D (new_AGEMA_signal_4180), .Q (new_AGEMA_signal_4181) ) ;
    buf_clk new_AGEMA_reg_buffer_2731 ( .C (CLK), .D (new_AGEMA_signal_4182), .Q (new_AGEMA_signal_4183) ) ;
    buf_clk new_AGEMA_reg_buffer_2741 ( .C (CLK), .D (new_AGEMA_signal_4192), .Q (new_AGEMA_signal_4193) ) ;
    buf_clk new_AGEMA_reg_buffer_2743 ( .C (CLK), .D (new_AGEMA_signal_4194), .Q (new_AGEMA_signal_4195) ) ;
    buf_clk new_AGEMA_reg_buffer_2747 ( .C (CLK), .D (new_AGEMA_signal_4198), .Q (new_AGEMA_signal_4199) ) ;
    buf_clk new_AGEMA_reg_buffer_2751 ( .C (CLK), .D (new_AGEMA_signal_4202), .Q (new_AGEMA_signal_4203) ) ;
    buf_clk new_AGEMA_reg_buffer_2755 ( .C (CLK), .D (new_AGEMA_signal_4206), .Q (new_AGEMA_signal_4207) ) ;
    buf_clk new_AGEMA_reg_buffer_2759 ( .C (CLK), .D (new_AGEMA_signal_4210), .Q (new_AGEMA_signal_4211) ) ;
    buf_clk new_AGEMA_reg_buffer_2761 ( .C (CLK), .D (new_AGEMA_signal_4212), .Q (new_AGEMA_signal_4213) ) ;
    buf_clk new_AGEMA_reg_buffer_2763 ( .C (CLK), .D (new_AGEMA_signal_4214), .Q (new_AGEMA_signal_4215) ) ;
    buf_clk new_AGEMA_reg_buffer_2773 ( .C (CLK), .D (new_AGEMA_signal_4224), .Q (new_AGEMA_signal_4225) ) ;
    buf_clk new_AGEMA_reg_buffer_2775 ( .C (CLK), .D (new_AGEMA_signal_4226), .Q (new_AGEMA_signal_4227) ) ;
    buf_clk new_AGEMA_reg_buffer_2779 ( .C (CLK), .D (new_AGEMA_signal_4230), .Q (new_AGEMA_signal_4231) ) ;
    buf_clk new_AGEMA_reg_buffer_2783 ( .C (CLK), .D (new_AGEMA_signal_4234), .Q (new_AGEMA_signal_4235) ) ;
    buf_clk new_AGEMA_reg_buffer_2785 ( .C (CLK), .D (new_AGEMA_signal_4236), .Q (new_AGEMA_signal_4237) ) ;
    buf_clk new_AGEMA_reg_buffer_2787 ( .C (CLK), .D (new_AGEMA_signal_4238), .Q (new_AGEMA_signal_4239) ) ;
    buf_clk new_AGEMA_reg_buffer_2797 ( .C (CLK), .D (new_AGEMA_signal_4248), .Q (new_AGEMA_signal_4249) ) ;
    buf_clk new_AGEMA_reg_buffer_2799 ( .C (CLK), .D (new_AGEMA_signal_4250), .Q (new_AGEMA_signal_4251) ) ;
    buf_clk new_AGEMA_reg_buffer_2803 ( .C (CLK), .D (new_AGEMA_signal_4254), .Q (new_AGEMA_signal_4255) ) ;
    buf_clk new_AGEMA_reg_buffer_2807 ( .C (CLK), .D (new_AGEMA_signal_4258), .Q (new_AGEMA_signal_4259) ) ;
    buf_clk new_AGEMA_reg_buffer_2809 ( .C (CLK), .D (new_AGEMA_signal_4260), .Q (new_AGEMA_signal_4261) ) ;
    buf_clk new_AGEMA_reg_buffer_2811 ( .C (CLK), .D (new_AGEMA_signal_4262), .Q (new_AGEMA_signal_4263) ) ;
    buf_clk new_AGEMA_reg_buffer_2813 ( .C (CLK), .D (new_AGEMA_signal_4264), .Q (new_AGEMA_signal_4265) ) ;
    buf_clk new_AGEMA_reg_buffer_2815 ( .C (CLK), .D (new_AGEMA_signal_4266), .Q (new_AGEMA_signal_4267) ) ;
    buf_clk new_AGEMA_reg_buffer_2817 ( .C (CLK), .D (new_AGEMA_signal_4268), .Q (new_AGEMA_signal_4269) ) ;
    buf_clk new_AGEMA_reg_buffer_2819 ( .C (CLK), .D (new_AGEMA_signal_4270), .Q (new_AGEMA_signal_4271) ) ;
    buf_clk new_AGEMA_reg_buffer_2821 ( .C (CLK), .D (new_AGEMA_signal_4272), .Q (new_AGEMA_signal_4273) ) ;
    buf_clk new_AGEMA_reg_buffer_2823 ( .C (CLK), .D (new_AGEMA_signal_4274), .Q (new_AGEMA_signal_4275) ) ;
    buf_clk new_AGEMA_reg_buffer_2825 ( .C (CLK), .D (new_AGEMA_signal_4276), .Q (new_AGEMA_signal_4277) ) ;
    buf_clk new_AGEMA_reg_buffer_2827 ( .C (CLK), .D (new_AGEMA_signal_4278), .Q (new_AGEMA_signal_4279) ) ;
    buf_clk new_AGEMA_reg_buffer_2829 ( .C (CLK), .D (new_AGEMA_signal_4280), .Q (new_AGEMA_signal_4281) ) ;
    buf_clk new_AGEMA_reg_buffer_2831 ( .C (CLK), .D (new_AGEMA_signal_4282), .Q (new_AGEMA_signal_4283) ) ;
    buf_clk new_AGEMA_reg_buffer_2833 ( .C (CLK), .D (new_AGEMA_signal_4284), .Q (new_AGEMA_signal_4285) ) ;
    buf_clk new_AGEMA_reg_buffer_2835 ( .C (CLK), .D (new_AGEMA_signal_4286), .Q (new_AGEMA_signal_4287) ) ;
    buf_clk new_AGEMA_reg_buffer_2837 ( .C (CLK), .D (new_AGEMA_signal_4288), .Q (new_AGEMA_signal_4289) ) ;
    buf_clk new_AGEMA_reg_buffer_2839 ( .C (CLK), .D (new_AGEMA_signal_4290), .Q (new_AGEMA_signal_4291) ) ;
    buf_clk new_AGEMA_reg_buffer_2841 ( .C (CLK), .D (new_AGEMA_signal_4292), .Q (new_AGEMA_signal_4293) ) ;
    buf_clk new_AGEMA_reg_buffer_2843 ( .C (CLK), .D (new_AGEMA_signal_4294), .Q (new_AGEMA_signal_4295) ) ;
    buf_clk new_AGEMA_reg_buffer_2845 ( .C (CLK), .D (new_AGEMA_signal_4296), .Q (new_AGEMA_signal_4297) ) ;
    buf_clk new_AGEMA_reg_buffer_2847 ( .C (CLK), .D (new_AGEMA_signal_4298), .Q (new_AGEMA_signal_4299) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (CLK), .D (new_AGEMA_signal_4300), .Q (new_AGEMA_signal_4301) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (CLK), .D (new_AGEMA_signal_4302), .Q (new_AGEMA_signal_4303) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (CLK), .D (new_AGEMA_signal_4304), .Q (new_AGEMA_signal_4305) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (CLK), .D (new_AGEMA_signal_4306), .Q (new_AGEMA_signal_4307) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (CLK), .D (new_AGEMA_signal_4308), .Q (new_AGEMA_signal_4309) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (CLK), .D (new_AGEMA_signal_4310), .Q (new_AGEMA_signal_4311) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (CLK), .D (new_AGEMA_signal_4312), .Q (new_AGEMA_signal_4313) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (CLK), .D (new_AGEMA_signal_4314), .Q (new_AGEMA_signal_4315) ) ;
    buf_clk new_AGEMA_reg_buffer_2865 ( .C (CLK), .D (new_AGEMA_signal_4316), .Q (new_AGEMA_signal_4317) ) ;
    buf_clk new_AGEMA_reg_buffer_2867 ( .C (CLK), .D (new_AGEMA_signal_4318), .Q (new_AGEMA_signal_4319) ) ;
    buf_clk new_AGEMA_reg_buffer_2869 ( .C (CLK), .D (new_AGEMA_signal_4320), .Q (new_AGEMA_signal_4321) ) ;
    buf_clk new_AGEMA_reg_buffer_2871 ( .C (CLK), .D (new_AGEMA_signal_4322), .Q (new_AGEMA_signal_4323) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (CLK), .D (new_AGEMA_signal_4324), .Q (new_AGEMA_signal_4325) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (CLK), .D (new_AGEMA_signal_4326), .Q (new_AGEMA_signal_4327) ) ;
    buf_clk new_AGEMA_reg_buffer_2879 ( .C (CLK), .D (new_AGEMA_signal_4330), .Q (new_AGEMA_signal_4331) ) ;
    buf_clk new_AGEMA_reg_buffer_2883 ( .C (CLK), .D (new_AGEMA_signal_4334), .Q (new_AGEMA_signal_4335) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (CLK), .D (new_AGEMA_signal_4338), .Q (new_AGEMA_signal_4339) ) ;
    buf_clk new_AGEMA_reg_buffer_2891 ( .C (CLK), .D (new_AGEMA_signal_4342), .Q (new_AGEMA_signal_4343) ) ;
    buf_clk new_AGEMA_reg_buffer_2895 ( .C (CLK), .D (new_AGEMA_signal_4346), .Q (new_AGEMA_signal_4347) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (CLK), .D (new_AGEMA_signal_4350), .Q (new_AGEMA_signal_4351) ) ;
    buf_clk new_AGEMA_reg_buffer_2903 ( .C (CLK), .D (new_AGEMA_signal_4354), .Q (new_AGEMA_signal_4355) ) ;
    buf_clk new_AGEMA_reg_buffer_2907 ( .C (CLK), .D (new_AGEMA_signal_4358), .Q (new_AGEMA_signal_4359) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (CLK), .D (new_AGEMA_signal_4362), .Q (new_AGEMA_signal_4363) ) ;
    buf_clk new_AGEMA_reg_buffer_2915 ( .C (CLK), .D (new_AGEMA_signal_4366), .Q (new_AGEMA_signal_4367) ) ;
    buf_clk new_AGEMA_reg_buffer_2919 ( .C (CLK), .D (new_AGEMA_signal_4370), .Q (new_AGEMA_signal_4371) ) ;

    /* register cells */
    DFF_X1 LED_128_Instance_ks_reg_0__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4331), .Q (LED_128_Instance_ks_reg_0__Q), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_1__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4335), .Q (LED_128_Instance_n26), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_2__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4339), .Q (LED_128_Instance_n25), .QN () ) ;
    DFF_X1 LED_128_Instance_ks_reg_3__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4343), .Q (LED_128_Instance_n2), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_0__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4347), .Q (roundconstant[0]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_1__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4351), .Q (roundconstant[1]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_2__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4355), .Q (roundconstant[2]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_3__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4359), .Q (roundconstant[3]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_4__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4363), .Q (roundconstant[4]), .QN () ) ;
    DFF_X1 LED_128_Instance_roundconstant_reg_5__FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4367), .Q (roundconstant[5]), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_0__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2201, LED_128_Instance_state1[0]}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_1__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2319, LED_128_Instance_state1[1]}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_2__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2227, LED_128_Instance_state1[2]}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_3__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2277, LED_128_Instance_state1[3]}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_4__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2229, LED_128_Instance_state1[4]}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_5__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2321, LED_128_Instance_state1[5]}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_6__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2231, LED_128_Instance_state1[6]}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_7__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2233, LED_128_Instance_state1[7]}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_8__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2235, LED_128_Instance_state1[8]}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_9__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2279, LED_128_Instance_state1[9]}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_10__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2237, LED_128_Instance_state1[10]}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_11__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2239, LED_128_Instance_state1[11]}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_12__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2241, LED_128_Instance_state1[12]}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_13__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2281, LED_128_Instance_state1[13]}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_14__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2243, LED_128_Instance_state1[14]}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_15__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2283, LED_128_Instance_state1[15]}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_16__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2368, LED_128_Instance_state1[16]}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_17__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2403, LED_128_Instance_state1[17]}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_18__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2405, LED_128_Instance_state1[18]}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_19__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2323, LED_128_Instance_state1[19]}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_20__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2325, LED_128_Instance_state1[20]}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_21__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2370, LED_128_Instance_state1[21]}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_22__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2407, LED_128_Instance_state1[22]}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_23__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2327, LED_128_Instance_state1[23]}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_24__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2329, LED_128_Instance_state1[24]}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_25__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2372, LED_128_Instance_state1[25]}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_26__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2374, LED_128_Instance_state1[26]}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_27__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2331, LED_128_Instance_state1[27]}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_28__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2376, LED_128_Instance_state1[28]}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_29__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2409, LED_128_Instance_state1[29]}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_30__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2378, LED_128_Instance_state1[30]}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_31__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2333, LED_128_Instance_state1[31]}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_32__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2411, LED_128_Instance_state1[32]}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_33__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2443, LED_128_Instance_state1[33]}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_34__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2413, LED_128_Instance_state1[34]}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_35__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2463, LED_128_Instance_state1[35]}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_36__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2415, LED_128_Instance_state1[36]}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_37__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2417, LED_128_Instance_state1[37]}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_38__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2380, LED_128_Instance_state1[38]}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_39__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2465, LED_128_Instance_state1[39]}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_40__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2419, LED_128_Instance_state1[40]}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_41__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2421, LED_128_Instance_state1[41]}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_42__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2382, LED_128_Instance_state1[42]}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_43__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2445, LED_128_Instance_state1[43]}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_44__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2423, LED_128_Instance_state1[44]}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_45__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2447, LED_128_Instance_state1[45]}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_46__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2425, LED_128_Instance_state1[46]}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_47__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2449, LED_128_Instance_state1[47]}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_48__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2505, LED_128_Instance_state1[48]}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_49__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2513, LED_128_Instance_state1[49]}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_50__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2467, LED_128_Instance_state1[50]}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_51__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2469, LED_128_Instance_state1[51]}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_52__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2507, LED_128_Instance_state1[52]}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_53__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2515, LED_128_Instance_state1[53]}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_54__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2451, LED_128_Instance_state1[54]}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_55__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2471, LED_128_Instance_state1[55]}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_56__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2497, LED_128_Instance_state1[56]}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_57__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2509, LED_128_Instance_state1[57]}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_58__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2453, LED_128_Instance_state1[58]}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_59__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2455, LED_128_Instance_state1[59]}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_60__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2499, LED_128_Instance_state1[60]}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_61__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2511, LED_128_Instance_state1[61]}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_62__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2473, LED_128_Instance_state1[62]}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) LED_128_Instance_cipherstate_reg_63__FF_FF ( .clk (CLK), .D ({new_AGEMA_signal_2475, LED_128_Instance_state1[63]}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 internal_done_reg_FF_FF ( .CK (CLK), .D (new_AGEMA_signal_4371), .Q (OUT_done), .QN () ) ;
endmodule
