/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [203:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_555 ;
    wire signal_556 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_560 ;
    wire signal_561 ;
    wire signal_562 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_569 ;
    wire signal_570 ;
    wire signal_571 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_136 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_283, signal_282, signal_281, signal_151}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_137 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_289, signal_288, signal_287, signal_152}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_138 ( .a ({X_s3[7], X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_295, signal_294, signal_293, signal_153}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_139 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_298, signal_297, signal_296, signal_154}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_140 ( .a ({X_s3[3], X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_304, signal_303, signal_302, signal_155}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_141 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_313, signal_312, signal_311, signal_156}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_142 ( .a ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_316, signal_315, signal_314, signal_157}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_143 ( .a ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s3[2], X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_319, signal_318, signal_317, signal_158}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_144 ( .a ({X_s3[4], X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_325, signal_324, signal_323, signal_159}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_145 ( .a ({X_s3[1], X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_328, signal_327, signal_326, signal_160}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_146 ( .a ({signal_283, signal_282, signal_281, signal_151}), .b ({signal_304, signal_303, signal_302, signal_155}), .c ({signal_331, signal_330, signal_329, signal_161}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_147 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_313, signal_312, signal_311, signal_156}), .c ({signal_334, signal_333, signal_332, signal_162}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_148 ( .a ({signal_295, signal_294, signal_293, signal_153}), .b ({signal_298, signal_297, signal_296, signal_154}), .c ({signal_337, signal_336, signal_335, signal_163}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_149 ( .a ({signal_304, signal_303, signal_302, signal_155}), .b ({signal_316, signal_315, signal_314, signal_157}), .c ({signal_340, signal_339, signal_338, signal_164}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_150 ( .a ({signal_304, signal_303, signal_302, signal_155}), .b ({signal_319, signal_318, signal_317, signal_158}), .c ({signal_343, signal_342, signal_341, signal_165}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_151 ( .a ({signal_313, signal_312, signal_311, signal_156}), .b ({signal_325, signal_324, signal_323, signal_159}), .c ({signal_346, signal_345, signal_344, signal_166}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_152 ( .a ({signal_313, signal_312, signal_311, signal_156}), .b ({signal_328, signal_327, signal_326, signal_160}), .c ({signal_349, signal_348, signal_347, signal_167}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_153 ( .a ({signal_283, signal_282, signal_281, signal_151}), .b ({signal_319, signal_318, signal_317, signal_158}), .c ({signal_352, signal_351, signal_350, signal_168}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_160 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_331, signal_330, signal_329, signal_161}), .c ({signal_373, signal_372, signal_371, signal_175}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_161 ( .a ({signal_313, signal_312, signal_311, signal_156}), .b ({signal_331, signal_330, signal_329, signal_161}), .c ({signal_376, signal_375, signal_374, signal_176}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_162 ( .a ({signal_316, signal_315, signal_314, signal_157}), .b ({signal_331, signal_330, signal_329, signal_161}), .c ({signal_379, signal_378, signal_377, signal_177}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_163 ( .a ({signal_334, signal_333, signal_332, signal_162}), .b ({signal_343, signal_342, signal_341, signal_165}), .c ({signal_382, signal_381, signal_380, signal_178}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_164 ( .a ({signal_283, signal_282, signal_281, signal_151}), .b ({signal_346, signal_345, signal_344, signal_166}), .c ({signal_385, signal_384, signal_383, signal_179}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_165 ( .a ({signal_289, signal_288, signal_287, signal_152}), .b ({signal_349, signal_348, signal_347, signal_167}), .c ({signal_388, signal_387, signal_386, signal_180}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_166 ( .a ({signal_295, signal_294, signal_293, signal_153}), .b ({signal_343, signal_342, signal_341, signal_165}), .c ({signal_391, signal_390, signal_389, signal_181}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_170 ( .a ({signal_289, signal_288, signal_287, signal_152}), .b ({signal_376, signal_375, signal_374, signal_176}), .c ({signal_403, signal_402, signal_401, signal_185}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_171 ( .a ({signal_382, signal_381, signal_380, signal_178}), .b ({signal_385, signal_384, signal_383, signal_179}), .c ({signal_406, signal_405, signal_404, signal_186}) ) ;

    /* cells in depth 1 */
    buf_clk cell_268 ( .C (clk), .D (signal_177), .Q (signal_923) ) ;
    buf_clk cell_270 ( .C (clk), .D (signal_377), .Q (signal_925) ) ;
    buf_clk cell_272 ( .C (clk), .D (signal_378), .Q (signal_927) ) ;
    buf_clk cell_274 ( .C (clk), .D (signal_379), .Q (signal_929) ) ;
    buf_clk cell_276 ( .C (clk), .D (signal_181), .Q (signal_931) ) ;
    buf_clk cell_278 ( .C (clk), .D (signal_389), .Q (signal_933) ) ;
    buf_clk cell_280 ( .C (clk), .D (signal_390), .Q (signal_935) ) ;
    buf_clk cell_282 ( .C (clk), .D (signal_391), .Q (signal_937) ) ;
    buf_clk cell_284 ( .C (clk), .D (signal_185), .Q (signal_939) ) ;
    buf_clk cell_286 ( .C (clk), .D (signal_401), .Q (signal_941) ) ;
    buf_clk cell_288 ( .C (clk), .D (signal_402), .Q (signal_943) ) ;
    buf_clk cell_290 ( .C (clk), .D (signal_403), .Q (signal_945) ) ;
    buf_clk cell_292 ( .C (clk), .D (signal_186), .Q (signal_947) ) ;
    buf_clk cell_294 ( .C (clk), .D (signal_404), .Q (signal_949) ) ;
    buf_clk cell_296 ( .C (clk), .D (signal_405), .Q (signal_951) ) ;
    buf_clk cell_298 ( .C (clk), .D (signal_406), .Q (signal_953) ) ;
    buf_clk cell_364 ( .C (clk), .D (signal_175), .Q (signal_1019) ) ;
    buf_clk cell_370 ( .C (clk), .D (signal_371), .Q (signal_1025) ) ;
    buf_clk cell_376 ( .C (clk), .D (signal_372), .Q (signal_1031) ) ;
    buf_clk cell_382 ( .C (clk), .D (signal_373), .Q (signal_1037) ) ;
    buf_clk cell_388 ( .C (clk), .D (X_s0[0]), .Q (signal_1043) ) ;
    buf_clk cell_394 ( .C (clk), .D (X_s1[0]), .Q (signal_1049) ) ;
    buf_clk cell_400 ( .C (clk), .D (X_s2[0]), .Q (signal_1055) ) ;
    buf_clk cell_406 ( .C (clk), .D (X_s3[0]), .Q (signal_1061) ) ;
    buf_clk cell_412 ( .C (clk), .D (signal_162), .Q (signal_1067) ) ;
    buf_clk cell_418 ( .C (clk), .D (signal_332), .Q (signal_1073) ) ;
    buf_clk cell_424 ( .C (clk), .D (signal_333), .Q (signal_1079) ) ;
    buf_clk cell_430 ( .C (clk), .D (signal_334), .Q (signal_1085) ) ;
    buf_clk cell_436 ( .C (clk), .D (signal_178), .Q (signal_1091) ) ;
    buf_clk cell_442 ( .C (clk), .D (signal_380), .Q (signal_1097) ) ;
    buf_clk cell_448 ( .C (clk), .D (signal_381), .Q (signal_1103) ) ;
    buf_clk cell_454 ( .C (clk), .D (signal_382), .Q (signal_1109) ) ;
    buf_clk cell_460 ( .C (clk), .D (signal_180), .Q (signal_1115) ) ;
    buf_clk cell_466 ( .C (clk), .D (signal_386), .Q (signal_1121) ) ;
    buf_clk cell_472 ( .C (clk), .D (signal_387), .Q (signal_1127) ) ;
    buf_clk cell_478 ( .C (clk), .D (signal_388), .Q (signal_1133) ) ;
    buf_clk cell_484 ( .C (clk), .D (signal_166), .Q (signal_1139) ) ;
    buf_clk cell_490 ( .C (clk), .D (signal_344), .Q (signal_1145) ) ;
    buf_clk cell_496 ( .C (clk), .D (signal_345), .Q (signal_1151) ) ;
    buf_clk cell_502 ( .C (clk), .D (signal_346), .Q (signal_1157) ) ;
    buf_clk cell_508 ( .C (clk), .D (signal_167), .Q (signal_1163) ) ;
    buf_clk cell_514 ( .C (clk), .D (signal_347), .Q (signal_1169) ) ;
    buf_clk cell_520 ( .C (clk), .D (signal_348), .Q (signal_1175) ) ;
    buf_clk cell_526 ( .C (clk), .D (signal_349), .Q (signal_1181) ) ;
    buf_clk cell_532 ( .C (clk), .D (signal_179), .Q (signal_1187) ) ;
    buf_clk cell_538 ( .C (clk), .D (signal_383), .Q (signal_1193) ) ;
    buf_clk cell_544 ( .C (clk), .D (signal_384), .Q (signal_1199) ) ;
    buf_clk cell_550 ( .C (clk), .D (signal_385), .Q (signal_1205) ) ;
    buf_clk cell_556 ( .C (clk), .D (signal_161), .Q (signal_1211) ) ;
    buf_clk cell_562 ( .C (clk), .D (signal_329), .Q (signal_1217) ) ;
    buf_clk cell_568 ( .C (clk), .D (signal_330), .Q (signal_1223) ) ;
    buf_clk cell_574 ( .C (clk), .D (signal_331), .Q (signal_1229) ) ;
    buf_clk cell_580 ( .C (clk), .D (signal_165), .Q (signal_1235) ) ;
    buf_clk cell_586 ( .C (clk), .D (signal_341), .Q (signal_1241) ) ;
    buf_clk cell_592 ( .C (clk), .D (signal_342), .Q (signal_1247) ) ;
    buf_clk cell_598 ( .C (clk), .D (signal_343), .Q (signal_1253) ) ;
    buf_clk cell_604 ( .C (clk), .D (signal_164), .Q (signal_1259) ) ;
    buf_clk cell_610 ( .C (clk), .D (signal_338), .Q (signal_1265) ) ;
    buf_clk cell_616 ( .C (clk), .D (signal_339), .Q (signal_1271) ) ;
    buf_clk cell_622 ( .C (clk), .D (signal_340), .Q (signal_1277) ) ;
    buf_clk cell_628 ( .C (clk), .D (signal_176), .Q (signal_1283) ) ;
    buf_clk cell_634 ( .C (clk), .D (signal_374), .Q (signal_1289) ) ;
    buf_clk cell_640 ( .C (clk), .D (signal_375), .Q (signal_1295) ) ;
    buf_clk cell_646 ( .C (clk), .D (signal_376), .Q (signal_1301) ) ;
    buf_clk cell_652 ( .C (clk), .D (signal_163), .Q (signal_1307) ) ;
    buf_clk cell_658 ( .C (clk), .D (signal_335), .Q (signal_1313) ) ;
    buf_clk cell_664 ( .C (clk), .D (signal_336), .Q (signal_1319) ) ;
    buf_clk cell_670 ( .C (clk), .D (signal_337), .Q (signal_1325) ) ;
    buf_clk cell_676 ( .C (clk), .D (signal_153), .Q (signal_1331) ) ;
    buf_clk cell_682 ( .C (clk), .D (signal_293), .Q (signal_1337) ) ;
    buf_clk cell_688 ( .C (clk), .D (signal_294), .Q (signal_1343) ) ;
    buf_clk cell_694 ( .C (clk), .D (signal_295), .Q (signal_1349) ) ;
    buf_clk cell_700 ( .C (clk), .D (signal_151), .Q (signal_1355) ) ;
    buf_clk cell_706 ( .C (clk), .D (signal_281), .Q (signal_1361) ) ;
    buf_clk cell_712 ( .C (clk), .D (signal_282), .Q (signal_1367) ) ;
    buf_clk cell_718 ( .C (clk), .D (signal_283), .Q (signal_1373) ) ;
    buf_clk cell_724 ( .C (clk), .D (signal_152), .Q (signal_1379) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_287), .Q (signal_1385) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_288), .Q (signal_1391) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_289), .Q (signal_1397) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_168), .Q (signal_1403) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_350), .Q (signal_1409) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_351), .Q (signal_1415) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_352), .Q (signal_1421) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_154), .Q (signal_1427) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_296), .Q (signal_1433) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_297), .Q (signal_1439) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_298), .Q (signal_1445) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_154 ( .a ({signal_331, signal_330, signal_329, signal_161}), .b ({signal_337, signal_336, signal_335, signal_163}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_355, signal_354, signal_353, signal_169}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_155 ( .a ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_346, signal_345, signal_344, signal_166}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_358, signal_357, signal_356, signal_170}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_156 ( .a ({signal_295, signal_294, signal_293, signal_153}), .b ({signal_343, signal_342, signal_341, signal_165}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_361, signal_360, signal_359, signal_171}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_157 ( .a ({signal_334, signal_333, signal_332, signal_162}), .b ({signal_349, signal_348, signal_347, signal_167}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_364, signal_363, signal_362, signal_172}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_158 ( .a ({signal_283, signal_282, signal_281, signal_151}), .b ({signal_340, signal_339, signal_338, signal_164}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_367, signal_366, signal_365, signal_173}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_159 ( .a ({signal_298, signal_297, signal_296, signal_154}), .b ({signal_352, signal_351, signal_350, signal_168}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_370, signal_369, signal_368, signal_174}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_167 ( .a ({signal_373, signal_372, signal_371, signal_175}), .b ({signal_388, signal_387, signal_386, signal_180}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_394, signal_393, signal_392, signal_182}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_168 ( .a ({signal_382, signal_381, signal_380, signal_178}), .b ({signal_385, signal_384, signal_383, signal_179}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_397, signal_396, signal_395, signal_183}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_169 ( .a ({signal_289, signal_288, signal_287, signal_152}), .b ({signal_376, signal_375, signal_374, signal_176}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_400, signal_399, signal_398, signal_184}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_172 ( .a ({signal_930, signal_928, signal_926, signal_924}), .b ({signal_355, signal_354, signal_353, signal_169}), .c ({signal_409, signal_408, signal_407, signal_187}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_173 ( .a ({signal_355, signal_354, signal_353, signal_169}), .b ({signal_358, signal_357, signal_356, signal_170}), .c ({signal_412, signal_411, signal_410, signal_188}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_174 ( .a ({signal_938, signal_936, signal_934, signal_932}), .b ({signal_361, signal_360, signal_359, signal_171}), .c ({signal_415, signal_414, signal_413, signal_189}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_175 ( .a ({signal_367, signal_366, signal_365, signal_173}), .b ({signal_370, signal_369, signal_368, signal_174}), .c ({signal_418, signal_417, signal_416, signal_190}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_176 ( .a ({signal_361, signal_360, signal_359, signal_171}), .b ({signal_397, signal_396, signal_395, signal_183}), .c ({signal_421, signal_420, signal_419, signal_191}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_177 ( .a ({signal_367, signal_366, signal_365, signal_173}), .b ({signal_400, signal_399, signal_398, signal_184}), .c ({signal_424, signal_423, signal_422, signal_192}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_178 ( .a ({signal_394, signal_393, signal_392, signal_182}), .b ({signal_409, signal_408, signal_407, signal_187}), .c ({signal_427, signal_426, signal_425, signal_193}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_179 ( .a ({signal_946, signal_944, signal_942, signal_940}), .b ({signal_412, signal_411, signal_410, signal_188}), .c ({signal_430, signal_429, signal_428, signal_194}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_180 ( .a ({signal_364, signal_363, signal_362, signal_172}), .b ({signal_415, signal_414, signal_413, signal_189}), .c ({signal_433, signal_432, signal_431, signal_195}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_181 ( .a ({signal_421, signal_420, signal_419, signal_191}), .b ({signal_424, signal_423, signal_422, signal_192}), .c ({signal_436, signal_435, signal_434, signal_196}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_182 ( .a ({signal_418, signal_417, signal_416, signal_190}), .b ({signal_427, signal_426, signal_425, signal_193}), .c ({signal_439, signal_438, signal_437, signal_197}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_183 ( .a ({signal_424, signal_423, signal_422, signal_192}), .b ({signal_430, signal_429, signal_428, signal_194}), .c ({signal_442, signal_441, signal_440, signal_198}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_184 ( .a ({signal_418, signal_417, signal_416, signal_190}), .b ({signal_433, signal_432, signal_431, signal_195}), .c ({signal_445, signal_444, signal_443, signal_199}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_187 ( .a ({signal_954, signal_952, signal_950, signal_948}), .b ({signal_436, signal_435, signal_434, signal_196}), .c ({signal_454, signal_453, signal_452, signal_202}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_188 ( .a ({signal_439, signal_438, signal_437, signal_197}), .b ({signal_442, signal_441, signal_440, signal_198}), .c ({signal_457, signal_456, signal_455, signal_203}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_190 ( .a ({signal_445, signal_444, signal_443, signal_199}), .b ({signal_454, signal_453, signal_452, signal_202}), .c ({signal_463, signal_462, signal_461, signal_205}) ) ;
    buf_clk cell_269 ( .C (clk), .D (signal_923), .Q (signal_924) ) ;
    buf_clk cell_271 ( .C (clk), .D (signal_925), .Q (signal_926) ) ;
    buf_clk cell_273 ( .C (clk), .D (signal_927), .Q (signal_928) ) ;
    buf_clk cell_275 ( .C (clk), .D (signal_929), .Q (signal_930) ) ;
    buf_clk cell_277 ( .C (clk), .D (signal_931), .Q (signal_932) ) ;
    buf_clk cell_279 ( .C (clk), .D (signal_933), .Q (signal_934) ) ;
    buf_clk cell_281 ( .C (clk), .D (signal_935), .Q (signal_936) ) ;
    buf_clk cell_283 ( .C (clk), .D (signal_937), .Q (signal_938) ) ;
    buf_clk cell_285 ( .C (clk), .D (signal_939), .Q (signal_940) ) ;
    buf_clk cell_287 ( .C (clk), .D (signal_941), .Q (signal_942) ) ;
    buf_clk cell_289 ( .C (clk), .D (signal_943), .Q (signal_944) ) ;
    buf_clk cell_291 ( .C (clk), .D (signal_945), .Q (signal_946) ) ;
    buf_clk cell_293 ( .C (clk), .D (signal_947), .Q (signal_948) ) ;
    buf_clk cell_295 ( .C (clk), .D (signal_949), .Q (signal_950) ) ;
    buf_clk cell_297 ( .C (clk), .D (signal_951), .Q (signal_952) ) ;
    buf_clk cell_299 ( .C (clk), .D (signal_953), .Q (signal_954) ) ;
    buf_clk cell_365 ( .C (clk), .D (signal_1019), .Q (signal_1020) ) ;
    buf_clk cell_371 ( .C (clk), .D (signal_1025), .Q (signal_1026) ) ;
    buf_clk cell_377 ( .C (clk), .D (signal_1031), .Q (signal_1032) ) ;
    buf_clk cell_383 ( .C (clk), .D (signal_1037), .Q (signal_1038) ) ;
    buf_clk cell_389 ( .C (clk), .D (signal_1043), .Q (signal_1044) ) ;
    buf_clk cell_395 ( .C (clk), .D (signal_1049), .Q (signal_1050) ) ;
    buf_clk cell_401 ( .C (clk), .D (signal_1055), .Q (signal_1056) ) ;
    buf_clk cell_407 ( .C (clk), .D (signal_1061), .Q (signal_1062) ) ;
    buf_clk cell_413 ( .C (clk), .D (signal_1067), .Q (signal_1068) ) ;
    buf_clk cell_419 ( .C (clk), .D (signal_1073), .Q (signal_1074) ) ;
    buf_clk cell_425 ( .C (clk), .D (signal_1079), .Q (signal_1080) ) ;
    buf_clk cell_431 ( .C (clk), .D (signal_1085), .Q (signal_1086) ) ;
    buf_clk cell_437 ( .C (clk), .D (signal_1091), .Q (signal_1092) ) ;
    buf_clk cell_443 ( .C (clk), .D (signal_1097), .Q (signal_1098) ) ;
    buf_clk cell_449 ( .C (clk), .D (signal_1103), .Q (signal_1104) ) ;
    buf_clk cell_455 ( .C (clk), .D (signal_1109), .Q (signal_1110) ) ;
    buf_clk cell_461 ( .C (clk), .D (signal_1115), .Q (signal_1116) ) ;
    buf_clk cell_467 ( .C (clk), .D (signal_1121), .Q (signal_1122) ) ;
    buf_clk cell_473 ( .C (clk), .D (signal_1127), .Q (signal_1128) ) ;
    buf_clk cell_479 ( .C (clk), .D (signal_1133), .Q (signal_1134) ) ;
    buf_clk cell_485 ( .C (clk), .D (signal_1139), .Q (signal_1140) ) ;
    buf_clk cell_491 ( .C (clk), .D (signal_1145), .Q (signal_1146) ) ;
    buf_clk cell_497 ( .C (clk), .D (signal_1151), .Q (signal_1152) ) ;
    buf_clk cell_503 ( .C (clk), .D (signal_1157), .Q (signal_1158) ) ;
    buf_clk cell_509 ( .C (clk), .D (signal_1163), .Q (signal_1164) ) ;
    buf_clk cell_515 ( .C (clk), .D (signal_1169), .Q (signal_1170) ) ;
    buf_clk cell_521 ( .C (clk), .D (signal_1175), .Q (signal_1176) ) ;
    buf_clk cell_527 ( .C (clk), .D (signal_1181), .Q (signal_1182) ) ;
    buf_clk cell_533 ( .C (clk), .D (signal_1187), .Q (signal_1188) ) ;
    buf_clk cell_539 ( .C (clk), .D (signal_1193), .Q (signal_1194) ) ;
    buf_clk cell_545 ( .C (clk), .D (signal_1199), .Q (signal_1200) ) ;
    buf_clk cell_551 ( .C (clk), .D (signal_1205), .Q (signal_1206) ) ;
    buf_clk cell_557 ( .C (clk), .D (signal_1211), .Q (signal_1212) ) ;
    buf_clk cell_563 ( .C (clk), .D (signal_1217), .Q (signal_1218) ) ;
    buf_clk cell_569 ( .C (clk), .D (signal_1223), .Q (signal_1224) ) ;
    buf_clk cell_575 ( .C (clk), .D (signal_1229), .Q (signal_1230) ) ;
    buf_clk cell_581 ( .C (clk), .D (signal_1235), .Q (signal_1236) ) ;
    buf_clk cell_587 ( .C (clk), .D (signal_1241), .Q (signal_1242) ) ;
    buf_clk cell_593 ( .C (clk), .D (signal_1247), .Q (signal_1248) ) ;
    buf_clk cell_599 ( .C (clk), .D (signal_1253), .Q (signal_1254) ) ;
    buf_clk cell_605 ( .C (clk), .D (signal_1259), .Q (signal_1260) ) ;
    buf_clk cell_611 ( .C (clk), .D (signal_1265), .Q (signal_1266) ) ;
    buf_clk cell_617 ( .C (clk), .D (signal_1271), .Q (signal_1272) ) ;
    buf_clk cell_623 ( .C (clk), .D (signal_1277), .Q (signal_1278) ) ;
    buf_clk cell_629 ( .C (clk), .D (signal_1283), .Q (signal_1284) ) ;
    buf_clk cell_635 ( .C (clk), .D (signal_1289), .Q (signal_1290) ) ;
    buf_clk cell_641 ( .C (clk), .D (signal_1295), .Q (signal_1296) ) ;
    buf_clk cell_647 ( .C (clk), .D (signal_1301), .Q (signal_1302) ) ;
    buf_clk cell_653 ( .C (clk), .D (signal_1307), .Q (signal_1308) ) ;
    buf_clk cell_659 ( .C (clk), .D (signal_1313), .Q (signal_1314) ) ;
    buf_clk cell_665 ( .C (clk), .D (signal_1319), .Q (signal_1320) ) ;
    buf_clk cell_671 ( .C (clk), .D (signal_1325), .Q (signal_1326) ) ;
    buf_clk cell_677 ( .C (clk), .D (signal_1331), .Q (signal_1332) ) ;
    buf_clk cell_683 ( .C (clk), .D (signal_1337), .Q (signal_1338) ) ;
    buf_clk cell_689 ( .C (clk), .D (signal_1343), .Q (signal_1344) ) ;
    buf_clk cell_695 ( .C (clk), .D (signal_1349), .Q (signal_1350) ) ;
    buf_clk cell_701 ( .C (clk), .D (signal_1355), .Q (signal_1356) ) ;
    buf_clk cell_707 ( .C (clk), .D (signal_1361), .Q (signal_1362) ) ;
    buf_clk cell_713 ( .C (clk), .D (signal_1367), .Q (signal_1368) ) ;
    buf_clk cell_719 ( .C (clk), .D (signal_1373), .Q (signal_1374) ) ;
    buf_clk cell_725 ( .C (clk), .D (signal_1379), .Q (signal_1380) ) ;
    buf_clk cell_731 ( .C (clk), .D (signal_1385), .Q (signal_1386) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_1391), .Q (signal_1392) ) ;
    buf_clk cell_743 ( .C (clk), .D (signal_1397), .Q (signal_1398) ) ;
    buf_clk cell_749 ( .C (clk), .D (signal_1403), .Q (signal_1404) ) ;
    buf_clk cell_755 ( .C (clk), .D (signal_1409), .Q (signal_1410) ) ;
    buf_clk cell_761 ( .C (clk), .D (signal_1415), .Q (signal_1416) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_1421), .Q (signal_1422) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_1427), .Q (signal_1428) ) ;
    buf_clk cell_779 ( .C (clk), .D (signal_1433), .Q (signal_1434) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_1439), .Q (signal_1440) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_1445), .Q (signal_1446) ) ;

    /* cells in depth 3 */
    buf_clk cell_300 ( .C (clk), .D (signal_198), .Q (signal_955) ) ;
    buf_clk cell_302 ( .C (clk), .D (signal_440), .Q (signal_957) ) ;
    buf_clk cell_304 ( .C (clk), .D (signal_441), .Q (signal_959) ) ;
    buf_clk cell_306 ( .C (clk), .D (signal_442), .Q (signal_961) ) ;
    buf_clk cell_308 ( .C (clk), .D (signal_202), .Q (signal_963) ) ;
    buf_clk cell_310 ( .C (clk), .D (signal_452), .Q (signal_965) ) ;
    buf_clk cell_312 ( .C (clk), .D (signal_453), .Q (signal_967) ) ;
    buf_clk cell_314 ( .C (clk), .D (signal_454), .Q (signal_969) ) ;
    buf_clk cell_316 ( .C (clk), .D (signal_203), .Q (signal_971) ) ;
    buf_clk cell_318 ( .C (clk), .D (signal_455), .Q (signal_973) ) ;
    buf_clk cell_320 ( .C (clk), .D (signal_456), .Q (signal_975) ) ;
    buf_clk cell_322 ( .C (clk), .D (signal_457), .Q (signal_977) ) ;
    buf_clk cell_324 ( .C (clk), .D (signal_205), .Q (signal_979) ) ;
    buf_clk cell_326 ( .C (clk), .D (signal_461), .Q (signal_981) ) ;
    buf_clk cell_328 ( .C (clk), .D (signal_462), .Q (signal_983) ) ;
    buf_clk cell_330 ( .C (clk), .D (signal_463), .Q (signal_985) ) ;
    buf_clk cell_366 ( .C (clk), .D (signal_1020), .Q (signal_1021) ) ;
    buf_clk cell_372 ( .C (clk), .D (signal_1026), .Q (signal_1027) ) ;
    buf_clk cell_378 ( .C (clk), .D (signal_1032), .Q (signal_1033) ) ;
    buf_clk cell_384 ( .C (clk), .D (signal_1038), .Q (signal_1039) ) ;
    buf_clk cell_390 ( .C (clk), .D (signal_1044), .Q (signal_1045) ) ;
    buf_clk cell_396 ( .C (clk), .D (signal_1050), .Q (signal_1051) ) ;
    buf_clk cell_402 ( .C (clk), .D (signal_1056), .Q (signal_1057) ) ;
    buf_clk cell_408 ( .C (clk), .D (signal_1062), .Q (signal_1063) ) ;
    buf_clk cell_414 ( .C (clk), .D (signal_1068), .Q (signal_1069) ) ;
    buf_clk cell_420 ( .C (clk), .D (signal_1074), .Q (signal_1075) ) ;
    buf_clk cell_426 ( .C (clk), .D (signal_1080), .Q (signal_1081) ) ;
    buf_clk cell_432 ( .C (clk), .D (signal_1086), .Q (signal_1087) ) ;
    buf_clk cell_438 ( .C (clk), .D (signal_1092), .Q (signal_1093) ) ;
    buf_clk cell_444 ( .C (clk), .D (signal_1098), .Q (signal_1099) ) ;
    buf_clk cell_450 ( .C (clk), .D (signal_1104), .Q (signal_1105) ) ;
    buf_clk cell_456 ( .C (clk), .D (signal_1110), .Q (signal_1111) ) ;
    buf_clk cell_462 ( .C (clk), .D (signal_1116), .Q (signal_1117) ) ;
    buf_clk cell_468 ( .C (clk), .D (signal_1122), .Q (signal_1123) ) ;
    buf_clk cell_474 ( .C (clk), .D (signal_1128), .Q (signal_1129) ) ;
    buf_clk cell_480 ( .C (clk), .D (signal_1134), .Q (signal_1135) ) ;
    buf_clk cell_486 ( .C (clk), .D (signal_1140), .Q (signal_1141) ) ;
    buf_clk cell_492 ( .C (clk), .D (signal_1146), .Q (signal_1147) ) ;
    buf_clk cell_498 ( .C (clk), .D (signal_1152), .Q (signal_1153) ) ;
    buf_clk cell_504 ( .C (clk), .D (signal_1158), .Q (signal_1159) ) ;
    buf_clk cell_510 ( .C (clk), .D (signal_1164), .Q (signal_1165) ) ;
    buf_clk cell_516 ( .C (clk), .D (signal_1170), .Q (signal_1171) ) ;
    buf_clk cell_522 ( .C (clk), .D (signal_1176), .Q (signal_1177) ) ;
    buf_clk cell_528 ( .C (clk), .D (signal_1182), .Q (signal_1183) ) ;
    buf_clk cell_534 ( .C (clk), .D (signal_1188), .Q (signal_1189) ) ;
    buf_clk cell_540 ( .C (clk), .D (signal_1194), .Q (signal_1195) ) ;
    buf_clk cell_546 ( .C (clk), .D (signal_1200), .Q (signal_1201) ) ;
    buf_clk cell_552 ( .C (clk), .D (signal_1206), .Q (signal_1207) ) ;
    buf_clk cell_558 ( .C (clk), .D (signal_1212), .Q (signal_1213) ) ;
    buf_clk cell_564 ( .C (clk), .D (signal_1218), .Q (signal_1219) ) ;
    buf_clk cell_570 ( .C (clk), .D (signal_1224), .Q (signal_1225) ) ;
    buf_clk cell_576 ( .C (clk), .D (signal_1230), .Q (signal_1231) ) ;
    buf_clk cell_582 ( .C (clk), .D (signal_1236), .Q (signal_1237) ) ;
    buf_clk cell_588 ( .C (clk), .D (signal_1242), .Q (signal_1243) ) ;
    buf_clk cell_594 ( .C (clk), .D (signal_1248), .Q (signal_1249) ) ;
    buf_clk cell_600 ( .C (clk), .D (signal_1254), .Q (signal_1255) ) ;
    buf_clk cell_606 ( .C (clk), .D (signal_1260), .Q (signal_1261) ) ;
    buf_clk cell_612 ( .C (clk), .D (signal_1266), .Q (signal_1267) ) ;
    buf_clk cell_618 ( .C (clk), .D (signal_1272), .Q (signal_1273) ) ;
    buf_clk cell_624 ( .C (clk), .D (signal_1278), .Q (signal_1279) ) ;
    buf_clk cell_630 ( .C (clk), .D (signal_1284), .Q (signal_1285) ) ;
    buf_clk cell_636 ( .C (clk), .D (signal_1290), .Q (signal_1291) ) ;
    buf_clk cell_642 ( .C (clk), .D (signal_1296), .Q (signal_1297) ) ;
    buf_clk cell_648 ( .C (clk), .D (signal_1302), .Q (signal_1303) ) ;
    buf_clk cell_654 ( .C (clk), .D (signal_1308), .Q (signal_1309) ) ;
    buf_clk cell_660 ( .C (clk), .D (signal_1314), .Q (signal_1315) ) ;
    buf_clk cell_666 ( .C (clk), .D (signal_1320), .Q (signal_1321) ) ;
    buf_clk cell_672 ( .C (clk), .D (signal_1326), .Q (signal_1327) ) ;
    buf_clk cell_678 ( .C (clk), .D (signal_1332), .Q (signal_1333) ) ;
    buf_clk cell_684 ( .C (clk), .D (signal_1338), .Q (signal_1339) ) ;
    buf_clk cell_690 ( .C (clk), .D (signal_1344), .Q (signal_1345) ) ;
    buf_clk cell_696 ( .C (clk), .D (signal_1350), .Q (signal_1351) ) ;
    buf_clk cell_702 ( .C (clk), .D (signal_1356), .Q (signal_1357) ) ;
    buf_clk cell_708 ( .C (clk), .D (signal_1362), .Q (signal_1363) ) ;
    buf_clk cell_714 ( .C (clk), .D (signal_1368), .Q (signal_1369) ) ;
    buf_clk cell_720 ( .C (clk), .D (signal_1374), .Q (signal_1375) ) ;
    buf_clk cell_726 ( .C (clk), .D (signal_1380), .Q (signal_1381) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_1386), .Q (signal_1387) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_1392), .Q (signal_1393) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_1398), .Q (signal_1399) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_1404), .Q (signal_1405) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_1410), .Q (signal_1411) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_1416), .Q (signal_1417) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_1422), .Q (signal_1423) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_1428), .Q (signal_1429) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_1434), .Q (signal_1435) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_1440), .Q (signal_1441) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_1446), .Q (signal_1447) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_185 ( .a ({signal_439, signal_438, signal_437, signal_197}), .b ({signal_445, signal_444, signal_443, signal_199}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_448, signal_447, signal_446, signal_200}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_186 ( .a ({signal_442, signal_441, signal_440, signal_198}), .b ({signal_445, signal_444, signal_443, signal_199}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_451, signal_450, signal_449, signal_201}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_189 ( .a ({signal_439, signal_438, signal_437, signal_197}), .b ({signal_454, signal_453, signal_452, signal_202}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_460, signal_459, signal_458, signal_204}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_191 ( .a ({signal_962, signal_960, signal_958, signal_956}), .b ({signal_448, signal_447, signal_446, signal_200}), .c ({signal_466, signal_465, signal_464, signal_206}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_192 ( .a ({signal_970, signal_968, signal_966, signal_964}), .b ({signal_448, signal_447, signal_446, signal_200}), .c ({signal_469, signal_468, signal_467, signal_207}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_193 ( .a ({signal_448, signal_447, signal_446, signal_200}), .b ({signal_978, signal_976, signal_974, signal_972}), .c ({signal_472, signal_471, signal_470, signal_208}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_198 ( .a ({signal_448, signal_447, signal_446, signal_200}), .b ({signal_986, signal_984, signal_982, signal_980}), .c ({signal_487, signal_486, signal_485, signal_213}) ) ;
    buf_clk cell_301 ( .C (clk), .D (signal_955), .Q (signal_956) ) ;
    buf_clk cell_303 ( .C (clk), .D (signal_957), .Q (signal_958) ) ;
    buf_clk cell_305 ( .C (clk), .D (signal_959), .Q (signal_960) ) ;
    buf_clk cell_307 ( .C (clk), .D (signal_961), .Q (signal_962) ) ;
    buf_clk cell_309 ( .C (clk), .D (signal_963), .Q (signal_964) ) ;
    buf_clk cell_311 ( .C (clk), .D (signal_965), .Q (signal_966) ) ;
    buf_clk cell_313 ( .C (clk), .D (signal_967), .Q (signal_968) ) ;
    buf_clk cell_315 ( .C (clk), .D (signal_969), .Q (signal_970) ) ;
    buf_clk cell_317 ( .C (clk), .D (signal_971), .Q (signal_972) ) ;
    buf_clk cell_319 ( .C (clk), .D (signal_973), .Q (signal_974) ) ;
    buf_clk cell_321 ( .C (clk), .D (signal_975), .Q (signal_976) ) ;
    buf_clk cell_323 ( .C (clk), .D (signal_977), .Q (signal_978) ) ;
    buf_clk cell_325 ( .C (clk), .D (signal_979), .Q (signal_980) ) ;
    buf_clk cell_327 ( .C (clk), .D (signal_981), .Q (signal_982) ) ;
    buf_clk cell_329 ( .C (clk), .D (signal_983), .Q (signal_984) ) ;
    buf_clk cell_331 ( .C (clk), .D (signal_985), .Q (signal_986) ) ;
    buf_clk cell_367 ( .C (clk), .D (signal_1021), .Q (signal_1022) ) ;
    buf_clk cell_373 ( .C (clk), .D (signal_1027), .Q (signal_1028) ) ;
    buf_clk cell_379 ( .C (clk), .D (signal_1033), .Q (signal_1034) ) ;
    buf_clk cell_385 ( .C (clk), .D (signal_1039), .Q (signal_1040) ) ;
    buf_clk cell_391 ( .C (clk), .D (signal_1045), .Q (signal_1046) ) ;
    buf_clk cell_397 ( .C (clk), .D (signal_1051), .Q (signal_1052) ) ;
    buf_clk cell_403 ( .C (clk), .D (signal_1057), .Q (signal_1058) ) ;
    buf_clk cell_409 ( .C (clk), .D (signal_1063), .Q (signal_1064) ) ;
    buf_clk cell_415 ( .C (clk), .D (signal_1069), .Q (signal_1070) ) ;
    buf_clk cell_421 ( .C (clk), .D (signal_1075), .Q (signal_1076) ) ;
    buf_clk cell_427 ( .C (clk), .D (signal_1081), .Q (signal_1082) ) ;
    buf_clk cell_433 ( .C (clk), .D (signal_1087), .Q (signal_1088) ) ;
    buf_clk cell_439 ( .C (clk), .D (signal_1093), .Q (signal_1094) ) ;
    buf_clk cell_445 ( .C (clk), .D (signal_1099), .Q (signal_1100) ) ;
    buf_clk cell_451 ( .C (clk), .D (signal_1105), .Q (signal_1106) ) ;
    buf_clk cell_457 ( .C (clk), .D (signal_1111), .Q (signal_1112) ) ;
    buf_clk cell_463 ( .C (clk), .D (signal_1117), .Q (signal_1118) ) ;
    buf_clk cell_469 ( .C (clk), .D (signal_1123), .Q (signal_1124) ) ;
    buf_clk cell_475 ( .C (clk), .D (signal_1129), .Q (signal_1130) ) ;
    buf_clk cell_481 ( .C (clk), .D (signal_1135), .Q (signal_1136) ) ;
    buf_clk cell_487 ( .C (clk), .D (signal_1141), .Q (signal_1142) ) ;
    buf_clk cell_493 ( .C (clk), .D (signal_1147), .Q (signal_1148) ) ;
    buf_clk cell_499 ( .C (clk), .D (signal_1153), .Q (signal_1154) ) ;
    buf_clk cell_505 ( .C (clk), .D (signal_1159), .Q (signal_1160) ) ;
    buf_clk cell_511 ( .C (clk), .D (signal_1165), .Q (signal_1166) ) ;
    buf_clk cell_517 ( .C (clk), .D (signal_1171), .Q (signal_1172) ) ;
    buf_clk cell_523 ( .C (clk), .D (signal_1177), .Q (signal_1178) ) ;
    buf_clk cell_529 ( .C (clk), .D (signal_1183), .Q (signal_1184) ) ;
    buf_clk cell_535 ( .C (clk), .D (signal_1189), .Q (signal_1190) ) ;
    buf_clk cell_541 ( .C (clk), .D (signal_1195), .Q (signal_1196) ) ;
    buf_clk cell_547 ( .C (clk), .D (signal_1201), .Q (signal_1202) ) ;
    buf_clk cell_553 ( .C (clk), .D (signal_1207), .Q (signal_1208) ) ;
    buf_clk cell_559 ( .C (clk), .D (signal_1213), .Q (signal_1214) ) ;
    buf_clk cell_565 ( .C (clk), .D (signal_1219), .Q (signal_1220) ) ;
    buf_clk cell_571 ( .C (clk), .D (signal_1225), .Q (signal_1226) ) ;
    buf_clk cell_577 ( .C (clk), .D (signal_1231), .Q (signal_1232) ) ;
    buf_clk cell_583 ( .C (clk), .D (signal_1237), .Q (signal_1238) ) ;
    buf_clk cell_589 ( .C (clk), .D (signal_1243), .Q (signal_1244) ) ;
    buf_clk cell_595 ( .C (clk), .D (signal_1249), .Q (signal_1250) ) ;
    buf_clk cell_601 ( .C (clk), .D (signal_1255), .Q (signal_1256) ) ;
    buf_clk cell_607 ( .C (clk), .D (signal_1261), .Q (signal_1262) ) ;
    buf_clk cell_613 ( .C (clk), .D (signal_1267), .Q (signal_1268) ) ;
    buf_clk cell_619 ( .C (clk), .D (signal_1273), .Q (signal_1274) ) ;
    buf_clk cell_625 ( .C (clk), .D (signal_1279), .Q (signal_1280) ) ;
    buf_clk cell_631 ( .C (clk), .D (signal_1285), .Q (signal_1286) ) ;
    buf_clk cell_637 ( .C (clk), .D (signal_1291), .Q (signal_1292) ) ;
    buf_clk cell_643 ( .C (clk), .D (signal_1297), .Q (signal_1298) ) ;
    buf_clk cell_649 ( .C (clk), .D (signal_1303), .Q (signal_1304) ) ;
    buf_clk cell_655 ( .C (clk), .D (signal_1309), .Q (signal_1310) ) ;
    buf_clk cell_661 ( .C (clk), .D (signal_1315), .Q (signal_1316) ) ;
    buf_clk cell_667 ( .C (clk), .D (signal_1321), .Q (signal_1322) ) ;
    buf_clk cell_673 ( .C (clk), .D (signal_1327), .Q (signal_1328) ) ;
    buf_clk cell_679 ( .C (clk), .D (signal_1333), .Q (signal_1334) ) ;
    buf_clk cell_685 ( .C (clk), .D (signal_1339), .Q (signal_1340) ) ;
    buf_clk cell_691 ( .C (clk), .D (signal_1345), .Q (signal_1346) ) ;
    buf_clk cell_697 ( .C (clk), .D (signal_1351), .Q (signal_1352) ) ;
    buf_clk cell_703 ( .C (clk), .D (signal_1357), .Q (signal_1358) ) ;
    buf_clk cell_709 ( .C (clk), .D (signal_1363), .Q (signal_1364) ) ;
    buf_clk cell_715 ( .C (clk), .D (signal_1369), .Q (signal_1370) ) ;
    buf_clk cell_721 ( .C (clk), .D (signal_1375), .Q (signal_1376) ) ;
    buf_clk cell_727 ( .C (clk), .D (signal_1381), .Q (signal_1382) ) ;
    buf_clk cell_733 ( .C (clk), .D (signal_1387), .Q (signal_1388) ) ;
    buf_clk cell_739 ( .C (clk), .D (signal_1393), .Q (signal_1394) ) ;
    buf_clk cell_745 ( .C (clk), .D (signal_1399), .Q (signal_1400) ) ;
    buf_clk cell_751 ( .C (clk), .D (signal_1405), .Q (signal_1406) ) ;
    buf_clk cell_757 ( .C (clk), .D (signal_1411), .Q (signal_1412) ) ;
    buf_clk cell_763 ( .C (clk), .D (signal_1417), .Q (signal_1418) ) ;
    buf_clk cell_769 ( .C (clk), .D (signal_1423), .Q (signal_1424) ) ;
    buf_clk cell_775 ( .C (clk), .D (signal_1429), .Q (signal_1430) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_1435), .Q (signal_1436) ) ;
    buf_clk cell_787 ( .C (clk), .D (signal_1441), .Q (signal_1442) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_1447), .Q (signal_1448) ) ;

    /* cells in depth 5 */
    buf_clk cell_332 ( .C (clk), .D (signal_956), .Q (signal_987) ) ;
    buf_clk cell_334 ( .C (clk), .D (signal_958), .Q (signal_989) ) ;
    buf_clk cell_336 ( .C (clk), .D (signal_960), .Q (signal_991) ) ;
    buf_clk cell_338 ( .C (clk), .D (signal_962), .Q (signal_993) ) ;
    buf_clk cell_340 ( .C (clk), .D (signal_208), .Q (signal_995) ) ;
    buf_clk cell_342 ( .C (clk), .D (signal_470), .Q (signal_997) ) ;
    buf_clk cell_344 ( .C (clk), .D (signal_471), .Q (signal_999) ) ;
    buf_clk cell_346 ( .C (clk), .D (signal_472), .Q (signal_1001) ) ;
    buf_clk cell_348 ( .C (clk), .D (signal_964), .Q (signal_1003) ) ;
    buf_clk cell_350 ( .C (clk), .D (signal_966), .Q (signal_1005) ) ;
    buf_clk cell_352 ( .C (clk), .D (signal_968), .Q (signal_1007) ) ;
    buf_clk cell_354 ( .C (clk), .D (signal_970), .Q (signal_1009) ) ;
    buf_clk cell_356 ( .C (clk), .D (signal_213), .Q (signal_1011) ) ;
    buf_clk cell_358 ( .C (clk), .D (signal_485), .Q (signal_1013) ) ;
    buf_clk cell_360 ( .C (clk), .D (signal_486), .Q (signal_1015) ) ;
    buf_clk cell_362 ( .C (clk), .D (signal_487), .Q (signal_1017) ) ;
    buf_clk cell_368 ( .C (clk), .D (signal_1022), .Q (signal_1023) ) ;
    buf_clk cell_374 ( .C (clk), .D (signal_1028), .Q (signal_1029) ) ;
    buf_clk cell_380 ( .C (clk), .D (signal_1034), .Q (signal_1035) ) ;
    buf_clk cell_386 ( .C (clk), .D (signal_1040), .Q (signal_1041) ) ;
    buf_clk cell_392 ( .C (clk), .D (signal_1046), .Q (signal_1047) ) ;
    buf_clk cell_398 ( .C (clk), .D (signal_1052), .Q (signal_1053) ) ;
    buf_clk cell_404 ( .C (clk), .D (signal_1058), .Q (signal_1059) ) ;
    buf_clk cell_410 ( .C (clk), .D (signal_1064), .Q (signal_1065) ) ;
    buf_clk cell_416 ( .C (clk), .D (signal_1070), .Q (signal_1071) ) ;
    buf_clk cell_422 ( .C (clk), .D (signal_1076), .Q (signal_1077) ) ;
    buf_clk cell_428 ( .C (clk), .D (signal_1082), .Q (signal_1083) ) ;
    buf_clk cell_434 ( .C (clk), .D (signal_1088), .Q (signal_1089) ) ;
    buf_clk cell_440 ( .C (clk), .D (signal_1094), .Q (signal_1095) ) ;
    buf_clk cell_446 ( .C (clk), .D (signal_1100), .Q (signal_1101) ) ;
    buf_clk cell_452 ( .C (clk), .D (signal_1106), .Q (signal_1107) ) ;
    buf_clk cell_458 ( .C (clk), .D (signal_1112), .Q (signal_1113) ) ;
    buf_clk cell_464 ( .C (clk), .D (signal_1118), .Q (signal_1119) ) ;
    buf_clk cell_470 ( .C (clk), .D (signal_1124), .Q (signal_1125) ) ;
    buf_clk cell_476 ( .C (clk), .D (signal_1130), .Q (signal_1131) ) ;
    buf_clk cell_482 ( .C (clk), .D (signal_1136), .Q (signal_1137) ) ;
    buf_clk cell_488 ( .C (clk), .D (signal_1142), .Q (signal_1143) ) ;
    buf_clk cell_494 ( .C (clk), .D (signal_1148), .Q (signal_1149) ) ;
    buf_clk cell_500 ( .C (clk), .D (signal_1154), .Q (signal_1155) ) ;
    buf_clk cell_506 ( .C (clk), .D (signal_1160), .Q (signal_1161) ) ;
    buf_clk cell_512 ( .C (clk), .D (signal_1166), .Q (signal_1167) ) ;
    buf_clk cell_518 ( .C (clk), .D (signal_1172), .Q (signal_1173) ) ;
    buf_clk cell_524 ( .C (clk), .D (signal_1178), .Q (signal_1179) ) ;
    buf_clk cell_530 ( .C (clk), .D (signal_1184), .Q (signal_1185) ) ;
    buf_clk cell_536 ( .C (clk), .D (signal_1190), .Q (signal_1191) ) ;
    buf_clk cell_542 ( .C (clk), .D (signal_1196), .Q (signal_1197) ) ;
    buf_clk cell_548 ( .C (clk), .D (signal_1202), .Q (signal_1203) ) ;
    buf_clk cell_554 ( .C (clk), .D (signal_1208), .Q (signal_1209) ) ;
    buf_clk cell_560 ( .C (clk), .D (signal_1214), .Q (signal_1215) ) ;
    buf_clk cell_566 ( .C (clk), .D (signal_1220), .Q (signal_1221) ) ;
    buf_clk cell_572 ( .C (clk), .D (signal_1226), .Q (signal_1227) ) ;
    buf_clk cell_578 ( .C (clk), .D (signal_1232), .Q (signal_1233) ) ;
    buf_clk cell_584 ( .C (clk), .D (signal_1238), .Q (signal_1239) ) ;
    buf_clk cell_590 ( .C (clk), .D (signal_1244), .Q (signal_1245) ) ;
    buf_clk cell_596 ( .C (clk), .D (signal_1250), .Q (signal_1251) ) ;
    buf_clk cell_602 ( .C (clk), .D (signal_1256), .Q (signal_1257) ) ;
    buf_clk cell_608 ( .C (clk), .D (signal_1262), .Q (signal_1263) ) ;
    buf_clk cell_614 ( .C (clk), .D (signal_1268), .Q (signal_1269) ) ;
    buf_clk cell_620 ( .C (clk), .D (signal_1274), .Q (signal_1275) ) ;
    buf_clk cell_626 ( .C (clk), .D (signal_1280), .Q (signal_1281) ) ;
    buf_clk cell_632 ( .C (clk), .D (signal_1286), .Q (signal_1287) ) ;
    buf_clk cell_638 ( .C (clk), .D (signal_1292), .Q (signal_1293) ) ;
    buf_clk cell_644 ( .C (clk), .D (signal_1298), .Q (signal_1299) ) ;
    buf_clk cell_650 ( .C (clk), .D (signal_1304), .Q (signal_1305) ) ;
    buf_clk cell_656 ( .C (clk), .D (signal_1310), .Q (signal_1311) ) ;
    buf_clk cell_662 ( .C (clk), .D (signal_1316), .Q (signal_1317) ) ;
    buf_clk cell_668 ( .C (clk), .D (signal_1322), .Q (signal_1323) ) ;
    buf_clk cell_674 ( .C (clk), .D (signal_1328), .Q (signal_1329) ) ;
    buf_clk cell_680 ( .C (clk), .D (signal_1334), .Q (signal_1335) ) ;
    buf_clk cell_686 ( .C (clk), .D (signal_1340), .Q (signal_1341) ) ;
    buf_clk cell_692 ( .C (clk), .D (signal_1346), .Q (signal_1347) ) ;
    buf_clk cell_698 ( .C (clk), .D (signal_1352), .Q (signal_1353) ) ;
    buf_clk cell_704 ( .C (clk), .D (signal_1358), .Q (signal_1359) ) ;
    buf_clk cell_710 ( .C (clk), .D (signal_1364), .Q (signal_1365) ) ;
    buf_clk cell_716 ( .C (clk), .D (signal_1370), .Q (signal_1371) ) ;
    buf_clk cell_722 ( .C (clk), .D (signal_1376), .Q (signal_1377) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_1382), .Q (signal_1383) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_1388), .Q (signal_1389) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_1394), .Q (signal_1395) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_1400), .Q (signal_1401) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_1406), .Q (signal_1407) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_1412), .Q (signal_1413) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_1418), .Q (signal_1419) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_1424), .Q (signal_1425) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_1430), .Q (signal_1431) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_1436), .Q (signal_1437) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_1442), .Q (signal_1443) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_1448), .Q (signal_1449) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_194 ( .a ({signal_978, signal_976, signal_974, signal_972}), .b ({signal_469, signal_468, signal_467, signal_207}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_475, signal_474, signal_473, signal_209}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_195 ( .a ({signal_986, signal_984, signal_982, signal_980}), .b ({signal_466, signal_465, signal_464, signal_206}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_478, signal_477, signal_476, signal_210}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_196 ( .a ({signal_978, signal_976, signal_974, signal_972}), .b ({signal_460, signal_459, signal_458, signal_204}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_481, signal_480, signal_479, signal_211}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_197 ( .a ({signal_451, signal_450, signal_449, signal_201}), .b ({signal_986, signal_984, signal_982, signal_980}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_484, signal_483, signal_482, signal_212}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_199 ( .a ({signal_994, signal_992, signal_990, signal_988}), .b ({signal_475, signal_474, signal_473, signal_209}), .c ({signal_490, signal_489, signal_488, signal_214}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_200 ( .a ({signal_1002, signal_1000, signal_998, signal_996}), .b ({signal_481, signal_480, signal_479, signal_211}), .c ({signal_493, signal_492, signal_491, signal_215}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_201 ( .a ({signal_1010, signal_1008, signal_1006, signal_1004}), .b ({signal_478, signal_477, signal_476, signal_210}), .c ({signal_496, signal_495, signal_494, signal_216}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_202 ( .a ({signal_484, signal_483, signal_482, signal_212}), .b ({signal_1018, signal_1016, signal_1014, signal_1012}), .c ({signal_499, signal_498, signal_497, signal_217}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_211 ( .a ({signal_493, signal_492, signal_491, signal_215}), .b ({signal_499, signal_498, signal_497, signal_217}), .c ({signal_526, signal_525, signal_524, signal_226}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_212 ( .a ({signal_490, signal_489, signal_488, signal_214}), .b ({signal_496, signal_495, signal_494, signal_216}), .c ({signal_529, signal_528, signal_527, signal_227}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_213 ( .a ({signal_490, signal_489, signal_488, signal_214}), .b ({signal_493, signal_492, signal_491, signal_215}), .c ({signal_532, signal_531, signal_530, signal_228}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_214 ( .a ({signal_496, signal_495, signal_494, signal_216}), .b ({signal_499, signal_498, signal_497, signal_217}), .c ({signal_535, signal_534, signal_533, signal_229}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_223 ( .a ({signal_526, signal_525, signal_524, signal_226}), .b ({signal_529, signal_528, signal_527, signal_227}), .c ({signal_562, signal_561, signal_560, signal_238}) ) ;
    buf_clk cell_333 ( .C (clk), .D (signal_987), .Q (signal_988) ) ;
    buf_clk cell_335 ( .C (clk), .D (signal_989), .Q (signal_990) ) ;
    buf_clk cell_337 ( .C (clk), .D (signal_991), .Q (signal_992) ) ;
    buf_clk cell_339 ( .C (clk), .D (signal_993), .Q (signal_994) ) ;
    buf_clk cell_341 ( .C (clk), .D (signal_995), .Q (signal_996) ) ;
    buf_clk cell_343 ( .C (clk), .D (signal_997), .Q (signal_998) ) ;
    buf_clk cell_345 ( .C (clk), .D (signal_999), .Q (signal_1000) ) ;
    buf_clk cell_347 ( .C (clk), .D (signal_1001), .Q (signal_1002) ) ;
    buf_clk cell_349 ( .C (clk), .D (signal_1003), .Q (signal_1004) ) ;
    buf_clk cell_351 ( .C (clk), .D (signal_1005), .Q (signal_1006) ) ;
    buf_clk cell_353 ( .C (clk), .D (signal_1007), .Q (signal_1008) ) ;
    buf_clk cell_355 ( .C (clk), .D (signal_1009), .Q (signal_1010) ) ;
    buf_clk cell_357 ( .C (clk), .D (signal_1011), .Q (signal_1012) ) ;
    buf_clk cell_359 ( .C (clk), .D (signal_1013), .Q (signal_1014) ) ;
    buf_clk cell_361 ( .C (clk), .D (signal_1015), .Q (signal_1016) ) ;
    buf_clk cell_363 ( .C (clk), .D (signal_1017), .Q (signal_1018) ) ;
    buf_clk cell_369 ( .C (clk), .D (signal_1023), .Q (signal_1024) ) ;
    buf_clk cell_375 ( .C (clk), .D (signal_1029), .Q (signal_1030) ) ;
    buf_clk cell_381 ( .C (clk), .D (signal_1035), .Q (signal_1036) ) ;
    buf_clk cell_387 ( .C (clk), .D (signal_1041), .Q (signal_1042) ) ;
    buf_clk cell_393 ( .C (clk), .D (signal_1047), .Q (signal_1048) ) ;
    buf_clk cell_399 ( .C (clk), .D (signal_1053), .Q (signal_1054) ) ;
    buf_clk cell_405 ( .C (clk), .D (signal_1059), .Q (signal_1060) ) ;
    buf_clk cell_411 ( .C (clk), .D (signal_1065), .Q (signal_1066) ) ;
    buf_clk cell_417 ( .C (clk), .D (signal_1071), .Q (signal_1072) ) ;
    buf_clk cell_423 ( .C (clk), .D (signal_1077), .Q (signal_1078) ) ;
    buf_clk cell_429 ( .C (clk), .D (signal_1083), .Q (signal_1084) ) ;
    buf_clk cell_435 ( .C (clk), .D (signal_1089), .Q (signal_1090) ) ;
    buf_clk cell_441 ( .C (clk), .D (signal_1095), .Q (signal_1096) ) ;
    buf_clk cell_447 ( .C (clk), .D (signal_1101), .Q (signal_1102) ) ;
    buf_clk cell_453 ( .C (clk), .D (signal_1107), .Q (signal_1108) ) ;
    buf_clk cell_459 ( .C (clk), .D (signal_1113), .Q (signal_1114) ) ;
    buf_clk cell_465 ( .C (clk), .D (signal_1119), .Q (signal_1120) ) ;
    buf_clk cell_471 ( .C (clk), .D (signal_1125), .Q (signal_1126) ) ;
    buf_clk cell_477 ( .C (clk), .D (signal_1131), .Q (signal_1132) ) ;
    buf_clk cell_483 ( .C (clk), .D (signal_1137), .Q (signal_1138) ) ;
    buf_clk cell_489 ( .C (clk), .D (signal_1143), .Q (signal_1144) ) ;
    buf_clk cell_495 ( .C (clk), .D (signal_1149), .Q (signal_1150) ) ;
    buf_clk cell_501 ( .C (clk), .D (signal_1155), .Q (signal_1156) ) ;
    buf_clk cell_507 ( .C (clk), .D (signal_1161), .Q (signal_1162) ) ;
    buf_clk cell_513 ( .C (clk), .D (signal_1167), .Q (signal_1168) ) ;
    buf_clk cell_519 ( .C (clk), .D (signal_1173), .Q (signal_1174) ) ;
    buf_clk cell_525 ( .C (clk), .D (signal_1179), .Q (signal_1180) ) ;
    buf_clk cell_531 ( .C (clk), .D (signal_1185), .Q (signal_1186) ) ;
    buf_clk cell_537 ( .C (clk), .D (signal_1191), .Q (signal_1192) ) ;
    buf_clk cell_543 ( .C (clk), .D (signal_1197), .Q (signal_1198) ) ;
    buf_clk cell_549 ( .C (clk), .D (signal_1203), .Q (signal_1204) ) ;
    buf_clk cell_555 ( .C (clk), .D (signal_1209), .Q (signal_1210) ) ;
    buf_clk cell_561 ( .C (clk), .D (signal_1215), .Q (signal_1216) ) ;
    buf_clk cell_567 ( .C (clk), .D (signal_1221), .Q (signal_1222) ) ;
    buf_clk cell_573 ( .C (clk), .D (signal_1227), .Q (signal_1228) ) ;
    buf_clk cell_579 ( .C (clk), .D (signal_1233), .Q (signal_1234) ) ;
    buf_clk cell_585 ( .C (clk), .D (signal_1239), .Q (signal_1240) ) ;
    buf_clk cell_591 ( .C (clk), .D (signal_1245), .Q (signal_1246) ) ;
    buf_clk cell_597 ( .C (clk), .D (signal_1251), .Q (signal_1252) ) ;
    buf_clk cell_603 ( .C (clk), .D (signal_1257), .Q (signal_1258) ) ;
    buf_clk cell_609 ( .C (clk), .D (signal_1263), .Q (signal_1264) ) ;
    buf_clk cell_615 ( .C (clk), .D (signal_1269), .Q (signal_1270) ) ;
    buf_clk cell_621 ( .C (clk), .D (signal_1275), .Q (signal_1276) ) ;
    buf_clk cell_627 ( .C (clk), .D (signal_1281), .Q (signal_1282) ) ;
    buf_clk cell_633 ( .C (clk), .D (signal_1287), .Q (signal_1288) ) ;
    buf_clk cell_639 ( .C (clk), .D (signal_1293), .Q (signal_1294) ) ;
    buf_clk cell_645 ( .C (clk), .D (signal_1299), .Q (signal_1300) ) ;
    buf_clk cell_651 ( .C (clk), .D (signal_1305), .Q (signal_1306) ) ;
    buf_clk cell_657 ( .C (clk), .D (signal_1311), .Q (signal_1312) ) ;
    buf_clk cell_663 ( .C (clk), .D (signal_1317), .Q (signal_1318) ) ;
    buf_clk cell_669 ( .C (clk), .D (signal_1323), .Q (signal_1324) ) ;
    buf_clk cell_675 ( .C (clk), .D (signal_1329), .Q (signal_1330) ) ;
    buf_clk cell_681 ( .C (clk), .D (signal_1335), .Q (signal_1336) ) ;
    buf_clk cell_687 ( .C (clk), .D (signal_1341), .Q (signal_1342) ) ;
    buf_clk cell_693 ( .C (clk), .D (signal_1347), .Q (signal_1348) ) ;
    buf_clk cell_699 ( .C (clk), .D (signal_1353), .Q (signal_1354) ) ;
    buf_clk cell_705 ( .C (clk), .D (signal_1359), .Q (signal_1360) ) ;
    buf_clk cell_711 ( .C (clk), .D (signal_1365), .Q (signal_1366) ) ;
    buf_clk cell_717 ( .C (clk), .D (signal_1371), .Q (signal_1372) ) ;
    buf_clk cell_723 ( .C (clk), .D (signal_1377), .Q (signal_1378) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_1383), .Q (signal_1384) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_1389), .Q (signal_1390) ) ;
    buf_clk cell_741 ( .C (clk), .D (signal_1395), .Q (signal_1396) ) ;
    buf_clk cell_747 ( .C (clk), .D (signal_1401), .Q (signal_1402) ) ;
    buf_clk cell_753 ( .C (clk), .D (signal_1407), .Q (signal_1408) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_1413), .Q (signal_1414) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_1419), .Q (signal_1420) ) ;
    buf_clk cell_771 ( .C (clk), .D (signal_1425), .Q (signal_1426) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_1431), .Q (signal_1432) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_1437), .Q (signal_1438) ) ;
    buf_clk cell_789 ( .C (clk), .D (signal_1443), .Q (signal_1444) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_1449), .Q (signal_1450) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_203 ( .a ({signal_1042, signal_1036, signal_1030, signal_1024}), .b ({signal_499, signal_498, signal_497, signal_217}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_502, signal_501, signal_500, signal_218}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_204 ( .a ({signal_1066, signal_1060, signal_1054, signal_1048}), .b ({signal_496, signal_495, signal_494, signal_216}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_505, signal_504, signal_503, signal_219}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_205 ( .a ({signal_1090, signal_1084, signal_1078, signal_1072}), .b ({signal_493, signal_492, signal_491, signal_215}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_508, signal_507, signal_506, signal_220}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_206 ( .a ({signal_1114, signal_1108, signal_1102, signal_1096}), .b ({signal_490, signal_489, signal_488, signal_214}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_511, signal_510, signal_509, signal_221}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_207 ( .a ({signal_1138, signal_1132, signal_1126, signal_1120}), .b ({signal_499, signal_498, signal_497, signal_217}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_514, signal_513, signal_512, signal_222}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_208 ( .a ({signal_1162, signal_1156, signal_1150, signal_1144}), .b ({signal_496, signal_495, signal_494, signal_216}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_517, signal_516, signal_515, signal_223}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_209 ( .a ({signal_1186, signal_1180, signal_1174, signal_1168}), .b ({signal_493, signal_492, signal_491, signal_215}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_520, signal_519, signal_518, signal_224}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_210 ( .a ({signal_1210, signal_1204, signal_1198, signal_1192}), .b ({signal_490, signal_489, signal_488, signal_214}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_523, signal_522, signal_521, signal_225}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_215 ( .a ({signal_1234, signal_1228, signal_1222, signal_1216}), .b ({signal_535, signal_534, signal_533, signal_229}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_538, signal_537, signal_536, signal_230}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_216 ( .a ({signal_1258, signal_1252, signal_1246, signal_1240}), .b ({signal_532, signal_531, signal_530, signal_228}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_541, signal_540, signal_539, signal_231}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_217 ( .a ({signal_1282, signal_1276, signal_1270, signal_1264}), .b ({signal_529, signal_528, signal_527, signal_227}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_544, signal_543, signal_542, signal_232}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_218 ( .a ({signal_1306, signal_1300, signal_1294, signal_1288}), .b ({signal_526, signal_525, signal_524, signal_226}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_547, signal_546, signal_545, signal_233}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_219 ( .a ({signal_1330, signal_1324, signal_1318, signal_1312}), .b ({signal_535, signal_534, signal_533, signal_229}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_550, signal_549, signal_548, signal_234}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_220 ( .a ({signal_1354, signal_1348, signal_1342, signal_1336}), .b ({signal_532, signal_531, signal_530, signal_228}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_553, signal_552, signal_551, signal_235}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_221 ( .a ({signal_1378, signal_1372, signal_1366, signal_1360}), .b ({signal_529, signal_528, signal_527, signal_227}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_556, signal_555, signal_554, signal_236}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_222 ( .a ({signal_1402, signal_1396, signal_1390, signal_1384}), .b ({signal_526, signal_525, signal_524, signal_226}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_559, signal_558, signal_557, signal_237}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_224 ( .a ({signal_508, signal_507, signal_506, signal_220}), .b ({signal_514, signal_513, signal_512, signal_222}), .c ({signal_565, signal_564, signal_563, signal_239}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_225 ( .a ({signal_511, signal_510, signal_509, signal_221}), .b ({signal_520, signal_519, signal_518, signal_224}), .c ({signal_568, signal_567, signal_566, signal_240}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_226 ( .a ({signal_505, signal_504, signal_503, signal_219}), .b ({signal_511, signal_510, signal_509, signal_221}), .c ({signal_571, signal_570, signal_569, signal_241}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_227 ( .a ({signal_1426, signal_1420, signal_1414, signal_1408}), .b ({signal_562, signal_561, signal_560, signal_238}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_574, signal_573, signal_572, signal_242}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(1)) cell_228 ( .a ({signal_1450, signal_1444, signal_1438, signal_1432}), .b ({signal_562, signal_561, signal_560, signal_238}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_577, signal_576, signal_575, signal_243}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_229 ( .a ({signal_505, signal_504, signal_503, signal_219}), .b ({signal_538, signal_537, signal_536, signal_230}), .c ({signal_580, signal_579, signal_578, signal_244}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_230 ( .a ({signal_502, signal_501, signal_500, signal_218}), .b ({signal_550, signal_549, signal_548, signal_234}), .c ({signal_583, signal_582, signal_581, signal_245}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_231 ( .a ({signal_547, signal_546, signal_545, signal_233}), .b ({signal_553, signal_552, signal_551, signal_235}), .c ({signal_586, signal_585, signal_584, signal_246}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_232 ( .a ({signal_541, signal_540, signal_539, signal_231}), .b ({signal_556, signal_555, signal_554, signal_236}), .c ({signal_589, signal_588, signal_587, signal_247}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_233 ( .a ({signal_544, signal_543, signal_542, signal_232}), .b ({signal_556, signal_555, signal_554, signal_236}), .c ({signal_592, signal_591, signal_590, signal_248}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_234 ( .a ({signal_550, signal_549, signal_548, signal_234}), .b ({signal_565, signal_564, signal_563, signal_239}), .c ({signal_595, signal_594, signal_593, signal_249}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_235 ( .a ({signal_517, signal_516, signal_515, signal_223}), .b ({signal_565, signal_564, signal_563, signal_239}), .c ({signal_598, signal_597, signal_596, signal_250}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_236 ( .a ({signal_553, signal_552, signal_551, signal_235}), .b ({signal_568, signal_567, signal_566, signal_240}), .c ({signal_601, signal_600, signal_599, signal_251}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_237 ( .a ({signal_556, signal_555, signal_554, signal_236}), .b ({signal_577, signal_576, signal_575, signal_243}), .c ({signal_604, signal_603, signal_602, signal_252}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_238 ( .a ({signal_577, signal_576, signal_575, signal_243}), .b ({signal_589, signal_588, signal_587, signal_247}), .c ({signal_607, signal_606, signal_605, signal_253}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_239 ( .a ({signal_538, signal_537, signal_536, signal_230}), .b ({signal_583, signal_582, signal_581, signal_245}), .c ({signal_610, signal_609, signal_608, signal_254}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_240 ( .a ({signal_544, signal_543, signal_542, signal_232}), .b ({signal_574, signal_573, signal_572, signal_242}), .c ({signal_613, signal_612, signal_611, signal_255}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_241 ( .a ({signal_574, signal_573, signal_572, signal_242}), .b ({signal_586, signal_585, signal_584, signal_246}), .c ({signal_616, signal_615, signal_614, signal_256}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_242 ( .a ({signal_523, signal_522, signal_521, signal_225}), .b ({signal_580, signal_579, signal_578, signal_244}), .c ({signal_619, signal_618, signal_617, signal_257}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_243 ( .a ({signal_559, signal_558, signal_557, signal_237}), .b ({signal_586, signal_585, signal_584, signal_246}), .c ({signal_622, signal_621, signal_620, signal_258}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_244 ( .a ({signal_571, signal_570, signal_569, signal_241}), .b ({signal_583, signal_582, signal_581, signal_245}), .c ({signal_625, signal_624, signal_623, signal_259}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_245 ( .a ({signal_580, signal_579, signal_578, signal_244}), .b ({signal_601, signal_600, signal_599, signal_251}), .c ({signal_628, signal_627, signal_626, signal_260}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_246 ( .a ({signal_508, signal_507, signal_506, signal_220}), .b ({signal_604, signal_603, signal_602, signal_252}), .c ({signal_631, signal_630, signal_629, signal_261}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_247 ( .a ({signal_514, signal_513, signal_512, signal_222}), .b ({signal_604, signal_603, signal_602, signal_252}), .c ({signal_634, signal_633, signal_632, signal_262}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_248 ( .a ({signal_565, signal_564, signal_563, signal_239}), .b ({signal_604, signal_603, signal_602, signal_252}), .c ({signal_637, signal_636, signal_635, signal_263}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_249 ( .a ({signal_565, signal_564, signal_563, signal_239}), .b ({signal_610, signal_609, signal_608, signal_254}), .c ({signal_640, signal_639, signal_638, signal_264}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_250 ( .a ({signal_595, signal_594, signal_593, signal_249}), .b ({signal_613, signal_612, signal_611, signal_255}), .c ({signal_643, signal_642, signal_641, signal_265}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_251 ( .a ({signal_607, signal_606, signal_605, signal_253}), .b ({signal_616, signal_615, signal_614, signal_256}), .c ({signal_646, signal_645, signal_644, signal_266}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_252 ( .a ({signal_610, signal_609, signal_608, signal_254}), .b ({signal_613, signal_612, signal_611, signal_255}), .c ({signal_649, signal_648, signal_647, signal_267}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_253 ( .a ({signal_568, signal_567, signal_566, signal_240}), .b ({signal_616, signal_615, signal_614, signal_256}), .c ({signal_652, signal_651, signal_650, signal_268}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_254 ( .a ({signal_592, signal_591, signal_590, signal_248}), .b ({signal_619, signal_618, signal_617, signal_257}), .c ({signal_655, signal_654, signal_653, signal_269}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_255 ( .a ({signal_598, signal_597, signal_596, signal_250}), .b ({signal_619, signal_618, signal_617, signal_257}), .c ({signal_658, signal_657, signal_656, signal_270}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_256 ( .a ({signal_607, signal_606, signal_605, signal_253}), .b ({signal_628, signal_627, signal_626, signal_260}), .c ({signal_661, signal_660, signal_659, signal_271}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_257 ( .a ({signal_661, signal_660, signal_659, signal_271}), .b ({signal_664, signal_663, signal_662, signal_150}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_258 ( .a ({signal_607, signal_606, signal_605, signal_253}), .b ({signal_643, signal_642, signal_641, signal_265}), .c ({signal_667, signal_666, signal_665, signal_143}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_259 ( .a ({signal_634, signal_633, signal_632, signal_262}), .b ({signal_649, signal_648, signal_647, signal_267}), .c ({signal_670, signal_669, signal_668, signal_272}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_260 ( .a ({signal_622, signal_621, signal_620, signal_258}), .b ({signal_655, signal_654, signal_653, signal_269}), .c ({signal_673, signal_672, signal_671, signal_273}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_261 ( .a ({signal_607, signal_606, signal_605, signal_253}), .b ({signal_640, signal_639, signal_638, signal_264}), .c ({signal_676, signal_675, signal_674, signal_146}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_262 ( .a ({signal_625, signal_624, signal_623, signal_259}), .b ({signal_637, signal_636, signal_635, signal_263}), .c ({signal_679, signal_678, signal_677, signal_147}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_263 ( .a ({signal_646, signal_645, signal_644, signal_266}), .b ({signal_658, signal_657, signal_656, signal_270}), .c ({signal_682, signal_681, signal_680, signal_148}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(1)) cell_264 ( .a ({signal_631, signal_630, signal_629, signal_261}), .b ({signal_652, signal_651, signal_650, signal_268}), .c ({signal_685, signal_684, signal_683, signal_274}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_265 ( .a ({signal_670, signal_669, signal_668, signal_272}), .b ({signal_688, signal_687, signal_686, signal_144}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_266 ( .a ({signal_673, signal_672, signal_671, signal_273}), .b ({signal_691, signal_690, signal_689, signal_145}) ) ;
    not_masked #(.security_order(3), .pipeline(1)) cell_267 ( .a ({signal_685, signal_684, signal_683, signal_274}), .b ({signal_694, signal_693, signal_692, signal_149}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_667, signal_666, signal_665, signal_143}), .Q ({Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_688, signal_687, signal_686, signal_144}), .Q ({Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_691, signal_690, signal_689, signal_145}), .Q ({Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_676, signal_675, signal_674, signal_146}), .Q ({Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_679, signal_678, signal_677, signal_147}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_682, signal_681, signal_680, signal_148}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_694, signal_693, signal_692, signal_149}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_664, signal_663, signal_662, signal_150}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
