
module SkinnyTop_HPC2_ClockGating_d1 ( Plaintext_s0, Key_s0, clk, rst, Key_s1, 
        Plaintext_s1, Fresh, Ciphertext_s0, done, Ciphertext_s1, Synch );
  input [63:0] Plaintext_s0;
  input [63:0] Key_s0;
  input [63:0] Key_s1;
  input [63:0] Plaintext_s1;
  input [63:0] Fresh;
  output [63:0] Ciphertext_s0;
  output [63:0] Ciphertext_s1;
  input clk, rst;
  output done, Synch;
  wire   SubCellInst_SboxInst_0_n3, new_AGEMA_signal_1167,
         SubCellInst_SboxInst_0_XX_1_, new_AGEMA_signal_1169,
         SubCellInst_SboxInst_0_XX_2_, new_AGEMA_signal_1453,
         SubCellInst_SboxInst_0_Q0, new_AGEMA_signal_1454,
         SubCellInst_SboxInst_0_Q1, new_AGEMA_signal_1455,
         SubCellInst_SboxInst_0_Q4, new_AGEMA_signal_1456,
         SubCellInst_SboxInst_0_Q6, new_AGEMA_signal_1550,
         SubCellInst_SboxInst_0_L1, new_AGEMA_signal_1457,
         SubCellInst_SboxInst_0_L2, SubCellInst_SboxInst_1_n3,
         new_AGEMA_signal_1173, SubCellInst_SboxInst_1_XX_1_,
         new_AGEMA_signal_1175, SubCellInst_SboxInst_1_XX_2_,
         new_AGEMA_signal_1459, SubCellInst_SboxInst_1_Q0,
         new_AGEMA_signal_1460, SubCellInst_SboxInst_1_Q1,
         new_AGEMA_signal_1461, SubCellInst_SboxInst_1_Q4,
         new_AGEMA_signal_1462, SubCellInst_SboxInst_1_Q6,
         new_AGEMA_signal_1553, SubCellInst_SboxInst_1_L1,
         new_AGEMA_signal_1463, SubCellInst_SboxInst_1_L2,
         SubCellInst_SboxInst_2_n3, new_AGEMA_signal_1179,
         SubCellInst_SboxInst_2_XX_1_, new_AGEMA_signal_1181,
         SubCellInst_SboxInst_2_XX_2_, new_AGEMA_signal_1465,
         SubCellInst_SboxInst_2_Q0, new_AGEMA_signal_1466,
         SubCellInst_SboxInst_2_Q1, new_AGEMA_signal_1467,
         SubCellInst_SboxInst_2_Q4, new_AGEMA_signal_1468,
         SubCellInst_SboxInst_2_Q6, new_AGEMA_signal_1556,
         SubCellInst_SboxInst_2_L1, new_AGEMA_signal_1469,
         SubCellInst_SboxInst_2_L2, SubCellInst_SboxInst_3_n3,
         new_AGEMA_signal_1185, SubCellInst_SboxInst_3_XX_1_,
         new_AGEMA_signal_1187, SubCellInst_SboxInst_3_XX_2_,
         new_AGEMA_signal_1471, SubCellInst_SboxInst_3_Q0,
         new_AGEMA_signal_1472, SubCellInst_SboxInst_3_Q1,
         new_AGEMA_signal_1473, SubCellInst_SboxInst_3_Q4,
         new_AGEMA_signal_1474, SubCellInst_SboxInst_3_Q6,
         new_AGEMA_signal_1559, SubCellInst_SboxInst_3_L1,
         new_AGEMA_signal_1475, SubCellInst_SboxInst_3_L2,
         SubCellInst_SboxInst_4_n3, new_AGEMA_signal_1191,
         SubCellInst_SboxInst_4_XX_1_, new_AGEMA_signal_1193,
         SubCellInst_SboxInst_4_XX_2_, new_AGEMA_signal_1477,
         SubCellInst_SboxInst_4_Q0, new_AGEMA_signal_1478,
         SubCellInst_SboxInst_4_Q1, new_AGEMA_signal_1479,
         SubCellInst_SboxInst_4_Q4, new_AGEMA_signal_1480,
         SubCellInst_SboxInst_4_Q6, new_AGEMA_signal_1562,
         SubCellInst_SboxInst_4_L1, new_AGEMA_signal_1481,
         SubCellInst_SboxInst_4_L2, SubCellInst_SboxInst_5_n3,
         new_AGEMA_signal_1197, SubCellInst_SboxInst_5_XX_1_,
         new_AGEMA_signal_1199, SubCellInst_SboxInst_5_XX_2_,
         new_AGEMA_signal_1483, SubCellInst_SboxInst_5_Q0,
         new_AGEMA_signal_1484, SubCellInst_SboxInst_5_Q1,
         new_AGEMA_signal_1485, SubCellInst_SboxInst_5_Q4,
         new_AGEMA_signal_1486, SubCellInst_SboxInst_5_Q6,
         new_AGEMA_signal_1565, SubCellInst_SboxInst_5_L1,
         new_AGEMA_signal_1487, SubCellInst_SboxInst_5_L2,
         SubCellInst_SboxInst_6_n3, new_AGEMA_signal_1203,
         SubCellInst_SboxInst_6_XX_1_, new_AGEMA_signal_1205,
         SubCellInst_SboxInst_6_XX_2_, new_AGEMA_signal_1489,
         SubCellInst_SboxInst_6_Q0, new_AGEMA_signal_1490,
         SubCellInst_SboxInst_6_Q1, new_AGEMA_signal_1491,
         SubCellInst_SboxInst_6_Q4, new_AGEMA_signal_1492,
         SubCellInst_SboxInst_6_Q6, new_AGEMA_signal_1568,
         SubCellInst_SboxInst_6_L1, new_AGEMA_signal_1493,
         SubCellInst_SboxInst_6_L2, SubCellInst_SboxInst_7_n3,
         new_AGEMA_signal_1209, SubCellInst_SboxInst_7_XX_1_,
         new_AGEMA_signal_1211, SubCellInst_SboxInst_7_XX_2_,
         new_AGEMA_signal_1495, SubCellInst_SboxInst_7_Q0,
         new_AGEMA_signal_1496, SubCellInst_SboxInst_7_Q1,
         new_AGEMA_signal_1497, SubCellInst_SboxInst_7_Q4,
         new_AGEMA_signal_1498, SubCellInst_SboxInst_7_Q6,
         new_AGEMA_signal_1571, SubCellInst_SboxInst_7_L1,
         new_AGEMA_signal_1499, SubCellInst_SboxInst_7_L2,
         SubCellInst_SboxInst_8_n3, new_AGEMA_signal_1215,
         SubCellInst_SboxInst_8_XX_1_, new_AGEMA_signal_1217,
         SubCellInst_SboxInst_8_XX_2_, new_AGEMA_signal_1501,
         SubCellInst_SboxInst_8_Q0, new_AGEMA_signal_1502,
         SubCellInst_SboxInst_8_Q1, new_AGEMA_signal_1503,
         SubCellInst_SboxInst_8_Q4, new_AGEMA_signal_1504,
         SubCellInst_SboxInst_8_Q6, new_AGEMA_signal_1574,
         SubCellInst_SboxInst_8_L1, new_AGEMA_signal_1505,
         SubCellInst_SboxInst_8_L2, SubCellInst_SboxInst_9_n3,
         new_AGEMA_signal_1221, SubCellInst_SboxInst_9_XX_1_,
         new_AGEMA_signal_1223, SubCellInst_SboxInst_9_XX_2_,
         new_AGEMA_signal_1507, SubCellInst_SboxInst_9_Q0,
         new_AGEMA_signal_1508, SubCellInst_SboxInst_9_Q1,
         new_AGEMA_signal_1509, SubCellInst_SboxInst_9_Q4,
         new_AGEMA_signal_1510, SubCellInst_SboxInst_9_Q6,
         new_AGEMA_signal_1577, SubCellInst_SboxInst_9_L1,
         new_AGEMA_signal_1511, SubCellInst_SboxInst_9_L2,
         SubCellInst_SboxInst_10_n3, new_AGEMA_signal_1227,
         SubCellInst_SboxInst_10_XX_1_, new_AGEMA_signal_1229,
         SubCellInst_SboxInst_10_XX_2_, new_AGEMA_signal_1513,
         SubCellInst_SboxInst_10_Q0, new_AGEMA_signal_1514,
         SubCellInst_SboxInst_10_Q1, new_AGEMA_signal_1515,
         SubCellInst_SboxInst_10_Q4, new_AGEMA_signal_1516,
         SubCellInst_SboxInst_10_Q6, new_AGEMA_signal_1580,
         SubCellInst_SboxInst_10_L1, new_AGEMA_signal_1517,
         SubCellInst_SboxInst_10_L2, SubCellInst_SboxInst_11_n3,
         new_AGEMA_signal_1233, SubCellInst_SboxInst_11_XX_1_,
         new_AGEMA_signal_1235, SubCellInst_SboxInst_11_XX_2_,
         new_AGEMA_signal_1519, SubCellInst_SboxInst_11_Q0,
         new_AGEMA_signal_1520, SubCellInst_SboxInst_11_Q1,
         new_AGEMA_signal_1521, SubCellInst_SboxInst_11_Q4,
         new_AGEMA_signal_1522, SubCellInst_SboxInst_11_Q6,
         new_AGEMA_signal_1583, SubCellInst_SboxInst_11_L1,
         new_AGEMA_signal_1523, SubCellInst_SboxInst_11_L2,
         SubCellInst_SboxInst_12_n3, new_AGEMA_signal_1239,
         SubCellInst_SboxInst_12_XX_1_, new_AGEMA_signal_1241,
         SubCellInst_SboxInst_12_XX_2_, new_AGEMA_signal_1525,
         SubCellInst_SboxInst_12_Q0, new_AGEMA_signal_1526,
         SubCellInst_SboxInst_12_Q1, new_AGEMA_signal_1527,
         SubCellInst_SboxInst_12_Q4, new_AGEMA_signal_1528,
         SubCellInst_SboxInst_12_Q6, new_AGEMA_signal_1586,
         SubCellInst_SboxInst_12_L1, new_AGEMA_signal_1529,
         SubCellInst_SboxInst_12_L2, SubCellInst_SboxInst_13_n3,
         new_AGEMA_signal_1245, SubCellInst_SboxInst_13_XX_1_,
         new_AGEMA_signal_1247, SubCellInst_SboxInst_13_XX_2_,
         new_AGEMA_signal_1531, SubCellInst_SboxInst_13_Q0,
         new_AGEMA_signal_1532, SubCellInst_SboxInst_13_Q1,
         new_AGEMA_signal_1533, SubCellInst_SboxInst_13_Q4,
         new_AGEMA_signal_1534, SubCellInst_SboxInst_13_Q6,
         new_AGEMA_signal_1589, SubCellInst_SboxInst_13_L1,
         new_AGEMA_signal_1535, SubCellInst_SboxInst_13_L2,
         SubCellInst_SboxInst_14_n3, new_AGEMA_signal_1251,
         SubCellInst_SboxInst_14_XX_1_, new_AGEMA_signal_1253,
         SubCellInst_SboxInst_14_XX_2_, new_AGEMA_signal_1537,
         SubCellInst_SboxInst_14_Q0, new_AGEMA_signal_1538,
         SubCellInst_SboxInst_14_Q1, new_AGEMA_signal_1539,
         SubCellInst_SboxInst_14_Q4, new_AGEMA_signal_1540,
         SubCellInst_SboxInst_14_Q6, new_AGEMA_signal_1592,
         SubCellInst_SboxInst_14_L1, new_AGEMA_signal_1541,
         SubCellInst_SboxInst_14_L2, SubCellInst_SboxInst_15_n3,
         new_AGEMA_signal_1257, SubCellInst_SboxInst_15_XX_1_,
         new_AGEMA_signal_1259, SubCellInst_SboxInst_15_XX_2_,
         new_AGEMA_signal_1543, SubCellInst_SboxInst_15_Q0,
         new_AGEMA_signal_1544, SubCellInst_SboxInst_15_Q1,
         new_AGEMA_signal_1545, SubCellInst_SboxInst_15_Q4,
         new_AGEMA_signal_1546, SubCellInst_SboxInst_15_Q6,
         new_AGEMA_signal_1595, SubCellInst_SboxInst_15_L1,
         new_AGEMA_signal_1547, SubCellInst_SboxInst_15_L2,
         new_AGEMA_signal_1262, new_AGEMA_signal_1260, new_AGEMA_signal_1265,
         new_AGEMA_signal_1263, new_AGEMA_signal_1268, new_AGEMA_signal_1266,
         new_AGEMA_signal_1271, new_AGEMA_signal_1269, new_AGEMA_signal_1274,
         new_AGEMA_signal_1272, new_AGEMA_signal_1277, new_AGEMA_signal_1275,
         new_AGEMA_signal_1280, new_AGEMA_signal_1278, new_AGEMA_signal_1283,
         new_AGEMA_signal_1281, new_AGEMA_signal_1286, new_AGEMA_signal_1284,
         new_AGEMA_signal_1289, new_AGEMA_signal_1287, new_AGEMA_signal_1292,
         new_AGEMA_signal_1290, new_AGEMA_signal_1295, new_AGEMA_signal_1293,
         new_AGEMA_signal_1298, new_AGEMA_signal_1296, new_AGEMA_signal_1301,
         new_AGEMA_signal_1299, new_AGEMA_signal_1304, new_AGEMA_signal_1302,
         new_AGEMA_signal_1307, new_AGEMA_signal_1305, new_AGEMA_signal_1310,
         new_AGEMA_signal_1308, new_AGEMA_signal_1313, new_AGEMA_signal_1311,
         new_AGEMA_signal_1316, new_AGEMA_signal_1314, new_AGEMA_signal_1319,
         new_AGEMA_signal_1317, new_AGEMA_signal_1322, new_AGEMA_signal_1320,
         new_AGEMA_signal_1325, new_AGEMA_signal_1323, new_AGEMA_signal_1328,
         new_AGEMA_signal_1326, new_AGEMA_signal_1331, new_AGEMA_signal_1329,
         new_AGEMA_signal_1334, new_AGEMA_signal_1332, new_AGEMA_signal_1337,
         new_AGEMA_signal_1335, new_AGEMA_signal_1340, new_AGEMA_signal_1338,
         new_AGEMA_signal_1343, new_AGEMA_signal_1341, new_AGEMA_signal_1346,
         new_AGEMA_signal_1344, new_AGEMA_signal_1349, new_AGEMA_signal_1347,
         new_AGEMA_signal_1352, new_AGEMA_signal_1350, new_AGEMA_signal_1355,
         new_AGEMA_signal_1353, new_AGEMA_signal_1358, new_AGEMA_signal_1356,
         new_AGEMA_signal_1361, new_AGEMA_signal_1359, new_AGEMA_signal_1364,
         new_AGEMA_signal_1362, new_AGEMA_signal_1367, new_AGEMA_signal_1365,
         new_AGEMA_signal_1370, new_AGEMA_signal_1368, new_AGEMA_signal_1373,
         new_AGEMA_signal_1371, new_AGEMA_signal_1376, new_AGEMA_signal_1374,
         new_AGEMA_signal_1379, new_AGEMA_signal_1377, new_AGEMA_signal_1382,
         new_AGEMA_signal_1380, new_AGEMA_signal_1385, new_AGEMA_signal_1383,
         new_AGEMA_signal_1388, new_AGEMA_signal_1386, new_AGEMA_signal_1391,
         new_AGEMA_signal_1389, new_AGEMA_signal_1394, new_AGEMA_signal_1392,
         new_AGEMA_signal_1397, new_AGEMA_signal_1395, new_AGEMA_signal_1400,
         new_AGEMA_signal_1398, new_AGEMA_signal_1403, new_AGEMA_signal_1401,
         new_AGEMA_signal_1406, new_AGEMA_signal_1404, new_AGEMA_signal_1409,
         new_AGEMA_signal_1407, new_AGEMA_signal_1412, new_AGEMA_signal_1410,
         new_AGEMA_signal_1415, new_AGEMA_signal_1413, new_AGEMA_signal_1418,
         new_AGEMA_signal_1416, new_AGEMA_signal_1421, new_AGEMA_signal_1419,
         new_AGEMA_signal_1424, new_AGEMA_signal_1422, new_AGEMA_signal_1427,
         new_AGEMA_signal_1425, new_AGEMA_signal_1430, new_AGEMA_signal_1428,
         new_AGEMA_signal_1433, new_AGEMA_signal_1431, new_AGEMA_signal_1436,
         new_AGEMA_signal_1434, new_AGEMA_signal_1439, new_AGEMA_signal_1437,
         new_AGEMA_signal_1442, new_AGEMA_signal_1440, new_AGEMA_signal_1445,
         new_AGEMA_signal_1443, new_AGEMA_signal_1448, new_AGEMA_signal_1446,
         new_AGEMA_signal_1451, new_AGEMA_signal_1449, FSM_1, clk_gated,
         new_AGEMA_signal_1922, new_AGEMA_signal_1915, new_AGEMA_signal_1982,
         new_AGEMA_signal_1975, new_AGEMA_signal_1924, new_AGEMA_signal_1917,
         new_AGEMA_signal_1984, new_AGEMA_signal_1977, new_AGEMA_signal_1926,
         new_AGEMA_signal_1919, new_AGEMA_signal_1986, new_AGEMA_signal_1979,
         new_AGEMA_signal_2042, new_AGEMA_signal_2033, new_AGEMA_signal_2085,
         new_AGEMA_signal_2077, new_AGEMA_signal_1928, new_AGEMA_signal_1909,
         new_AGEMA_signal_1988, new_AGEMA_signal_1968, new_AGEMA_signal_1930,
         new_AGEMA_signal_1911, new_AGEMA_signal_1990, new_AGEMA_signal_1970,
         new_AGEMA_signal_2048, new_AGEMA_signal_2023, new_AGEMA_signal_2091,
         new_AGEMA_signal_2071, new_AGEMA_signal_1932, new_AGEMA_signal_1913,
         new_AGEMA_signal_1992, new_AGEMA_signal_1973, new_AGEMA_signal_1821,
         new_AGEMA_signal_1810, new_AGEMA_signal_1874, new_AGEMA_signal_1854,
         new_AGEMA_signal_1823, new_AGEMA_signal_1812, new_AGEMA_signal_1876,
         new_AGEMA_signal_1856, new_AGEMA_signal_1825, new_AGEMA_signal_1814,
         new_AGEMA_signal_1878, new_AGEMA_signal_1858, new_AGEMA_signal_1940,
         new_AGEMA_signal_1898, new_AGEMA_signal_2000, new_AGEMA_signal_1958,
         new_AGEMA_signal_1942, new_AGEMA_signal_1901, new_AGEMA_signal_2002,
         new_AGEMA_signal_1960, new_AGEMA_signal_1944, new_AGEMA_signal_1903,
         new_AGEMA_signal_2004, new_AGEMA_signal_1963, new_AGEMA_signal_1946,
         new_AGEMA_signal_1906, new_AGEMA_signal_2006, new_AGEMA_signal_1965,
         new_AGEMA_signal_2060, new_AGEMA_signal_2017, new_AGEMA_signal_2103,
         new_AGEMA_signal_2067, new_AGEMA_signal_1724,
         SubCellInst_SboxInst_0_YY_1_, new_AGEMA_signal_1660,
         SubCellInst_SboxInst_0_YY_0_, new_AGEMA_signal_1548,
         SubCellInst_SboxInst_0_T0, new_AGEMA_signal_1596,
         SubCellInst_SboxInst_0_Q2, new_AGEMA_signal_1549,
         SubCellInst_SboxInst_0_T2, new_AGEMA_signal_1597,
         SubCellInst_SboxInst_0_Q7, new_AGEMA_signal_1598,
         SubCellInst_SboxInst_0_L3, new_AGEMA_signal_1726,
         SubCellInst_SboxInst_1_YY_1_, new_AGEMA_signal_1664,
         SubCellInst_SboxInst_1_YY_0_, new_AGEMA_signal_1551,
         SubCellInst_SboxInst_1_T0, new_AGEMA_signal_1600,
         SubCellInst_SboxInst_1_Q2, new_AGEMA_signal_1552,
         SubCellInst_SboxInst_1_T2, new_AGEMA_signal_1601,
         SubCellInst_SboxInst_1_Q7, new_AGEMA_signal_1602,
         SubCellInst_SboxInst_1_L3, new_AGEMA_signal_1728,
         SubCellInst_SboxInst_2_YY_1_, new_AGEMA_signal_1668,
         SubCellInst_SboxInst_2_YY_0_, new_AGEMA_signal_1554,
         SubCellInst_SboxInst_2_T0, new_AGEMA_signal_1604,
         SubCellInst_SboxInst_2_Q2, new_AGEMA_signal_1555,
         SubCellInst_SboxInst_2_T2, new_AGEMA_signal_1605,
         SubCellInst_SboxInst_2_Q7, new_AGEMA_signal_1606,
         SubCellInst_SboxInst_2_L3, new_AGEMA_signal_1730,
         SubCellInst_SboxInst_3_YY_1_, new_AGEMA_signal_1672,
         SubCellInst_SboxInst_3_YY_0_, new_AGEMA_signal_1557,
         SubCellInst_SboxInst_3_T0, new_AGEMA_signal_1608,
         SubCellInst_SboxInst_3_Q2, new_AGEMA_signal_1558,
         SubCellInst_SboxInst_3_T2, new_AGEMA_signal_1609,
         SubCellInst_SboxInst_3_Q7, new_AGEMA_signal_1610,
         SubCellInst_SboxInst_3_L3, new_AGEMA_signal_1732,
         SubCellInst_SboxInst_4_YY_1_, new_AGEMA_signal_1676,
         SubCellInst_SboxInst_4_YY_0_, new_AGEMA_signal_1560,
         SubCellInst_SboxInst_4_T0, new_AGEMA_signal_1612,
         SubCellInst_SboxInst_4_Q2, new_AGEMA_signal_1561,
         SubCellInst_SboxInst_4_T2, new_AGEMA_signal_1613,
         SubCellInst_SboxInst_4_Q7, new_AGEMA_signal_1614,
         SubCellInst_SboxInst_4_L3, new_AGEMA_signal_1734,
         SubCellInst_SboxInst_5_YY_1_, new_AGEMA_signal_1680,
         SubCellInst_SboxInst_5_YY_0_, new_AGEMA_signal_1563,
         SubCellInst_SboxInst_5_T0, new_AGEMA_signal_1616,
         SubCellInst_SboxInst_5_Q2, new_AGEMA_signal_1564,
         SubCellInst_SboxInst_5_T2, new_AGEMA_signal_1617,
         SubCellInst_SboxInst_5_Q7, new_AGEMA_signal_1618,
         SubCellInst_SboxInst_5_L3, new_AGEMA_signal_1736,
         SubCellInst_SboxInst_6_YY_1_, new_AGEMA_signal_1684,
         SubCellInst_SboxInst_6_YY_0_, new_AGEMA_signal_1566,
         SubCellInst_SboxInst_6_T0, new_AGEMA_signal_1620,
         SubCellInst_SboxInst_6_Q2, new_AGEMA_signal_1567,
         SubCellInst_SboxInst_6_T2, new_AGEMA_signal_1621,
         SubCellInst_SboxInst_6_Q7, new_AGEMA_signal_1622,
         SubCellInst_SboxInst_6_L3, new_AGEMA_signal_1738,
         SubCellInst_SboxInst_7_YY_1_, new_AGEMA_signal_1688,
         SubCellInst_SboxInst_7_YY_0_, new_AGEMA_signal_1569,
         SubCellInst_SboxInst_7_T0, new_AGEMA_signal_1624,
         SubCellInst_SboxInst_7_Q2, new_AGEMA_signal_1570,
         SubCellInst_SboxInst_7_T2, new_AGEMA_signal_1625,
         SubCellInst_SboxInst_7_Q7, new_AGEMA_signal_1626,
         SubCellInst_SboxInst_7_L3, new_AGEMA_signal_1740,
         SubCellInst_SboxInst_8_YY_1_, new_AGEMA_signal_1692,
         SubCellInst_SboxInst_8_YY_0_, new_AGEMA_signal_1572,
         SubCellInst_SboxInst_8_T0, new_AGEMA_signal_1628,
         SubCellInst_SboxInst_8_Q2, new_AGEMA_signal_1573,
         SubCellInst_SboxInst_8_T2, new_AGEMA_signal_1629,
         SubCellInst_SboxInst_8_Q7, new_AGEMA_signal_1630,
         SubCellInst_SboxInst_8_L3, new_AGEMA_signal_1742,
         SubCellInst_SboxInst_9_YY_1_, new_AGEMA_signal_1696,
         SubCellInst_SboxInst_9_YY_0_, new_AGEMA_signal_1575,
         SubCellInst_SboxInst_9_T0, new_AGEMA_signal_1632,
         SubCellInst_SboxInst_9_Q2, new_AGEMA_signal_1576,
         SubCellInst_SboxInst_9_T2, new_AGEMA_signal_1633,
         SubCellInst_SboxInst_9_Q7, new_AGEMA_signal_1634,
         SubCellInst_SboxInst_9_L3, new_AGEMA_signal_1744,
         SubCellInst_SboxInst_10_YY_1_, new_AGEMA_signal_1700,
         SubCellInst_SboxInst_10_YY_0_, new_AGEMA_signal_1578,
         SubCellInst_SboxInst_10_T0, new_AGEMA_signal_1636,
         SubCellInst_SboxInst_10_Q2, new_AGEMA_signal_1579,
         SubCellInst_SboxInst_10_T2, new_AGEMA_signal_1637,
         SubCellInst_SboxInst_10_Q7, new_AGEMA_signal_1638,
         SubCellInst_SboxInst_10_L3, SubCellOutput_47, SubCellOutput_46,
         SubCellOutput_45, SubCellOutput_44, SubCellOutput_29,
         new_AGEMA_signal_1746, SubCellInst_SboxInst_11_YY_1_,
         new_AGEMA_signal_1704, SubCellInst_SboxInst_11_YY_0_,
         new_AGEMA_signal_1581, SubCellInst_SboxInst_11_T0,
         new_AGEMA_signal_1640, SubCellInst_SboxInst_11_Q2,
         new_AGEMA_signal_1582, SubCellInst_SboxInst_11_T2,
         new_AGEMA_signal_1641, SubCellInst_SboxInst_11_Q7,
         new_AGEMA_signal_1642, SubCellInst_SboxInst_11_L3,
         new_AGEMA_signal_1748, SubCellInst_SboxInst_12_YY_1_,
         new_AGEMA_signal_1708, SubCellInst_SboxInst_12_YY_0_,
         new_AGEMA_signal_1584, SubCellInst_SboxInst_12_T0,
         new_AGEMA_signal_1644, SubCellInst_SboxInst_12_Q2,
         new_AGEMA_signal_1585, SubCellInst_SboxInst_12_T2,
         new_AGEMA_signal_1645, SubCellInst_SboxInst_12_Q7,
         new_AGEMA_signal_1646, SubCellInst_SboxInst_12_L3,
         new_AGEMA_signal_1750, SubCellInst_SboxInst_13_YY_1_,
         new_AGEMA_signal_1712, SubCellInst_SboxInst_13_YY_0_,
         new_AGEMA_signal_1587, SubCellInst_SboxInst_13_T0,
         new_AGEMA_signal_1648, SubCellInst_SboxInst_13_Q2,
         new_AGEMA_signal_1588, SubCellInst_SboxInst_13_T2,
         new_AGEMA_signal_1649, SubCellInst_SboxInst_13_Q7,
         new_AGEMA_signal_1650, SubCellInst_SboxInst_13_L3,
         new_AGEMA_signal_1752, SubCellInst_SboxInst_14_YY_1_,
         new_AGEMA_signal_1716, SubCellInst_SboxInst_14_YY_0_,
         new_AGEMA_signal_1590, SubCellInst_SboxInst_14_T0,
         new_AGEMA_signal_1652, SubCellInst_SboxInst_14_Q2,
         new_AGEMA_signal_1591, SubCellInst_SboxInst_14_T2,
         new_AGEMA_signal_1653, SubCellInst_SboxInst_14_Q7,
         new_AGEMA_signal_1654, SubCellInst_SboxInst_14_L3,
         new_AGEMA_signal_1754, SubCellInst_SboxInst_15_YY_1_,
         new_AGEMA_signal_1720, SubCellInst_SboxInst_15_YY_0_,
         new_AGEMA_signal_1593, SubCellInst_SboxInst_15_T0,
         new_AGEMA_signal_1656, SubCellInst_SboxInst_15_Q2,
         new_AGEMA_signal_1594, SubCellInst_SboxInst_15_T2,
         new_AGEMA_signal_1657, SubCellInst_SboxInst_15_Q7,
         new_AGEMA_signal_1658, SubCellInst_SboxInst_15_L3,
         new_AGEMA_signal_1800, new_AGEMA_signal_1756,
         AddConstXOR_AddConstXOR_XORInst_0_2_n1, new_AGEMA_signal_1843,
         new_AGEMA_signal_1801, AddConstXOR_AddConstXOR_XORInst_0_3_n1,
         new_AGEMA_signal_1802, new_AGEMA_signal_1757,
         AddConstXOR_AddConstXOR_XORInst_1_2_n1, new_AGEMA_signal_1845,
         new_AGEMA_signal_1803, AddConstXOR_AddConstXOR_XORInst_1_3_n1,
         new_AGEMA_signal_1804, new_AGEMA_signal_1758,
         AddRoundTweakeyXOR_XORInst_0_2_n1, new_AGEMA_signal_1847,
         new_AGEMA_signal_1805, AddRoundTweakeyXOR_XORInst_0_3_n1,
         new_AGEMA_signal_1806, new_AGEMA_signal_1759,
         AddRoundTweakeyXOR_XORInst_1_2_n1, new_AGEMA_signal_1849,
         new_AGEMA_signal_1807, AddRoundTweakeyXOR_XORInst_1_3_n1,
         new_AGEMA_signal_1808, new_AGEMA_signal_1760,
         AddRoundTweakeyXOR_XORInst_2_2_n1, new_AGEMA_signal_1851,
         new_AGEMA_signal_1809, AddRoundTweakeyXOR_XORInst_2_3_n1,
         new_AGEMA_signal_1890, new_AGEMA_signal_1852,
         AddRoundTweakeyXOR_XORInst_3_2_n1, new_AGEMA_signal_1953,
         new_AGEMA_signal_1891, AddRoundTweakeyXOR_XORInst_3_3_n1,
         new_AGEMA_signal_1761, AddRoundTweakeyXOR_XORInst_4_2_n1,
         new_AGEMA_signal_1811, AddRoundTweakeyXOR_XORInst_4_3_n1,
         new_AGEMA_signal_1762, AddRoundTweakeyXOR_XORInst_5_2_n1,
         new_AGEMA_signal_1813, AddRoundTweakeyXOR_XORInst_5_3_n1,
         new_AGEMA_signal_1763, AddRoundTweakeyXOR_XORInst_6_2_n1,
         new_AGEMA_signal_1815, AddRoundTweakeyXOR_XORInst_6_3_n1,
         new_AGEMA_signal_1859, AddRoundTweakeyXOR_XORInst_7_2_n1,
         new_AGEMA_signal_1899, AddRoundTweakeyXOR_XORInst_7_3_n1,
         new_AGEMA_signal_1764, MCInst_MCR0_XORInst_0_2_n1,
         new_AGEMA_signal_1861, MCInst_MCR0_XORInst_0_2_n2,
         new_AGEMA_signal_1816, MCInst_MCR0_XORInst_0_3_n1,
         new_AGEMA_signal_1902, MCInst_MCR0_XORInst_0_3_n2,
         new_AGEMA_signal_1765, MCInst_MCR0_XORInst_1_2_n1,
         new_AGEMA_signal_1863, MCInst_MCR0_XORInst_1_2_n2,
         new_AGEMA_signal_1817, MCInst_MCR0_XORInst_1_3_n1,
         new_AGEMA_signal_1904, MCInst_MCR0_XORInst_1_3_n2,
         new_AGEMA_signal_1766, MCInst_MCR0_XORInst_2_2_n1,
         new_AGEMA_signal_1865, MCInst_MCR0_XORInst_2_2_n2,
         new_AGEMA_signal_1818, MCInst_MCR0_XORInst_2_3_n1,
         new_AGEMA_signal_1907, MCInst_MCR0_XORInst_2_3_n2,
         new_AGEMA_signal_1767, MCInst_MCR0_XORInst_3_2_n1,
         new_AGEMA_signal_1966, MCInst_MCR0_XORInst_3_2_n2,
         new_AGEMA_signal_1819, MCInst_MCR0_XORInst_3_3_n1,
         new_AGEMA_signal_2018, MCInst_MCR0_XORInst_3_3_n2,
         new_AGEMA_signal_1867, MCInst_MCR2_XORInst_0_2_n1,
         new_AGEMA_signal_1910, MCInst_MCR2_XORInst_0_3_n1,
         new_AGEMA_signal_1868, MCInst_MCR2_XORInst_1_2_n1,
         new_AGEMA_signal_1912, MCInst_MCR2_XORInst_1_3_n1,
         new_AGEMA_signal_1971, MCInst_MCR2_XORInst_2_2_n1,
         new_AGEMA_signal_2024, MCInst_MCR2_XORInst_2_3_n1,
         new_AGEMA_signal_1869, MCInst_MCR2_XORInst_3_2_n1,
         new_AGEMA_signal_1914, MCInst_MCR2_XORInst_3_3_n1,
         new_AGEMA_signal_1870, MCInst_MCR3_XORInst_0_2_n1,
         new_AGEMA_signal_1916, MCInst_MCR3_XORInst_0_3_n1,
         new_AGEMA_signal_1871, MCInst_MCR3_XORInst_1_2_n1,
         new_AGEMA_signal_1918, MCInst_MCR3_XORInst_1_3_n1,
         new_AGEMA_signal_1872, MCInst_MCR3_XORInst_2_2_n1,
         new_AGEMA_signal_1920, MCInst_MCR3_XORInst_2_3_n1,
         new_AGEMA_signal_1980, MCInst_MCR3_XORInst_3_2_n1,
         new_AGEMA_signal_2034, MCInst_MCR3_XORInst_3_3_n1,
         new_AGEMA_signal_2036, new_AGEMA_signal_2027, new_AGEMA_signal_2079,
         new_AGEMA_signal_2073, new_AGEMA_signal_2038, new_AGEMA_signal_2029,
         new_AGEMA_signal_2081, new_AGEMA_signal_2074, new_AGEMA_signal_2040,
         new_AGEMA_signal_2031, new_AGEMA_signal_2083, new_AGEMA_signal_2075,
         new_AGEMA_signal_2111, new_AGEMA_signal_2108, new_AGEMA_signal_2120,
         new_AGEMA_signal_2118, new_AGEMA_signal_2044, new_AGEMA_signal_2019,
         new_AGEMA_signal_2087, new_AGEMA_signal_2068, new_AGEMA_signal_2046,
         new_AGEMA_signal_2021, new_AGEMA_signal_2089, new_AGEMA_signal_2069,
         new_AGEMA_signal_2113, new_AGEMA_signal_2106, new_AGEMA_signal_2122,
         new_AGEMA_signal_2117, new_AGEMA_signal_2050, new_AGEMA_signal_2025,
         new_AGEMA_signal_2093, new_AGEMA_signal_2072, new_AGEMA_signal_1934,
         new_AGEMA_signal_1892, new_AGEMA_signal_1994, new_AGEMA_signal_1954,
         new_AGEMA_signal_1936, new_AGEMA_signal_1894, new_AGEMA_signal_1996,
         new_AGEMA_signal_1955, new_AGEMA_signal_1938, new_AGEMA_signal_1896,
         new_AGEMA_signal_1998, new_AGEMA_signal_1956, new_AGEMA_signal_2052,
         new_AGEMA_signal_2009, new_AGEMA_signal_2095, new_AGEMA_signal_2062,
         new_AGEMA_signal_2054, new_AGEMA_signal_2011, new_AGEMA_signal_2097,
         new_AGEMA_signal_2063, new_AGEMA_signal_2056, new_AGEMA_signal_2013,
         new_AGEMA_signal_2099, new_AGEMA_signal_2064, new_AGEMA_signal_2058,
         new_AGEMA_signal_2015, new_AGEMA_signal_2101, new_AGEMA_signal_2065,
         new_AGEMA_signal_2115, new_AGEMA_signal_2104, new_AGEMA_signal_2124,
         new_AGEMA_signal_2116, new_AGEMA_signal_1661,
         SubCellInst_SboxInst_0_T1, new_AGEMA_signal_1725,
         SubCellInst_SboxInst_0_L0, new_AGEMA_signal_1662,
         SubCellInst_SboxInst_0_T3, new_AGEMA_signal_1768,
         SubCellInst_SboxInst_0_YY_3, new_AGEMA_signal_1769,
         new_AGEMA_signal_1826, new_AGEMA_signal_1665,
         SubCellInst_SboxInst_1_T1, new_AGEMA_signal_1727,
         SubCellInst_SboxInst_1_L0, new_AGEMA_signal_1666,
         SubCellInst_SboxInst_1_T3, new_AGEMA_signal_1770,
         SubCellInst_SboxInst_1_YY_3, new_AGEMA_signal_1771,
         new_AGEMA_signal_1827, new_AGEMA_signal_1669,
         SubCellInst_SboxInst_2_T1, new_AGEMA_signal_1729,
         SubCellInst_SboxInst_2_L0, new_AGEMA_signal_1670,
         SubCellInst_SboxInst_2_T3, new_AGEMA_signal_1772,
         SubCellInst_SboxInst_2_YY_3, new_AGEMA_signal_1773,
         new_AGEMA_signal_1828, new_AGEMA_signal_1673,
         SubCellInst_SboxInst_3_T1, new_AGEMA_signal_1731,
         SubCellInst_SboxInst_3_L0, new_AGEMA_signal_1674,
         SubCellInst_SboxInst_3_T3, new_AGEMA_signal_1774,
         SubCellInst_SboxInst_3_YY_3, new_AGEMA_signal_1775,
         new_AGEMA_signal_1829, new_AGEMA_signal_1677,
         SubCellInst_SboxInst_4_T1, new_AGEMA_signal_1733,
         SubCellInst_SboxInst_4_L0, new_AGEMA_signal_1678,
         SubCellInst_SboxInst_4_T3, new_AGEMA_signal_1776,
         SubCellInst_SboxInst_4_YY_3, new_AGEMA_signal_1777,
         new_AGEMA_signal_1830, new_AGEMA_signal_1681,
         SubCellInst_SboxInst_5_T1, new_AGEMA_signal_1735,
         SubCellInst_SboxInst_5_L0, new_AGEMA_signal_1682,
         SubCellInst_SboxInst_5_T3, new_AGEMA_signal_1778,
         SubCellInst_SboxInst_5_YY_3, new_AGEMA_signal_1779,
         new_AGEMA_signal_1831, new_AGEMA_signal_1685,
         SubCellInst_SboxInst_6_T1, new_AGEMA_signal_1737,
         SubCellInst_SboxInst_6_L0, new_AGEMA_signal_1686,
         SubCellInst_SboxInst_6_T3, new_AGEMA_signal_1780,
         SubCellInst_SboxInst_6_YY_3, new_AGEMA_signal_1781,
         new_AGEMA_signal_1832, new_AGEMA_signal_1689,
         SubCellInst_SboxInst_7_T1, new_AGEMA_signal_1739,
         SubCellInst_SboxInst_7_L0, new_AGEMA_signal_1690,
         SubCellInst_SboxInst_7_T3, new_AGEMA_signal_1782,
         SubCellInst_SboxInst_7_YY_3, new_AGEMA_signal_1783,
         new_AGEMA_signal_1693, SubCellInst_SboxInst_8_T1,
         new_AGEMA_signal_1741, SubCellInst_SboxInst_8_L0,
         new_AGEMA_signal_1694, SubCellInst_SboxInst_8_T3,
         new_AGEMA_signal_1784, SubCellInst_SboxInst_8_YY_3,
         new_AGEMA_signal_1785, new_AGEMA_signal_1834, new_AGEMA_signal_1697,
         SubCellInst_SboxInst_9_T1, new_AGEMA_signal_1743,
         SubCellInst_SboxInst_9_L0, new_AGEMA_signal_1698,
         SubCellInst_SboxInst_9_T3, new_AGEMA_signal_1786,
         SubCellInst_SboxInst_9_YY_3, new_AGEMA_signal_1787,
         new_AGEMA_signal_1835, new_AGEMA_signal_1701,
         SubCellInst_SboxInst_10_T1, new_AGEMA_signal_1745,
         SubCellInst_SboxInst_10_L0, new_AGEMA_signal_1702,
         SubCellInst_SboxInst_10_T3, new_AGEMA_signal_1788,
         SubCellInst_SboxInst_10_YY_3, new_AGEMA_signal_1789,
         new_AGEMA_signal_1836, new_AGEMA_signal_1705,
         SubCellInst_SboxInst_11_T1, new_AGEMA_signal_1747,
         SubCellInst_SboxInst_11_L0, new_AGEMA_signal_1706,
         SubCellInst_SboxInst_11_T3, new_AGEMA_signal_1790,
         SubCellInst_SboxInst_11_YY_3, new_AGEMA_signal_1791,
         new_AGEMA_signal_1837, new_AGEMA_signal_1709,
         SubCellInst_SboxInst_12_T1, new_AGEMA_signal_1749,
         SubCellInst_SboxInst_12_L0, new_AGEMA_signal_1710,
         SubCellInst_SboxInst_12_T3, new_AGEMA_signal_1792,
         SubCellInst_SboxInst_12_YY_3, new_AGEMA_signal_1793,
         new_AGEMA_signal_1838, new_AGEMA_signal_1713,
         SubCellInst_SboxInst_13_T1, new_AGEMA_signal_1751,
         SubCellInst_SboxInst_13_L0, new_AGEMA_signal_1714,
         SubCellInst_SboxInst_13_T3, new_AGEMA_signal_1794,
         SubCellInst_SboxInst_13_YY_3, new_AGEMA_signal_1795,
         new_AGEMA_signal_1839, new_AGEMA_signal_1717,
         SubCellInst_SboxInst_14_T1, new_AGEMA_signal_1753,
         SubCellInst_SboxInst_14_L0, new_AGEMA_signal_1718,
         SubCellInst_SboxInst_14_T3, new_AGEMA_signal_1796,
         SubCellInst_SboxInst_14_YY_3, new_AGEMA_signal_1797,
         new_AGEMA_signal_1840, new_AGEMA_signal_1721,
         SubCellInst_SboxInst_15_T1, new_AGEMA_signal_1755,
         SubCellInst_SboxInst_15_L0, new_AGEMA_signal_1722,
         SubCellInst_SboxInst_15_T3, new_AGEMA_signal_1798,
         SubCellInst_SboxInst_15_YY_3, new_AGEMA_signal_1799,
         new_AGEMA_signal_1841, new_AGEMA_signal_1879, new_AGEMA_signal_1880,
         new_AGEMA_signal_1842, AddConstXOR_AddConstXOR_XORInst_0_0_n1,
         new_AGEMA_signal_1947, new_AGEMA_signal_1881,
         AddConstXOR_AddConstXOR_XORInst_0_1_n1, new_AGEMA_signal_1882,
         new_AGEMA_signal_1844, AddConstXOR_AddConstXOR_XORInst_1_0_n1,
         new_AGEMA_signal_1948, new_AGEMA_signal_1883,
         AddConstXOR_AddConstXOR_XORInst_1_1_n1, new_AGEMA_signal_1884,
         new_AGEMA_signal_1846, AddRoundTweakeyXOR_XORInst_0_0_n1,
         new_AGEMA_signal_1949, new_AGEMA_signal_1885,
         AddRoundTweakeyXOR_XORInst_0_1_n1, new_AGEMA_signal_1886,
         new_AGEMA_signal_1848, AddRoundTweakeyXOR_XORInst_1_0_n1,
         new_AGEMA_signal_1950, new_AGEMA_signal_1887,
         AddRoundTweakeyXOR_XORInst_1_1_n1, new_AGEMA_signal_1888,
         new_AGEMA_signal_1850, AddRoundTweakeyXOR_XORInst_2_0_n1,
         new_AGEMA_signal_1951, new_AGEMA_signal_1889,
         AddRoundTweakeyXOR_XORInst_2_1_n1, new_AGEMA_signal_2007,
         new_AGEMA_signal_1952, AddRoundTweakeyXOR_XORInst_3_0_n1,
         new_AGEMA_signal_2061, new_AGEMA_signal_2008,
         AddRoundTweakeyXOR_XORInst_3_1_n1, new_AGEMA_signal_1853,
         AddRoundTweakeyXOR_XORInst_4_0_n1, new_AGEMA_signal_1893,
         AddRoundTweakeyXOR_XORInst_4_1_n1, new_AGEMA_signal_1855,
         AddRoundTweakeyXOR_XORInst_5_0_n1, new_AGEMA_signal_1895,
         AddRoundTweakeyXOR_XORInst_5_1_n1, new_AGEMA_signal_1857,
         AddRoundTweakeyXOR_XORInst_6_0_n1, new_AGEMA_signal_1897,
         AddRoundTweakeyXOR_XORInst_6_1_n1, new_AGEMA_signal_1957,
         AddRoundTweakeyXOR_XORInst_7_0_n1, new_AGEMA_signal_2010,
         AddRoundTweakeyXOR_XORInst_7_1_n1, new_AGEMA_signal_1860,
         MCInst_MCR0_XORInst_0_0_n1, new_AGEMA_signal_1959,
         MCInst_MCR0_XORInst_0_0_n2, new_AGEMA_signal_1900,
         MCInst_MCR0_XORInst_0_1_n1, new_AGEMA_signal_2012,
         MCInst_MCR0_XORInst_0_1_n2, new_AGEMA_signal_1862,
         MCInst_MCR0_XORInst_1_0_n1, new_AGEMA_signal_1961,
         MCInst_MCR0_XORInst_1_0_n2, new_AGEMA_signal_1962,
         MCInst_MCR0_XORInst_1_1_n1, new_AGEMA_signal_2014,
         MCInst_MCR0_XORInst_1_1_n2, new_AGEMA_signal_1864,
         MCInst_MCR0_XORInst_2_0_n1, new_AGEMA_signal_1964,
         MCInst_MCR0_XORInst_2_0_n2, new_AGEMA_signal_1905,
         MCInst_MCR0_XORInst_2_1_n1, new_AGEMA_signal_2016,
         MCInst_MCR0_XORInst_2_1_n2, new_AGEMA_signal_1866,
         MCInst_MCR0_XORInst_3_0_n1, new_AGEMA_signal_2066,
         MCInst_MCR0_XORInst_3_0_n2, new_AGEMA_signal_1908,
         MCInst_MCR0_XORInst_3_1_n1, new_AGEMA_signal_2105,
         MCInst_MCR0_XORInst_3_1_n2, new_AGEMA_signal_1967,
         MCInst_MCR2_XORInst_0_0_n1, new_AGEMA_signal_2020,
         MCInst_MCR2_XORInst_0_1_n1, new_AGEMA_signal_1969,
         MCInst_MCR2_XORInst_1_0_n1, new_AGEMA_signal_2022,
         MCInst_MCR2_XORInst_1_1_n1, new_AGEMA_signal_2070,
         MCInst_MCR2_XORInst_2_0_n1, new_AGEMA_signal_2107,
         MCInst_MCR2_XORInst_2_1_n1, new_AGEMA_signal_1972,
         MCInst_MCR2_XORInst_3_0_n1, new_AGEMA_signal_2026,
         MCInst_MCR2_XORInst_3_1_n1, new_AGEMA_signal_1974,
         MCInst_MCR3_XORInst_0_0_n1, new_AGEMA_signal_2028,
         MCInst_MCR3_XORInst_0_1_n1, new_AGEMA_signal_1976,
         MCInst_MCR3_XORInst_1_0_n1, new_AGEMA_signal_2030,
         MCInst_MCR3_XORInst_1_1_n1, new_AGEMA_signal_1978,
         MCInst_MCR3_XORInst_2_0_n1, new_AGEMA_signal_2032,
         MCInst_MCR3_XORInst_2_1_n1, new_AGEMA_signal_2076,
         MCInst_MCR3_XORInst_3_0_n1, new_AGEMA_signal_2109,
         MCInst_MCR3_XORInst_3_1_n1, n13, n14, n15, n16, n17, n18, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, ClockGatingInst_n11,
         ClockGatingInst_n10, ClockGatingInst_n9, ClockGatingInst_n8,
         ClockGatingInst_n7, ClockGatingInst_n6, ClockGatingInst_n4,
         ClockGatingInst_n3, ClockGatingInst_n2, ClockGatingInst_n1,
         ClockGatingInst_LatchedEnable, ClockGatingInst_N7,
         ClockGatingInst_ShiftRegister_5_, SubCellInst_SboxInst_0_AND1_U1_n9,
         SubCellInst_SboxInst_0_AND1_U1_n8, SubCellInst_SboxInst_0_AND1_U1_n7,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_0_AND3_U1_n9, SubCellInst_SboxInst_0_AND3_U1_n8,
         SubCellInst_SboxInst_0_AND3_U1_n7,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND1_U1_n9, SubCellInst_SboxInst_1_AND1_U1_n8,
         SubCellInst_SboxInst_1_AND1_U1_n7,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND3_U1_n9, SubCellInst_SboxInst_1_AND3_U1_n8,
         SubCellInst_SboxInst_1_AND3_U1_n7,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND1_U1_n9, SubCellInst_SboxInst_2_AND1_U1_n8,
         SubCellInst_SboxInst_2_AND1_U1_n7,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND3_U1_n9, SubCellInst_SboxInst_2_AND3_U1_n8,
         SubCellInst_SboxInst_2_AND3_U1_n7,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND1_U1_n9, SubCellInst_SboxInst_3_AND1_U1_n8,
         SubCellInst_SboxInst_3_AND1_U1_n7,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND3_U1_n9, SubCellInst_SboxInst_3_AND3_U1_n8,
         SubCellInst_SboxInst_3_AND3_U1_n7,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND1_U1_n9, SubCellInst_SboxInst_4_AND1_U1_n8,
         SubCellInst_SboxInst_4_AND1_U1_n7,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND3_U1_n9, SubCellInst_SboxInst_4_AND3_U1_n8,
         SubCellInst_SboxInst_4_AND3_U1_n7,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND1_U1_n9, SubCellInst_SboxInst_5_AND1_U1_n8,
         SubCellInst_SboxInst_5_AND1_U1_n7,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND3_U1_n9, SubCellInst_SboxInst_5_AND3_U1_n8,
         SubCellInst_SboxInst_5_AND3_U1_n7,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND1_U1_n9, SubCellInst_SboxInst_6_AND1_U1_n8,
         SubCellInst_SboxInst_6_AND1_U1_n7,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND3_U1_n9, SubCellInst_SboxInst_6_AND3_U1_n8,
         SubCellInst_SboxInst_6_AND3_U1_n7,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND1_U1_n9, SubCellInst_SboxInst_7_AND1_U1_n8,
         SubCellInst_SboxInst_7_AND1_U1_n7,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND3_U1_n9, SubCellInst_SboxInst_7_AND3_U1_n8,
         SubCellInst_SboxInst_7_AND3_U1_n7,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND1_U1_n9, SubCellInst_SboxInst_8_AND1_U1_n8,
         SubCellInst_SboxInst_8_AND1_U1_n7,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND3_U1_n9, SubCellInst_SboxInst_8_AND3_U1_n8,
         SubCellInst_SboxInst_8_AND3_U1_n7,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND1_U1_n9, SubCellInst_SboxInst_9_AND1_U1_n8,
         SubCellInst_SboxInst_9_AND1_U1_n7,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND3_U1_n9, SubCellInst_SboxInst_9_AND3_U1_n8,
         SubCellInst_SboxInst_9_AND3_U1_n7,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND1_U1_n9,
         SubCellInst_SboxInst_10_AND1_U1_n8,
         SubCellInst_SboxInst_10_AND1_U1_n7,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND3_U1_n9,
         SubCellInst_SboxInst_10_AND3_U1_n8,
         SubCellInst_SboxInst_10_AND3_U1_n7,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND1_U1_n9,
         SubCellInst_SboxInst_11_AND1_U1_n8,
         SubCellInst_SboxInst_11_AND1_U1_n7,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND3_U1_n9,
         SubCellInst_SboxInst_11_AND3_U1_n8,
         SubCellInst_SboxInst_11_AND3_U1_n7,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND1_U1_n9,
         SubCellInst_SboxInst_12_AND1_U1_n8,
         SubCellInst_SboxInst_12_AND1_U1_n7,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND3_U1_n9,
         SubCellInst_SboxInst_12_AND3_U1_n8,
         SubCellInst_SboxInst_12_AND3_U1_n7,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND1_U1_n9,
         SubCellInst_SboxInst_13_AND1_U1_n8,
         SubCellInst_SboxInst_13_AND1_U1_n7,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND3_U1_n9,
         SubCellInst_SboxInst_13_AND3_U1_n8,
         SubCellInst_SboxInst_13_AND3_U1_n7,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND1_U1_n9,
         SubCellInst_SboxInst_14_AND1_U1_n8,
         SubCellInst_SboxInst_14_AND1_U1_n7,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND3_U1_n9,
         SubCellInst_SboxInst_14_AND3_U1_n8,
         SubCellInst_SboxInst_14_AND3_U1_n7,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND1_U1_n9,
         SubCellInst_SboxInst_15_AND1_U1_n8,
         SubCellInst_SboxInst_15_AND1_U1_n7,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND1_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND1_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND3_U1_n9,
         SubCellInst_SboxInst_15_AND3_U1_n8,
         SubCellInst_SboxInst_15_AND3_U1_n7,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND3_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND3_U1_z_1__1_,
         SubCellInst_SboxInst_0_AND2_U1_n9, SubCellInst_SboxInst_0_AND2_U1_n8,
         SubCellInst_SboxInst_0_AND2_U1_n7,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_0_AND4_U1_n9, SubCellInst_SboxInst_0_AND4_U1_n8,
         SubCellInst_SboxInst_0_AND4_U1_n7,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_0_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_0_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND2_U1_n9, SubCellInst_SboxInst_1_AND2_U1_n8,
         SubCellInst_SboxInst_1_AND2_U1_n7,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_1_AND4_U1_n9, SubCellInst_SboxInst_1_AND4_U1_n8,
         SubCellInst_SboxInst_1_AND4_U1_n7,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_1_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_1_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND2_U1_n9, SubCellInst_SboxInst_2_AND2_U1_n8,
         SubCellInst_SboxInst_2_AND2_U1_n7,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_2_AND4_U1_n9, SubCellInst_SboxInst_2_AND4_U1_n8,
         SubCellInst_SboxInst_2_AND4_U1_n7,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_2_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_2_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND2_U1_n9, SubCellInst_SboxInst_3_AND2_U1_n8,
         SubCellInst_SboxInst_3_AND2_U1_n7,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_3_AND4_U1_n9, SubCellInst_SboxInst_3_AND4_U1_n8,
         SubCellInst_SboxInst_3_AND4_U1_n7,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_3_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_3_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND2_U1_n9, SubCellInst_SboxInst_4_AND2_U1_n8,
         SubCellInst_SboxInst_4_AND2_U1_n7,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_4_AND4_U1_n9, SubCellInst_SboxInst_4_AND4_U1_n8,
         SubCellInst_SboxInst_4_AND4_U1_n7,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_4_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_4_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND2_U1_n9, SubCellInst_SboxInst_5_AND2_U1_n8,
         SubCellInst_SboxInst_5_AND2_U1_n7,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_5_AND4_U1_n9, SubCellInst_SboxInst_5_AND4_U1_n8,
         SubCellInst_SboxInst_5_AND4_U1_n7,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_5_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_5_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND2_U1_n9, SubCellInst_SboxInst_6_AND2_U1_n8,
         SubCellInst_SboxInst_6_AND2_U1_n7,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_6_AND4_U1_n9, SubCellInst_SboxInst_6_AND4_U1_n8,
         SubCellInst_SboxInst_6_AND4_U1_n7,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_6_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_6_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND2_U1_n9, SubCellInst_SboxInst_7_AND2_U1_n8,
         SubCellInst_SboxInst_7_AND2_U1_n7,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_7_AND4_U1_n9, SubCellInst_SboxInst_7_AND4_U1_n8,
         SubCellInst_SboxInst_7_AND4_U1_n7,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_7_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_7_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND2_U1_n9, SubCellInst_SboxInst_8_AND2_U1_n8,
         SubCellInst_SboxInst_8_AND2_U1_n7,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_8_AND4_U1_n9, SubCellInst_SboxInst_8_AND4_U1_n8,
         SubCellInst_SboxInst_8_AND4_U1_n7,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_8_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_8_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND2_U1_n9, SubCellInst_SboxInst_9_AND2_U1_n8,
         SubCellInst_SboxInst_9_AND2_U1_n7,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_9_AND4_U1_n9, SubCellInst_SboxInst_9_AND4_U1_n8,
         SubCellInst_SboxInst_9_AND4_U1_n7,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_9_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_9_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND2_U1_n9,
         SubCellInst_SboxInst_10_AND2_U1_n8,
         SubCellInst_SboxInst_10_AND2_U1_n7,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_10_AND4_U1_n9,
         SubCellInst_SboxInst_10_AND4_U1_n8,
         SubCellInst_SboxInst_10_AND4_U1_n7,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_10_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_10_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND2_U1_n9,
         SubCellInst_SboxInst_11_AND2_U1_n8,
         SubCellInst_SboxInst_11_AND2_U1_n7,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_11_AND4_U1_n9,
         SubCellInst_SboxInst_11_AND4_U1_n8,
         SubCellInst_SboxInst_11_AND4_U1_n7,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_11_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_11_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND2_U1_n9,
         SubCellInst_SboxInst_12_AND2_U1_n8,
         SubCellInst_SboxInst_12_AND2_U1_n7,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_12_AND4_U1_n9,
         SubCellInst_SboxInst_12_AND4_U1_n8,
         SubCellInst_SboxInst_12_AND4_U1_n7,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_12_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_12_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND2_U1_n9,
         SubCellInst_SboxInst_13_AND2_U1_n8,
         SubCellInst_SboxInst_13_AND2_U1_n7,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_13_AND4_U1_n9,
         SubCellInst_SboxInst_13_AND4_U1_n8,
         SubCellInst_SboxInst_13_AND4_U1_n7,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_13_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_13_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND2_U1_n9,
         SubCellInst_SboxInst_14_AND2_U1_n8,
         SubCellInst_SboxInst_14_AND2_U1_n7,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_14_AND4_U1_n9,
         SubCellInst_SboxInst_14_AND4_U1_n8,
         SubCellInst_SboxInst_14_AND4_U1_n7,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_14_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_14_AND4_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND2_U1_n9,
         SubCellInst_SboxInst_15_AND2_U1_n8,
         SubCellInst_SboxInst_15_AND2_U1_n7,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND2_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND2_U1_z_1__1_,
         SubCellInst_SboxInst_15_AND4_U1_n9,
         SubCellInst_SboxInst_15_AND4_U1_n8,
         SubCellInst_SboxInst_15_AND4_U1_n7,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_,
         SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_,
         SubCellInst_SboxInst_15_AND4_U1_z_0__0_,
         SubCellInst_SboxInst_15_AND4_U1_z_1__1_;
  wire   [63:0] TweakeyGeneration_StateRegInput;
  wire   [63:0] TweakeyGeneration_key_Feedback;
  wire   [4:1] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [5:4] FSM;
  wire   [63:0] StateRegInput;
  wire   [63:0] MCOutput;
  wire   [47:0] ShiftRowsOutput;
  wire   [63:32] AddRoundConstantOutput;
  wire   [63:60] SubCellOutput;
  wire   [1:0] SubCellInst_SboxInst_0_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_0_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND1_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND1_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND1_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND3_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND3_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND3_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_0_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_0_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_0_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_0_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_1_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_1_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_1_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_2_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_2_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_2_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_3_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_3_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_3_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_4_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_4_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_4_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_5_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_5_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_5_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_6_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_6_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_6_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_7_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_7_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_7_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_8_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_8_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_8_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_9_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_9_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_9_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_10_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_10_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_10_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_11_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_11_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_11_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_12_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_12_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_12_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_13_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_13_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_13_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_14_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_14_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_14_AND4_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND2_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND2_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND2_U1_mul;
  wire   [1:0] SubCellInst_SboxInst_15_AND4_U1_a_reg;
  wire   [1:0] SubCellInst_SboxInst_15_AND4_U1_mul_s1_out;
  wire   [1:0] SubCellInst_SboxInst_15_AND4_U1_mul;

  DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .D(FSMSelected[3]), .CK(
        clk_gated), .Q(FSMUpdate[4]), .QN(n16) );
  DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .D(FSMSelected[4]), .CK(
        clk_gated), .Q(FSM[4]), .QN(n14) );
  DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .D(FSMSelected[1]), .CK(
        clk_gated), .Q(FSM_1), .QN(n15) );
  DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .D(FSMSelected[0]), .CK(
        clk_gated), .Q(FSMUpdate[1]), .QN(n18) );
  DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .D(FSMSelected[5]), .CK(
        clk_gated), .Q(FSM[5]), .QN(n13) );
  DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .D(FSMSelected[2]), .CK(
        clk_gated), .Q(FSMUpdate[3]), .QN(n17) );
  INV_X1 U39 ( .A(rst), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n16), .A2(n17), .A3(FSM_1), .ZN(n36) );
  NOR2_X1 U41 ( .A1(n18), .A2(n36), .ZN(n31) );
  OAI21_X1 U42 ( .B1(n13), .B2(n31), .A(n14), .ZN(n32) );
  OAI211_X1 U43 ( .C1(n13), .C2(n14), .A(n30), .B(n32), .ZN(FSMSelected[0]) );
  NOR2_X1 U44 ( .A1(rst), .A2(n18), .ZN(FSMSelected[1]) );
  NOR2_X1 U45 ( .A1(rst), .A2(n16), .ZN(FSMSelected[4]) );
  NOR2_X1 U46 ( .A1(rst), .A2(n17), .ZN(FSMSelected[3]) );
  NOR2_X1 U47 ( .A1(FSMSelected[4]), .A2(FSMSelected[3]), .ZN(n35) );
  NAND2_X1 U48 ( .A1(n14), .A2(FSM[5]), .ZN(n33) );
  OAI21_X1 U49 ( .B1(n18), .B2(n33), .A(n30), .ZN(n34) );
  AOI21_X1 U50 ( .B1(n35), .B2(n34), .A(n15), .ZN(FSMSelected[2]) );
  NAND2_X1 U51 ( .A1(FSMSelected[1]), .A2(FSM[5]), .ZN(n37) );
  OAI22_X1 U52 ( .A1(rst), .A2(n14), .B1(n37), .B2(n36), .ZN(FSMSelected[5])
         );
  NAND4_X1 U53 ( .A1(n15), .A2(n16), .A3(n17), .A4(FSM[5]), .ZN(n38) );
  NOR3_X1 U54 ( .A1(n14), .A2(n18), .A3(n38), .ZN(done) );
  INV_X1 SubCellInst_SboxInst_0_U1_U1 ( .A(Ciphertext_s0[2]), .ZN(
        SubCellInst_SboxInst_0_n3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[2]), 
        .B(Ciphertext_s0[3]), .Z(SubCellInst_SboxInst_0_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[2]), 
        .B(Ciphertext_s1[3]), .Z(new_AGEMA_signal_1167) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[0]), 
        .B(Ciphertext_s0[2]), .Z(SubCellInst_SboxInst_0_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[0]), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1169) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_2_), .Z(SubCellInst_SboxInst_0_Q0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1169), .Z(new_AGEMA_signal_1453) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_XX_1_), .Z(SubCellInst_SboxInst_0_Q1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        new_AGEMA_signal_1167), .Z(new_AGEMA_signal_1454) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .ZN(SubCellInst_SboxInst_0_Q4) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1455) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_n3), .Z(
        SubCellInst_SboxInst_0_Q6) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1169), 
        .B(Ciphertext_s1[2]), .Z(new_AGEMA_signal_1456) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_Q1), .B(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_L1) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1454), 
        .B(new_AGEMA_signal_1456), .Z(new_AGEMA_signal_1550) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[1]), .B(
        SubCellInst_SboxInst_0_n3), .Z(SubCellInst_SboxInst_0_L2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[1]), .B(
        Ciphertext_s1[2]), .Z(new_AGEMA_signal_1457) );
  INV_X1 SubCellInst_SboxInst_1_U1_U1 ( .A(Ciphertext_s0[6]), .ZN(
        SubCellInst_SboxInst_1_n3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[6]), 
        .B(Ciphertext_s0[7]), .Z(SubCellInst_SboxInst_1_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[6]), 
        .B(Ciphertext_s1[7]), .Z(new_AGEMA_signal_1173) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[4]), 
        .B(Ciphertext_s0[6]), .Z(SubCellInst_SboxInst_1_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[4]), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1175) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_2_), .Z(SubCellInst_SboxInst_1_Q0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1175), .Z(new_AGEMA_signal_1459) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_XX_1_), .Z(SubCellInst_SboxInst_1_Q1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        new_AGEMA_signal_1173), .Z(new_AGEMA_signal_1460) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .ZN(SubCellInst_SboxInst_1_Q4) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1461) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_n3), .Z(
        SubCellInst_SboxInst_1_Q6) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1175), 
        .B(Ciphertext_s1[6]), .Z(new_AGEMA_signal_1462) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_Q1), .B(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_L1) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1460), 
        .B(new_AGEMA_signal_1462), .Z(new_AGEMA_signal_1553) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[5]), .B(
        SubCellInst_SboxInst_1_n3), .Z(SubCellInst_SboxInst_1_L2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[5]), .B(
        Ciphertext_s1[6]), .Z(new_AGEMA_signal_1463) );
  INV_X1 SubCellInst_SboxInst_2_U1_U1 ( .A(Ciphertext_s0[10]), .ZN(
        SubCellInst_SboxInst_2_n3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[10]), 
        .B(Ciphertext_s0[11]), .Z(SubCellInst_SboxInst_2_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[10]), 
        .B(Ciphertext_s1[11]), .Z(new_AGEMA_signal_1179) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[8]), 
        .B(Ciphertext_s0[10]), .Z(SubCellInst_SboxInst_2_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[8]), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1181) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_2_), .Z(SubCellInst_SboxInst_2_Q0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1181), .Z(new_AGEMA_signal_1465) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_XX_1_), .Z(SubCellInst_SboxInst_2_Q1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        new_AGEMA_signal_1179), .Z(new_AGEMA_signal_1466) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .ZN(SubCellInst_SboxInst_2_Q4) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1467) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_n3), .Z(
        SubCellInst_SboxInst_2_Q6) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1181), 
        .B(Ciphertext_s1[10]), .Z(new_AGEMA_signal_1468) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_Q1), .B(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_L1) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1466), 
        .B(new_AGEMA_signal_1468), .Z(new_AGEMA_signal_1556) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[9]), .B(
        SubCellInst_SboxInst_2_n3), .Z(SubCellInst_SboxInst_2_L2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[9]), .B(
        Ciphertext_s1[10]), .Z(new_AGEMA_signal_1469) );
  INV_X1 SubCellInst_SboxInst_3_U1_U1 ( .A(Ciphertext_s0[14]), .ZN(
        SubCellInst_SboxInst_3_n3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[14]), 
        .B(Ciphertext_s0[15]), .Z(SubCellInst_SboxInst_3_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[14]), 
        .B(Ciphertext_s1[15]), .Z(new_AGEMA_signal_1185) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[12]), 
        .B(Ciphertext_s0[14]), .Z(SubCellInst_SboxInst_3_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[12]), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1187) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_2_), .Z(SubCellInst_SboxInst_3_Q0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1187), .Z(new_AGEMA_signal_1471) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_XX_1_), .Z(SubCellInst_SboxInst_3_Q1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        new_AGEMA_signal_1185), .Z(new_AGEMA_signal_1472) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .ZN(SubCellInst_SboxInst_3_Q4) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1473) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_n3), .Z(
        SubCellInst_SboxInst_3_Q6) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1187), 
        .B(Ciphertext_s1[14]), .Z(new_AGEMA_signal_1474) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_Q1), .B(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_L1) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1472), 
        .B(new_AGEMA_signal_1474), .Z(new_AGEMA_signal_1559) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[13]), .B(
        SubCellInst_SboxInst_3_n3), .Z(SubCellInst_SboxInst_3_L2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[13]), .B(
        Ciphertext_s1[14]), .Z(new_AGEMA_signal_1475) );
  INV_X1 SubCellInst_SboxInst_4_U1_U1 ( .A(Ciphertext_s0[18]), .ZN(
        SubCellInst_SboxInst_4_n3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[18]), 
        .B(Ciphertext_s0[19]), .Z(SubCellInst_SboxInst_4_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[18]), 
        .B(Ciphertext_s1[19]), .Z(new_AGEMA_signal_1191) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[16]), 
        .B(Ciphertext_s0[18]), .Z(SubCellInst_SboxInst_4_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[16]), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1193) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_2_), .Z(SubCellInst_SboxInst_4_Q0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1193), .Z(new_AGEMA_signal_1477) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_XX_1_), .Z(SubCellInst_SboxInst_4_Q1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        new_AGEMA_signal_1191), .Z(new_AGEMA_signal_1478) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .ZN(SubCellInst_SboxInst_4_Q4) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1479) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_n3), .Z(
        SubCellInst_SboxInst_4_Q6) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1193), 
        .B(Ciphertext_s1[18]), .Z(new_AGEMA_signal_1480) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_Q1), .B(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_L1) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1478), 
        .B(new_AGEMA_signal_1480), .Z(new_AGEMA_signal_1562) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[17]), .B(
        SubCellInst_SboxInst_4_n3), .Z(SubCellInst_SboxInst_4_L2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[17]), .B(
        Ciphertext_s1[18]), .Z(new_AGEMA_signal_1481) );
  INV_X1 SubCellInst_SboxInst_5_U1_U1 ( .A(Ciphertext_s0[22]), .ZN(
        SubCellInst_SboxInst_5_n3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[22]), 
        .B(Ciphertext_s0[23]), .Z(SubCellInst_SboxInst_5_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[22]), 
        .B(Ciphertext_s1[23]), .Z(new_AGEMA_signal_1197) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[20]), 
        .B(Ciphertext_s0[22]), .Z(SubCellInst_SboxInst_5_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[20]), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1199) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_2_), .Z(SubCellInst_SboxInst_5_Q0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1199), .Z(new_AGEMA_signal_1483) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_XX_1_), .Z(SubCellInst_SboxInst_5_Q1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        new_AGEMA_signal_1197), .Z(new_AGEMA_signal_1484) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .ZN(SubCellInst_SboxInst_5_Q4) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1485) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_n3), .Z(
        SubCellInst_SboxInst_5_Q6) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1199), 
        .B(Ciphertext_s1[22]), .Z(new_AGEMA_signal_1486) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_Q1), .B(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_L1) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1484), 
        .B(new_AGEMA_signal_1486), .Z(new_AGEMA_signal_1565) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[21]), .B(
        SubCellInst_SboxInst_5_n3), .Z(SubCellInst_SboxInst_5_L2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[21]), .B(
        Ciphertext_s1[22]), .Z(new_AGEMA_signal_1487) );
  INV_X1 SubCellInst_SboxInst_6_U1_U1 ( .A(Ciphertext_s0[26]), .ZN(
        SubCellInst_SboxInst_6_n3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[26]), 
        .B(Ciphertext_s0[27]), .Z(SubCellInst_SboxInst_6_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[26]), 
        .B(Ciphertext_s1[27]), .Z(new_AGEMA_signal_1203) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[24]), 
        .B(Ciphertext_s0[26]), .Z(SubCellInst_SboxInst_6_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[24]), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1205) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_2_), .Z(SubCellInst_SboxInst_6_Q0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1205), .Z(new_AGEMA_signal_1489) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_XX_1_), .Z(SubCellInst_SboxInst_6_Q1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        new_AGEMA_signal_1203), .Z(new_AGEMA_signal_1490) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .ZN(SubCellInst_SboxInst_6_Q4) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1491) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_n3), .Z(
        SubCellInst_SboxInst_6_Q6) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1205), 
        .B(Ciphertext_s1[26]), .Z(new_AGEMA_signal_1492) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_Q1), .B(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_L1) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1490), 
        .B(new_AGEMA_signal_1492), .Z(new_AGEMA_signal_1568) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[25]), .B(
        SubCellInst_SboxInst_6_n3), .Z(SubCellInst_SboxInst_6_L2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[25]), .B(
        Ciphertext_s1[26]), .Z(new_AGEMA_signal_1493) );
  INV_X1 SubCellInst_SboxInst_7_U1_U1 ( .A(Ciphertext_s0[30]), .ZN(
        SubCellInst_SboxInst_7_n3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[30]), 
        .B(Ciphertext_s0[31]), .Z(SubCellInst_SboxInst_7_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[30]), 
        .B(Ciphertext_s1[31]), .Z(new_AGEMA_signal_1209) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[28]), 
        .B(Ciphertext_s0[30]), .Z(SubCellInst_SboxInst_7_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[28]), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1211) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_2_), .Z(SubCellInst_SboxInst_7_Q0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1211), .Z(new_AGEMA_signal_1495) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_XX_1_), .Z(SubCellInst_SboxInst_7_Q1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        new_AGEMA_signal_1209), .Z(new_AGEMA_signal_1496) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .ZN(SubCellInst_SboxInst_7_Q4) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1497) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_n3), .Z(
        SubCellInst_SboxInst_7_Q6) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1211), 
        .B(Ciphertext_s1[30]), .Z(new_AGEMA_signal_1498) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_Q1), .B(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_L1) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1496), 
        .B(new_AGEMA_signal_1498), .Z(new_AGEMA_signal_1571) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[29]), .B(
        SubCellInst_SboxInst_7_n3), .Z(SubCellInst_SboxInst_7_L2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[29]), .B(
        Ciphertext_s1[30]), .Z(new_AGEMA_signal_1499) );
  INV_X1 SubCellInst_SboxInst_8_U1_U1 ( .A(Ciphertext_s0[34]), .ZN(
        SubCellInst_SboxInst_8_n3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[34]), 
        .B(Ciphertext_s0[35]), .Z(SubCellInst_SboxInst_8_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[34]), 
        .B(Ciphertext_s1[35]), .Z(new_AGEMA_signal_1215) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[32]), 
        .B(Ciphertext_s0[34]), .Z(SubCellInst_SboxInst_8_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[32]), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1217) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_2_), .Z(SubCellInst_SboxInst_8_Q0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1217), .Z(new_AGEMA_signal_1501) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_XX_1_), .Z(SubCellInst_SboxInst_8_Q1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        new_AGEMA_signal_1215), .Z(new_AGEMA_signal_1502) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .ZN(SubCellInst_SboxInst_8_Q4) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1503) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_n3), .Z(
        SubCellInst_SboxInst_8_Q6) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1217), 
        .B(Ciphertext_s1[34]), .Z(new_AGEMA_signal_1504) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_Q1), .B(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_L1) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1502), 
        .B(new_AGEMA_signal_1504), .Z(new_AGEMA_signal_1574) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[33]), .B(
        SubCellInst_SboxInst_8_n3), .Z(SubCellInst_SboxInst_8_L2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[33]), .B(
        Ciphertext_s1[34]), .Z(new_AGEMA_signal_1505) );
  INV_X1 SubCellInst_SboxInst_9_U1_U1 ( .A(Ciphertext_s0[38]), .ZN(
        SubCellInst_SboxInst_9_n3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[38]), 
        .B(Ciphertext_s0[39]), .Z(SubCellInst_SboxInst_9_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[38]), 
        .B(Ciphertext_s1[39]), .Z(new_AGEMA_signal_1221) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[36]), 
        .B(Ciphertext_s0[38]), .Z(SubCellInst_SboxInst_9_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[36]), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1223) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_2_), .Z(SubCellInst_SboxInst_9_Q0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1223), .Z(new_AGEMA_signal_1507) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_XX_1_), .Z(SubCellInst_SboxInst_9_Q1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        new_AGEMA_signal_1221), .Z(new_AGEMA_signal_1508) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .ZN(SubCellInst_SboxInst_9_Q4) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1509) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_n3), .Z(
        SubCellInst_SboxInst_9_Q6) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1223), 
        .B(Ciphertext_s1[38]), .Z(new_AGEMA_signal_1510) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_Q1), .B(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_L1) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1508), 
        .B(new_AGEMA_signal_1510), .Z(new_AGEMA_signal_1577) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[37]), .B(
        SubCellInst_SboxInst_9_n3), .Z(SubCellInst_SboxInst_9_L2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[37]), .B(
        Ciphertext_s1[38]), .Z(new_AGEMA_signal_1511) );
  INV_X1 SubCellInst_SboxInst_10_U1_U1 ( .A(Ciphertext_s0[42]), .ZN(
        SubCellInst_SboxInst_10_n3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[42]), 
        .B(Ciphertext_s0[43]), .Z(SubCellInst_SboxInst_10_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[42]), 
        .B(Ciphertext_s1[43]), .Z(new_AGEMA_signal_1227) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[40]), 
        .B(Ciphertext_s0[42]), .Z(SubCellInst_SboxInst_10_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[40]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1229) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_2_), .Z(SubCellInst_SboxInst_10_Q0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1229), .Z(new_AGEMA_signal_1513) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_XX_1_), .Z(SubCellInst_SboxInst_10_Q1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(new_AGEMA_signal_1227), .Z(new_AGEMA_signal_1514) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .ZN(SubCellInst_SboxInst_10_Q4) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1515) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_n3), .Z(
        SubCellInst_SboxInst_10_Q6) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1229), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1516) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_Q1), .B(SubCellInst_SboxInst_10_Q6), .ZN(
        SubCellInst_SboxInst_10_L1) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1514), 
        .B(new_AGEMA_signal_1516), .Z(new_AGEMA_signal_1580) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[41]), 
        .B(SubCellInst_SboxInst_10_n3), .Z(SubCellInst_SboxInst_10_L2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[41]), 
        .B(Ciphertext_s1[42]), .Z(new_AGEMA_signal_1517) );
  INV_X1 SubCellInst_SboxInst_11_U1_U1 ( .A(Ciphertext_s0[46]), .ZN(
        SubCellInst_SboxInst_11_n3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[46]), 
        .B(Ciphertext_s0[47]), .Z(SubCellInst_SboxInst_11_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[46]), 
        .B(Ciphertext_s1[47]), .Z(new_AGEMA_signal_1233) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[44]), 
        .B(Ciphertext_s0[46]), .Z(SubCellInst_SboxInst_11_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[44]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1235) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_2_), .Z(SubCellInst_SboxInst_11_Q0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1235), .Z(new_AGEMA_signal_1519) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_XX_1_), .Z(SubCellInst_SboxInst_11_Q1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(new_AGEMA_signal_1233), .Z(new_AGEMA_signal_1520) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .ZN(SubCellInst_SboxInst_11_Q4) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1521) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_n3), .Z(
        SubCellInst_SboxInst_11_Q6) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1235), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1522) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_Q1), .B(SubCellInst_SboxInst_11_Q6), .ZN(
        SubCellInst_SboxInst_11_L1) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1520), 
        .B(new_AGEMA_signal_1522), .Z(new_AGEMA_signal_1583) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[45]), 
        .B(SubCellInst_SboxInst_11_n3), .Z(SubCellInst_SboxInst_11_L2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[45]), 
        .B(Ciphertext_s1[46]), .Z(new_AGEMA_signal_1523) );
  INV_X1 SubCellInst_SboxInst_12_U1_U1 ( .A(Ciphertext_s0[50]), .ZN(
        SubCellInst_SboxInst_12_n3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[50]), 
        .B(Ciphertext_s0[51]), .Z(SubCellInst_SboxInst_12_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[50]), 
        .B(Ciphertext_s1[51]), .Z(new_AGEMA_signal_1239) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[48]), 
        .B(Ciphertext_s0[50]), .Z(SubCellInst_SboxInst_12_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[48]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1241) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_2_), .Z(SubCellInst_SboxInst_12_Q0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1241), .Z(new_AGEMA_signal_1525) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_XX_1_), .Z(SubCellInst_SboxInst_12_Q1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(new_AGEMA_signal_1239), .Z(new_AGEMA_signal_1526) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .ZN(SubCellInst_SboxInst_12_Q4) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1527) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_n3), .Z(
        SubCellInst_SboxInst_12_Q6) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1241), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1528) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_Q1), .B(SubCellInst_SboxInst_12_Q6), .ZN(
        SubCellInst_SboxInst_12_L1) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1526), 
        .B(new_AGEMA_signal_1528), .Z(new_AGEMA_signal_1586) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[49]), 
        .B(SubCellInst_SboxInst_12_n3), .Z(SubCellInst_SboxInst_12_L2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[49]), 
        .B(Ciphertext_s1[50]), .Z(new_AGEMA_signal_1529) );
  INV_X1 SubCellInst_SboxInst_13_U1_U1 ( .A(Ciphertext_s0[54]), .ZN(
        SubCellInst_SboxInst_13_n3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[54]), 
        .B(Ciphertext_s0[55]), .Z(SubCellInst_SboxInst_13_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[54]), 
        .B(Ciphertext_s1[55]), .Z(new_AGEMA_signal_1245) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[52]), 
        .B(Ciphertext_s0[54]), .Z(SubCellInst_SboxInst_13_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[52]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1247) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_2_), .Z(SubCellInst_SboxInst_13_Q0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1247), .Z(new_AGEMA_signal_1531) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_XX_1_), .Z(SubCellInst_SboxInst_13_Q1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(new_AGEMA_signal_1245), .Z(new_AGEMA_signal_1532) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .ZN(SubCellInst_SboxInst_13_Q4) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1533) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_n3), .Z(
        SubCellInst_SboxInst_13_Q6) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1247), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1534) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_Q1), .B(SubCellInst_SboxInst_13_Q6), .ZN(
        SubCellInst_SboxInst_13_L1) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1532), 
        .B(new_AGEMA_signal_1534), .Z(new_AGEMA_signal_1589) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[53]), 
        .B(SubCellInst_SboxInst_13_n3), .Z(SubCellInst_SboxInst_13_L2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[53]), 
        .B(Ciphertext_s1[54]), .Z(new_AGEMA_signal_1535) );
  INV_X1 SubCellInst_SboxInst_14_U1_U1 ( .A(Ciphertext_s0[58]), .ZN(
        SubCellInst_SboxInst_14_n3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[58]), 
        .B(Ciphertext_s0[59]), .Z(SubCellInst_SboxInst_14_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[58]), 
        .B(Ciphertext_s1[59]), .Z(new_AGEMA_signal_1251) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[56]), 
        .B(Ciphertext_s0[58]), .Z(SubCellInst_SboxInst_14_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[56]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1253) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_2_), .Z(SubCellInst_SboxInst_14_Q0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1253), .Z(new_AGEMA_signal_1537) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_XX_1_), .Z(SubCellInst_SboxInst_14_Q1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(new_AGEMA_signal_1251), .Z(new_AGEMA_signal_1538) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .ZN(SubCellInst_SboxInst_14_Q4) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1539) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_n3), .Z(
        SubCellInst_SboxInst_14_Q6) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1253), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1540) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_Q1), .B(SubCellInst_SboxInst_14_Q6), .ZN(
        SubCellInst_SboxInst_14_L1) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1538), 
        .B(new_AGEMA_signal_1540), .Z(new_AGEMA_signal_1592) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[57]), 
        .B(SubCellInst_SboxInst_14_n3), .Z(SubCellInst_SboxInst_14_L2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[57]), 
        .B(Ciphertext_s1[58]), .Z(new_AGEMA_signal_1541) );
  INV_X1 SubCellInst_SboxInst_15_U1_U1 ( .A(Ciphertext_s0[62]), .ZN(
        SubCellInst_SboxInst_15_n3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_0_U1 ( .A(Ciphertext_s0[62]), 
        .B(Ciphertext_s0[63]), .Z(SubCellInst_SboxInst_15_XX_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i1_U1_Ins_1_U1 ( .A(Ciphertext_s1[62]), 
        .B(Ciphertext_s1[63]), .Z(new_AGEMA_signal_1257) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_0_U1 ( .A(Ciphertext_s0[60]), 
        .B(Ciphertext_s0[62]), .Z(SubCellInst_SboxInst_15_XX_2_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_i2_U1_Ins_1_U1 ( .A(Ciphertext_s1[60]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1259) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_2_), .Z(SubCellInst_SboxInst_15_Q0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR0_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1259), .Z(new_AGEMA_signal_1543) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_XX_1_), .Z(SubCellInst_SboxInst_15_Q1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR1_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(new_AGEMA_signal_1257), .Z(new_AGEMA_signal_1544) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .ZN(SubCellInst_SboxInst_15_Q4) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR3_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1545) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_n3), .Z(
        SubCellInst_SboxInst_15_Q6) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1259), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1546) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_Q1), .B(SubCellInst_SboxInst_15_Q6), .ZN(
        SubCellInst_SboxInst_15_L1) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1544), 
        .B(new_AGEMA_signal_1546), .Z(new_AGEMA_signal_1595) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_0_U1 ( .A(Ciphertext_s0[61]), 
        .B(SubCellInst_SboxInst_15_n3), .Z(SubCellInst_SboxInst_15_L2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR8_U1_Ins_1_U1 ( .A(Ciphertext_s1[61]), 
        .B(Ciphertext_s1[62]), .Z(new_AGEMA_signal_1547) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[0]), .B(Key_s0[0]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[0]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_0_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1260), .B(Key_s1[0]), .S(rst), .Z(
        new_AGEMA_signal_1262) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[1]), .B(Key_s0[1]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[1]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1263), .B(Key_s1[1]), .S(rst), .Z(
        new_AGEMA_signal_1265) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[2]), .B(Key_s0[2]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[2]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_2_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1266), .B(Key_s1[2]), .S(rst), .Z(
        new_AGEMA_signal_1268) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[3]), .B(Key_s0[3]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[3]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_3_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1269), .B(Key_s1[3]), .S(rst), .Z(
        new_AGEMA_signal_1271) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[4]), .B(Key_s0[4]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[4]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_4_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1272), .B(Key_s1[4]), .S(rst), .Z(
        new_AGEMA_signal_1274) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[5]), .B(Key_s0[5]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[5]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_5_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1275), .B(Key_s1[5]), .S(rst), .Z(
        new_AGEMA_signal_1277) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[6]), .B(Key_s0[6]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[6]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_6_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1278), .B(Key_s1[6]), .S(rst), .Z(
        new_AGEMA_signal_1280) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[7]), .B(Key_s0[7]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[7]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_7_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1281), .B(Key_s1[7]), .S(rst), .Z(
        new_AGEMA_signal_1283) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[8]), .B(Key_s0[8]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[8]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_8_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1284), .B(Key_s1[8]), .S(rst), .Z(
        new_AGEMA_signal_1286) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[9]), .B(Key_s0[9]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[9]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_9_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1287), .B(Key_s1[9]), .S(rst), .Z(
        new_AGEMA_signal_1289) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[10]), .B(Key_s0[10]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[10]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_10_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1290), .B(Key_s1[10]), .S(rst), .Z(
        new_AGEMA_signal_1292) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[11]), .B(Key_s0[11]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[11]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_11_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1293), .B(Key_s1[11]), .S(rst), .Z(
        new_AGEMA_signal_1295) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[12]), .B(Key_s0[12]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[12]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_12_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1296), .B(Key_s1[12]), .S(rst), .Z(
        new_AGEMA_signal_1298) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[13]), .B(Key_s0[13]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[13]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_13_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1299), .B(Key_s1[13]), .S(rst), .Z(
        new_AGEMA_signal_1301) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[14]), .B(Key_s0[14]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[14]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_14_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1302), .B(Key_s1[14]), .S(rst), .Z(
        new_AGEMA_signal_1304) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[15]), .B(Key_s0[15]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[15]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_15_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1305), .B(Key_s1[15]), .S(rst), .Z(
        new_AGEMA_signal_1307) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[16]), .B(Key_s0[16]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[16]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_16_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1308), .B(Key_s1[16]), .S(rst), .Z(
        new_AGEMA_signal_1310) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[17]), .B(Key_s0[17]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[17]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_17_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1311), .B(Key_s1[17]), .S(rst), .Z(
        new_AGEMA_signal_1313) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[18]), .B(Key_s0[18]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[18]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_18_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1314), .B(Key_s1[18]), .S(rst), .Z(
        new_AGEMA_signal_1316) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[19]), .B(Key_s0[19]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[19]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_19_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1317), .B(Key_s1[19]), .S(rst), .Z(
        new_AGEMA_signal_1319) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[20]), .B(Key_s0[20]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[20]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_20_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1320), .B(Key_s1[20]), .S(rst), .Z(
        new_AGEMA_signal_1322) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[21]), .B(Key_s0[21]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[21]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_21_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1323), .B(Key_s1[21]), .S(rst), .Z(
        new_AGEMA_signal_1325) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[22]), .B(Key_s0[22]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[22]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_22_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1326), .B(Key_s1[22]), .S(rst), .Z(
        new_AGEMA_signal_1328) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[23]), .B(Key_s0[23]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[23]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_23_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1329), .B(Key_s1[23]), .S(rst), .Z(
        new_AGEMA_signal_1331) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[24]), .B(Key_s0[24]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[24]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_24_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1332), .B(Key_s1[24]), .S(rst), .Z(
        new_AGEMA_signal_1334) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[25]), .B(Key_s0[25]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[25]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_25_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1335), .B(Key_s1[25]), .S(rst), .Z(
        new_AGEMA_signal_1337) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[26]), .B(Key_s0[26]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[26]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_26_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1338), .B(Key_s1[26]), .S(rst), .Z(
        new_AGEMA_signal_1340) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[27]), .B(Key_s0[27]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[27]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_27_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1341), .B(Key_s1[27]), .S(rst), .Z(
        new_AGEMA_signal_1343) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[28]), .B(Key_s0[28]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[28]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_28_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1344), .B(Key_s1[28]), .S(rst), .Z(
        new_AGEMA_signal_1346) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[29]), .B(Key_s0[29]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[29]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_29_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1347), .B(Key_s1[29]), .S(rst), .Z(
        new_AGEMA_signal_1349) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[30]), .B(Key_s0[30]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[30]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_30_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1350), .B(Key_s1[30]), .S(rst), .Z(
        new_AGEMA_signal_1352) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[31]), .B(Key_s0[31]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[31]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_31_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1353), .B(Key_s1[31]), .S(rst), .Z(
        new_AGEMA_signal_1355) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[32]), .B(Key_s0[32]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[32]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_32_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1356), .B(Key_s1[32]), .S(rst), .Z(
        new_AGEMA_signal_1358) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[33]), .B(Key_s0[33]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[33]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_33_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1359), .B(Key_s1[33]), .S(rst), .Z(
        new_AGEMA_signal_1361) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[34]), .B(Key_s0[34]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[34]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_34_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1362), .B(Key_s1[34]), .S(rst), .Z(
        new_AGEMA_signal_1364) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[35]), .B(Key_s0[35]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[35]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_35_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1365), .B(Key_s1[35]), .S(rst), .Z(
        new_AGEMA_signal_1367) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[36]), .B(Key_s0[36]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[36]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_36_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1368), .B(Key_s1[36]), .S(rst), .Z(
        new_AGEMA_signal_1370) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[37]), .B(Key_s0[37]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[37]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_37_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1371), .B(Key_s1[37]), .S(rst), .Z(
        new_AGEMA_signal_1373) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[38]), .B(Key_s0[38]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[38]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_38_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1374), .B(Key_s1[38]), .S(rst), .Z(
        new_AGEMA_signal_1376) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[39]), .B(Key_s0[39]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[39]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_39_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1377), .B(Key_s1[39]), .S(rst), .Z(
        new_AGEMA_signal_1379) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[40]), .B(Key_s0[40]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[40]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_40_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1380), .B(Key_s1[40]), .S(rst), .Z(
        new_AGEMA_signal_1382) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[41]), .B(Key_s0[41]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[41]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_41_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1383), .B(Key_s1[41]), .S(rst), .Z(
        new_AGEMA_signal_1385) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[42]), .B(Key_s0[42]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[42]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_42_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1386), .B(Key_s1[42]), .S(rst), .Z(
        new_AGEMA_signal_1388) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[43]), .B(Key_s0[43]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[43]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_43_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1389), .B(Key_s1[43]), .S(rst), .Z(
        new_AGEMA_signal_1391) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[44]), .B(Key_s0[44]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[44]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_44_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1392), .B(Key_s1[44]), .S(rst), .Z(
        new_AGEMA_signal_1394) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[45]), .B(Key_s0[45]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[45]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_45_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1395), .B(Key_s1[45]), .S(rst), .Z(
        new_AGEMA_signal_1397) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[46]), .B(Key_s0[46]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[46]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_46_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1398), .B(Key_s1[46]), .S(rst), .Z(
        new_AGEMA_signal_1400) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[47]), .B(Key_s0[47]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[47]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_47_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1401), .B(Key_s1[47]), .S(rst), .Z(
        new_AGEMA_signal_1403) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[48]), .B(Key_s0[48]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[48]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_48_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1404), .B(Key_s1[48]), .S(rst), .Z(
        new_AGEMA_signal_1406) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[49]), .B(Key_s0[49]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[49]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_49_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1407), .B(Key_s1[49]), .S(rst), .Z(
        new_AGEMA_signal_1409) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[50]), .B(Key_s0[50]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[50]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_50_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1410), .B(Key_s1[50]), .S(rst), .Z(
        new_AGEMA_signal_1412) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[51]), .B(Key_s0[51]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[51]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_51_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1413), .B(Key_s1[51]), .S(rst), .Z(
        new_AGEMA_signal_1415) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[52]), .B(Key_s0[52]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[52]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_52_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1416), .B(Key_s1[52]), .S(rst), .Z(
        new_AGEMA_signal_1418) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[53]), .B(Key_s0[53]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[53]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_53_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1419), .B(Key_s1[53]), .S(rst), .Z(
        new_AGEMA_signal_1421) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[54]), .B(Key_s0[54]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[54]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_54_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1422), .B(Key_s1[54]), .S(rst), .Z(
        new_AGEMA_signal_1424) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[55]), .B(Key_s0[55]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[55]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_55_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1425), .B(Key_s1[55]), .S(rst), .Z(
        new_AGEMA_signal_1427) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[56]), .B(Key_s0[56]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[56]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_56_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1428), .B(Key_s1[56]), .S(rst), .Z(
        new_AGEMA_signal_1430) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[57]), .B(Key_s0[57]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[57]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_57_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1431), .B(Key_s1[57]), .S(rst), .Z(
        new_AGEMA_signal_1433) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[58]), .B(Key_s0[58]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[58]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_58_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1434), .B(Key_s1[58]), .S(rst), .Z(
        new_AGEMA_signal_1436) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[59]), .B(Key_s0[59]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[59]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_59_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1437), .B(Key_s1[59]), .S(rst), .Z(
        new_AGEMA_signal_1439) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[60]), .B(Key_s0[60]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[60]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_60_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1440), .B(Key_s1[60]), .S(rst), .Z(
        new_AGEMA_signal_1442) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[61]), .B(Key_s0[61]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[61]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_61_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1443), .B(Key_s1[61]), .S(rst), .Z(
        new_AGEMA_signal_1445) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[62]), .B(Key_s0[62]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[62]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_62_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1446), .B(Key_s1[62]), .S(rst), .Z(
        new_AGEMA_signal_1448) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_0_U1 ( .A(
        TweakeyGeneration_key_Feedback[63]), .B(Key_s0[63]), .S(rst), .Z(
        TweakeyGeneration_StateRegInput[63]) );
  MUX2_X1 TweakeyGeneration_KEYMUX_MUXInst_63_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1449), .B(Key_s1[63]), .S(rst), .Z(
        new_AGEMA_signal_1451) );
  NOR2_X1 ClockGatingInst_U9 ( .A1(rst), .A2(ClockGatingInst_n9), .ZN(
        ClockGatingInst_n4) );
  NOR2_X1 ClockGatingInst_U8 ( .A1(rst), .A2(ClockGatingInst_n8), .ZN(
        ClockGatingInst_n3) );
  NOR2_X1 ClockGatingInst_U7 ( .A1(rst), .A2(ClockGatingInst_n7), .ZN(
        ClockGatingInst_n2) );
  NOR2_X1 ClockGatingInst_U6 ( .A1(rst), .A2(ClockGatingInst_n6), .ZN(
        ClockGatingInst_n1) );
  NAND2_X1 ClockGatingInst_U5 ( .A1(ClockGatingInst_n10), .A2(
        ClockGatingInst_n11), .ZN(ClockGatingInst_N7) );
  AND2_X1 ClockGatingInst_U4 ( .A1(ClockGatingInst_LatchedEnable), .A2(clk), 
        .ZN(clk_gated) );
  INV_X1 ClockGatingInst_U3 ( .A(rst), .ZN(ClockGatingInst_n11) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_2_ ( .D(ClockGatingInst_n1), .CK(
        clk), .Q(), .QN(ClockGatingInst_n7) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_3_ ( .D(ClockGatingInst_n2), .CK(
        clk), .Q(), .QN(ClockGatingInst_n8) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_4_ ( .D(ClockGatingInst_n3), .CK(
        clk), .Q(), .QN(ClockGatingInst_n9) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_5_ ( .D(ClockGatingInst_n4), .CK(
        clk), .Q(ClockGatingInst_ShiftRegister_5_), .QN(ClockGatingInst_n10)
         );
  DLL_X1 ClockGatingInst_LatchedEnable_reg ( .D(ClockGatingInst_N7), .GN(clk), 
        .Q(ClockGatingInst_LatchedEnable) );
  DLL_X1 ClockGatingInst_Synch_reg ( .D(ClockGatingInst_ShiftRegister_5_), 
        .GN(clk), .Q(Synch) );
  DFF_X1 ClockGatingInst_ShiftRegister_reg_1_ ( .D(ClockGatingInst_N7), .CK(
        clk), .Q(), .QN(ClockGatingInst_n6) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_0_U1 ( .A(MCOutput[2]), .B(
        Plaintext_s0[2]), .S(rst), .Z(StateRegInput[2]) );
  MUX2_X1 PlaintextMUX_MUXInst_2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1915), .B(
        Plaintext_s1[2]), .S(rst), .Z(new_AGEMA_signal_1922) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_0_U1 ( .A(MCOutput[3]), .B(
        Plaintext_s0[3]), .S(rst), .Z(StateRegInput[3]) );
  MUX2_X1 PlaintextMUX_MUXInst_3_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1975), .B(
        Plaintext_s1[3]), .S(rst), .Z(new_AGEMA_signal_1982) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_0_U1 ( .A(MCOutput[6]), .B(
        Plaintext_s0[6]), .S(rst), .Z(StateRegInput[6]) );
  MUX2_X1 PlaintextMUX_MUXInst_6_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1917), .B(
        Plaintext_s1[6]), .S(rst), .Z(new_AGEMA_signal_1924) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_0_U1 ( .A(MCOutput[7]), .B(
        Plaintext_s0[7]), .S(rst), .Z(StateRegInput[7]) );
  MUX2_X1 PlaintextMUX_MUXInst_7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1977), .B(
        Plaintext_s1[7]), .S(rst), .Z(new_AGEMA_signal_1984) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_0_U1 ( .A(MCOutput[10]), .B(
        Plaintext_s0[10]), .S(rst), .Z(StateRegInput[10]) );
  MUX2_X1 PlaintextMUX_MUXInst_10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1919), .B(
        Plaintext_s1[10]), .S(rst), .Z(new_AGEMA_signal_1926) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_0_U1 ( .A(MCOutput[11]), .B(
        Plaintext_s0[11]), .S(rst), .Z(StateRegInput[11]) );
  MUX2_X1 PlaintextMUX_MUXInst_11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1979), .B(
        Plaintext_s1[11]), .S(rst), .Z(new_AGEMA_signal_1986) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_0_U1 ( .A(MCOutput[14]), .B(
        Plaintext_s0[14]), .S(rst), .Z(StateRegInput[14]) );
  MUX2_X1 PlaintextMUX_MUXInst_14_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2033), .B(
        Plaintext_s1[14]), .S(rst), .Z(new_AGEMA_signal_2042) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_0_U1 ( .A(MCOutput[15]), .B(
        Plaintext_s0[15]), .S(rst), .Z(StateRegInput[15]) );
  MUX2_X1 PlaintextMUX_MUXInst_15_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2077), .B(
        Plaintext_s1[15]), .S(rst), .Z(new_AGEMA_signal_2085) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_0_U1 ( .A(MCOutput[18]), .B(
        Plaintext_s0[18]), .S(rst), .Z(StateRegInput[18]) );
  MUX2_X1 PlaintextMUX_MUXInst_18_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1909), .B(
        Plaintext_s1[18]), .S(rst), .Z(new_AGEMA_signal_1928) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_0_U1 ( .A(MCOutput[19]), .B(
        Plaintext_s0[19]), .S(rst), .Z(StateRegInput[19]) );
  MUX2_X1 PlaintextMUX_MUXInst_19_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1968), .B(
        Plaintext_s1[19]), .S(rst), .Z(new_AGEMA_signal_1988) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_0_U1 ( .A(MCOutput[22]), .B(
        Plaintext_s0[22]), .S(rst), .Z(StateRegInput[22]) );
  MUX2_X1 PlaintextMUX_MUXInst_22_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1911), .B(
        Plaintext_s1[22]), .S(rst), .Z(new_AGEMA_signal_1930) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_0_U1 ( .A(MCOutput[23]), .B(
        Plaintext_s0[23]), .S(rst), .Z(StateRegInput[23]) );
  MUX2_X1 PlaintextMUX_MUXInst_23_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1970), .B(
        Plaintext_s1[23]), .S(rst), .Z(new_AGEMA_signal_1990) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_0_U1 ( .A(MCOutput[26]), .B(
        Plaintext_s0[26]), .S(rst), .Z(StateRegInput[26]) );
  MUX2_X1 PlaintextMUX_MUXInst_26_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2023), .B(
        Plaintext_s1[26]), .S(rst), .Z(new_AGEMA_signal_2048) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_0_U1 ( .A(MCOutput[27]), .B(
        Plaintext_s0[27]), .S(rst), .Z(StateRegInput[27]) );
  MUX2_X1 PlaintextMUX_MUXInst_27_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2071), .B(
        Plaintext_s1[27]), .S(rst), .Z(new_AGEMA_signal_2091) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_0_U1 ( .A(MCOutput[30]), .B(
        Plaintext_s0[30]), .S(rst), .Z(StateRegInput[30]) );
  MUX2_X1 PlaintextMUX_MUXInst_30_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1913), .B(
        Plaintext_s1[30]), .S(rst), .Z(new_AGEMA_signal_1932) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_0_U1 ( .A(MCOutput[31]), .B(
        Plaintext_s0[31]), .S(rst), .Z(StateRegInput[31]) );
  MUX2_X1 PlaintextMUX_MUXInst_31_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1973), .B(
        Plaintext_s1[31]), .S(rst), .Z(new_AGEMA_signal_1992) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_0_U1 ( .A(MCOutput[34]), .B(
        Plaintext_s0[34]), .S(rst), .Z(StateRegInput[34]) );
  MUX2_X1 PlaintextMUX_MUXInst_34_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1810), .B(
        Plaintext_s1[34]), .S(rst), .Z(new_AGEMA_signal_1821) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_0_U1 ( .A(MCOutput[35]), .B(
        Plaintext_s0[35]), .S(rst), .Z(StateRegInput[35]) );
  MUX2_X1 PlaintextMUX_MUXInst_35_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1854), .B(
        Plaintext_s1[35]), .S(rst), .Z(new_AGEMA_signal_1874) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_0_U1 ( .A(MCOutput[38]), .B(
        Plaintext_s0[38]), .S(rst), .Z(StateRegInput[38]) );
  MUX2_X1 PlaintextMUX_MUXInst_38_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1812), .B(
        Plaintext_s1[38]), .S(rst), .Z(new_AGEMA_signal_1823) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_0_U1 ( .A(MCOutput[39]), .B(
        Plaintext_s0[39]), .S(rst), .Z(StateRegInput[39]) );
  MUX2_X1 PlaintextMUX_MUXInst_39_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1856), .B(
        Plaintext_s1[39]), .S(rst), .Z(new_AGEMA_signal_1876) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_0_U1 ( .A(MCOutput[42]), .B(
        Plaintext_s0[42]), .S(rst), .Z(StateRegInput[42]) );
  MUX2_X1 PlaintextMUX_MUXInst_42_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1814), .B(
        Plaintext_s1[42]), .S(rst), .Z(new_AGEMA_signal_1825) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_0_U1 ( .A(MCOutput[43]), .B(
        Plaintext_s0[43]), .S(rst), .Z(StateRegInput[43]) );
  MUX2_X1 PlaintextMUX_MUXInst_43_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1858), .B(
        Plaintext_s1[43]), .S(rst), .Z(new_AGEMA_signal_1878) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_0_U1 ( .A(MCOutput[46]), .B(
        Plaintext_s0[46]), .S(rst), .Z(StateRegInput[46]) );
  MUX2_X1 PlaintextMUX_MUXInst_46_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1898), .B(
        Plaintext_s1[46]), .S(rst), .Z(new_AGEMA_signal_1940) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_0_U1 ( .A(MCOutput[47]), .B(
        Plaintext_s0[47]), .S(rst), .Z(StateRegInput[47]) );
  MUX2_X1 PlaintextMUX_MUXInst_47_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1958), .B(
        Plaintext_s1[47]), .S(rst), .Z(new_AGEMA_signal_2000) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_0_U1 ( .A(MCOutput[50]), .B(
        Plaintext_s0[50]), .S(rst), .Z(StateRegInput[50]) );
  MUX2_X1 PlaintextMUX_MUXInst_50_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1901), .B(
        Plaintext_s1[50]), .S(rst), .Z(new_AGEMA_signal_1942) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_0_U1 ( .A(MCOutput[51]), .B(
        Plaintext_s0[51]), .S(rst), .Z(StateRegInput[51]) );
  MUX2_X1 PlaintextMUX_MUXInst_51_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1960), .B(
        Plaintext_s1[51]), .S(rst), .Z(new_AGEMA_signal_2002) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_0_U1 ( .A(MCOutput[54]), .B(
        Plaintext_s0[54]), .S(rst), .Z(StateRegInput[54]) );
  MUX2_X1 PlaintextMUX_MUXInst_54_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1903), .B(
        Plaintext_s1[54]), .S(rst), .Z(new_AGEMA_signal_1944) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_0_U1 ( .A(MCOutput[55]), .B(
        Plaintext_s0[55]), .S(rst), .Z(StateRegInput[55]) );
  MUX2_X1 PlaintextMUX_MUXInst_55_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1963), .B(
        Plaintext_s1[55]), .S(rst), .Z(new_AGEMA_signal_2004) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_0_U1 ( .A(MCOutput[58]), .B(
        Plaintext_s0[58]), .S(rst), .Z(StateRegInput[58]) );
  MUX2_X1 PlaintextMUX_MUXInst_58_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1906), .B(
        Plaintext_s1[58]), .S(rst), .Z(new_AGEMA_signal_1946) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_0_U1 ( .A(MCOutput[59]), .B(
        Plaintext_s0[59]), .S(rst), .Z(StateRegInput[59]) );
  MUX2_X1 PlaintextMUX_MUXInst_59_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1965), .B(
        Plaintext_s1[59]), .S(rst), .Z(new_AGEMA_signal_2006) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_0_U1 ( .A(MCOutput[62]), .B(
        Plaintext_s0[62]), .S(rst), .Z(StateRegInput[62]) );
  MUX2_X1 PlaintextMUX_MUXInst_62_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2017), .B(
        Plaintext_s1[62]), .S(rst), .Z(new_AGEMA_signal_2060) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_0_U1 ( .A(MCOutput[63]), .B(
        Plaintext_s0[63]), .S(rst), .Z(StateRegInput[63]) );
  MUX2_X1 PlaintextMUX_MUXInst_63_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2067), .B(
        Plaintext_s1[63]), .S(rst), .Z(new_AGEMA_signal_2103) );
  INV_X1 SubCellInst_SboxInst_0_U3_U1 ( .A(SubCellInst_SboxInst_0_YY_1_), .ZN(
        ShiftRowsOutput[7]) );
  INV_X1 SubCellInst_SboxInst_0_U2_U1 ( .A(SubCellInst_SboxInst_0_YY_0_), .ZN(
        ShiftRowsOutput[6]) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U14 ( .A(Fresh[0]), .B(
        SubCellInst_SboxInst_0_Q1), .Z(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U13 ( .A(Fresh[0]), .B(
        new_AGEMA_signal_1454), .Z(SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U10 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND1_U1_U8 ( .A(Fresh[0]), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U7 ( .A1(new_AGEMA_signal_1454), .A2(
        Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q1), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n8), .B(
        SubCellInst_SboxInst_0_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1548) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_n7), .B(
        SubCellInst_SboxInst_0_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T0) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_Q0), .B(SubCellInst_SboxInst_0_T0), .Z(
        SubCellInst_SboxInst_0_Q2) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1453), 
        .B(new_AGEMA_signal_1548), .Z(new_AGEMA_signal_1596) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U14 ( .A(Fresh[1]), .B(
        SubCellInst_SboxInst_0_Q4), .Z(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U13 ( .A(Fresh[1]), .B(
        new_AGEMA_signal_1455), .Z(SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U10 ( .A1(Ciphertext_s1[2]), .A2(
        SubCellInst_SboxInst_0_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_0_n3), 
        .A2(SubCellInst_SboxInst_0_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND3_U1_U8 ( .A(Fresh[1]), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U7 ( .A1(new_AGEMA_signal_1455), .A2(
        Ciphertext_s1[2]), .ZN(SubCellInst_SboxInst_0_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q4), 
        .A2(SubCellInst_SboxInst_0_n3), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n8), .B(
        SubCellInst_SboxInst_0_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1549) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_n7), .B(
        SubCellInst_SboxInst_0_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T2) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[2]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L1), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_Q7) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1550), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1597) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_2_), .B(SubCellInst_SboxInst_0_T0), .Z(
        SubCellInst_SboxInst_0_L3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1169), 
        .B(new_AGEMA_signal_1548), .Z(new_AGEMA_signal_1598) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L3), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1598), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1724) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_XX_1_), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1167), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1660) );
  INV_X1 SubCellInst_SboxInst_1_U3_U1 ( .A(SubCellInst_SboxInst_1_YY_1_), .ZN(
        ShiftRowsOutput[11]) );
  INV_X1 SubCellInst_SboxInst_1_U2_U1 ( .A(SubCellInst_SboxInst_1_YY_0_), .ZN(
        ShiftRowsOutput[10]) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U14 ( .A(Fresh[2]), .B(
        SubCellInst_SboxInst_1_Q1), .Z(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U13 ( .A(Fresh[2]), .B(
        new_AGEMA_signal_1460), .Z(SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U10 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND1_U1_U8 ( .A(Fresh[2]), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U7 ( .A1(new_AGEMA_signal_1460), .A2(
        Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q1), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n8), .B(
        SubCellInst_SboxInst_1_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1551) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_n7), .B(
        SubCellInst_SboxInst_1_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T0) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_Q0), .B(SubCellInst_SboxInst_1_T0), .Z(
        SubCellInst_SboxInst_1_Q2) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1459), 
        .B(new_AGEMA_signal_1551), .Z(new_AGEMA_signal_1600) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U14 ( .A(Fresh[3]), .B(
        SubCellInst_SboxInst_1_Q4), .Z(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U13 ( .A(Fresh[3]), .B(
        new_AGEMA_signal_1461), .Z(SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U10 ( .A1(Ciphertext_s1[6]), .A2(
        SubCellInst_SboxInst_1_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_1_n3), 
        .A2(SubCellInst_SboxInst_1_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND3_U1_U8 ( .A(Fresh[3]), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U7 ( .A1(new_AGEMA_signal_1461), .A2(
        Ciphertext_s1[6]), .ZN(SubCellInst_SboxInst_1_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q4), 
        .A2(SubCellInst_SboxInst_1_n3), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n8), .B(
        SubCellInst_SboxInst_1_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1552) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_n7), .B(
        SubCellInst_SboxInst_1_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T2) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[6]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L1), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_Q7) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1553), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1601) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_2_), .B(SubCellInst_SboxInst_1_T0), .Z(
        SubCellInst_SboxInst_1_L3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1175), 
        .B(new_AGEMA_signal_1551), .Z(new_AGEMA_signal_1602) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L3), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1602), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1726) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_XX_1_), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1173), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1664) );
  INV_X1 SubCellInst_SboxInst_2_U3_U1 ( .A(SubCellInst_SboxInst_2_YY_1_), .ZN(
        ShiftRowsOutput[15]) );
  INV_X1 SubCellInst_SboxInst_2_U2_U1 ( .A(SubCellInst_SboxInst_2_YY_0_), .ZN(
        ShiftRowsOutput[14]) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U14 ( .A(Fresh[4]), .B(
        SubCellInst_SboxInst_2_Q1), .Z(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U13 ( .A(Fresh[4]), .B(
        new_AGEMA_signal_1466), .Z(SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U10 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND1_U1_U8 ( .A(Fresh[4]), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U7 ( .A1(new_AGEMA_signal_1466), .A2(
        Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q1), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n8), .B(
        SubCellInst_SboxInst_2_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1554) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_n7), .B(
        SubCellInst_SboxInst_2_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T0) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_Q0), .B(SubCellInst_SboxInst_2_T0), .Z(
        SubCellInst_SboxInst_2_Q2) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1465), 
        .B(new_AGEMA_signal_1554), .Z(new_AGEMA_signal_1604) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U14 ( .A(Fresh[5]), .B(
        SubCellInst_SboxInst_2_Q4), .Z(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U13 ( .A(Fresh[5]), .B(
        new_AGEMA_signal_1467), .Z(SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U10 ( .A1(Ciphertext_s1[10]), .A2(
        SubCellInst_SboxInst_2_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_2_n3), 
        .A2(SubCellInst_SboxInst_2_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND3_U1_U8 ( .A(Fresh[5]), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U7 ( .A1(new_AGEMA_signal_1467), .A2(
        Ciphertext_s1[10]), .ZN(SubCellInst_SboxInst_2_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q4), 
        .A2(SubCellInst_SboxInst_2_n3), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n8), .B(
        SubCellInst_SboxInst_2_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1555) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_n7), .B(
        SubCellInst_SboxInst_2_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T2) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[10]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L1), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_Q7) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1556), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1605) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_2_), .B(SubCellInst_SboxInst_2_T0), .Z(
        SubCellInst_SboxInst_2_L3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1181), 
        .B(new_AGEMA_signal_1554), .Z(new_AGEMA_signal_1606) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L3), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1606), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1728) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_XX_1_), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1179), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1668) );
  INV_X1 SubCellInst_SboxInst_3_U3_U1 ( .A(SubCellInst_SboxInst_3_YY_1_), .ZN(
        ShiftRowsOutput[3]) );
  INV_X1 SubCellInst_SboxInst_3_U2_U1 ( .A(SubCellInst_SboxInst_3_YY_0_), .ZN(
        ShiftRowsOutput[2]) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U14 ( .A(Fresh[6]), .B(
        SubCellInst_SboxInst_3_Q1), .Z(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U13 ( .A(Fresh[6]), .B(
        new_AGEMA_signal_1472), .Z(SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U10 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND1_U1_U8 ( .A(Fresh[6]), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U7 ( .A1(new_AGEMA_signal_1472), .A2(
        Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q1), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n8), .B(
        SubCellInst_SboxInst_3_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1557) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_n7), .B(
        SubCellInst_SboxInst_3_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T0) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_Q0), .B(SubCellInst_SboxInst_3_T0), .Z(
        SubCellInst_SboxInst_3_Q2) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1471), 
        .B(new_AGEMA_signal_1557), .Z(new_AGEMA_signal_1608) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U14 ( .A(Fresh[7]), .B(
        SubCellInst_SboxInst_3_Q4), .Z(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U13 ( .A(Fresh[7]), .B(
        new_AGEMA_signal_1473), .Z(SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U10 ( .A1(Ciphertext_s1[14]), .A2(
        SubCellInst_SboxInst_3_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_3_n3), 
        .A2(SubCellInst_SboxInst_3_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND3_U1_U8 ( .A(Fresh[7]), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U7 ( .A1(new_AGEMA_signal_1473), .A2(
        Ciphertext_s1[14]), .ZN(SubCellInst_SboxInst_3_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q4), 
        .A2(SubCellInst_SboxInst_3_n3), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n8), .B(
        SubCellInst_SboxInst_3_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1558) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_n7), .B(
        SubCellInst_SboxInst_3_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T2) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[14]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L1), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_Q7) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1559), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1609) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_2_), .B(SubCellInst_SboxInst_3_T0), .Z(
        SubCellInst_SboxInst_3_L3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1187), 
        .B(new_AGEMA_signal_1557), .Z(new_AGEMA_signal_1610) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L3), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1610), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1730) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_XX_1_), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1185), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1672) );
  INV_X1 SubCellInst_SboxInst_4_U3_U1 ( .A(SubCellInst_SboxInst_4_YY_1_), .ZN(
        ShiftRowsOutput[27]) );
  INV_X1 SubCellInst_SboxInst_4_U2_U1 ( .A(SubCellInst_SboxInst_4_YY_0_), .ZN(
        ShiftRowsOutput[26]) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U14 ( .A(Fresh[8]), .B(
        SubCellInst_SboxInst_4_Q1), .Z(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U13 ( .A(Fresh[8]), .B(
        new_AGEMA_signal_1478), .Z(SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U10 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND1_U1_U8 ( .A(Fresh[8]), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U7 ( .A1(new_AGEMA_signal_1478), .A2(
        Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q1), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n8), .B(
        SubCellInst_SboxInst_4_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1560) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_n7), .B(
        SubCellInst_SboxInst_4_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T0) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_Q0), .B(SubCellInst_SboxInst_4_T0), .Z(
        SubCellInst_SboxInst_4_Q2) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1477), 
        .B(new_AGEMA_signal_1560), .Z(new_AGEMA_signal_1612) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U14 ( .A(Fresh[9]), .B(
        SubCellInst_SboxInst_4_Q4), .Z(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U13 ( .A(Fresh[9]), .B(
        new_AGEMA_signal_1479), .Z(SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U10 ( .A1(Ciphertext_s1[18]), .A2(
        SubCellInst_SboxInst_4_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_4_n3), 
        .A2(SubCellInst_SboxInst_4_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND3_U1_U8 ( .A(Fresh[9]), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U7 ( .A1(new_AGEMA_signal_1479), .A2(
        Ciphertext_s1[18]), .ZN(SubCellInst_SboxInst_4_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q4), 
        .A2(SubCellInst_SboxInst_4_n3), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n8), .B(
        SubCellInst_SboxInst_4_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1561) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_n7), .B(
        SubCellInst_SboxInst_4_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T2) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[18]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L1), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_Q7) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1562), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1613) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_2_), .B(SubCellInst_SboxInst_4_T0), .Z(
        SubCellInst_SboxInst_4_L3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1193), 
        .B(new_AGEMA_signal_1560), .Z(new_AGEMA_signal_1614) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L3), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1614), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1732) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_XX_1_), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1191), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1676) );
  INV_X1 SubCellInst_SboxInst_5_U3_U1 ( .A(SubCellInst_SboxInst_5_YY_1_), .ZN(
        ShiftRowsOutput[31]) );
  INV_X1 SubCellInst_SboxInst_5_U2_U1 ( .A(SubCellInst_SboxInst_5_YY_0_), .ZN(
        ShiftRowsOutput[30]) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U14 ( .A(Fresh[10]), .B(
        SubCellInst_SboxInst_5_Q1), .Z(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U13 ( .A(Fresh[10]), .B(
        new_AGEMA_signal_1484), .Z(SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U10 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND1_U1_U8 ( .A(Fresh[10]), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U7 ( .A1(new_AGEMA_signal_1484), .A2(
        Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q1), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n8), .B(
        SubCellInst_SboxInst_5_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1563) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_n7), .B(
        SubCellInst_SboxInst_5_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T0) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_Q0), .B(SubCellInst_SboxInst_5_T0), .Z(
        SubCellInst_SboxInst_5_Q2) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1483), 
        .B(new_AGEMA_signal_1563), .Z(new_AGEMA_signal_1616) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U14 ( .A(Fresh[11]), .B(
        SubCellInst_SboxInst_5_Q4), .Z(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U13 ( .A(Fresh[11]), .B(
        new_AGEMA_signal_1485), .Z(SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U10 ( .A1(Ciphertext_s1[22]), .A2(
        SubCellInst_SboxInst_5_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_5_n3), 
        .A2(SubCellInst_SboxInst_5_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND3_U1_U8 ( .A(Fresh[11]), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U7 ( .A1(new_AGEMA_signal_1485), .A2(
        Ciphertext_s1[22]), .ZN(SubCellInst_SboxInst_5_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q4), 
        .A2(SubCellInst_SboxInst_5_n3), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n8), .B(
        SubCellInst_SboxInst_5_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1564) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_n7), .B(
        SubCellInst_SboxInst_5_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T2) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[22]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L1), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_Q7) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1565), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1617) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_2_), .B(SubCellInst_SboxInst_5_T0), .Z(
        SubCellInst_SboxInst_5_L3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1199), 
        .B(new_AGEMA_signal_1563), .Z(new_AGEMA_signal_1618) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L3), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1618), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1734) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_XX_1_), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1197), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1680) );
  INV_X1 SubCellInst_SboxInst_6_U3_U1 ( .A(SubCellInst_SboxInst_6_YY_1_), .ZN(
        ShiftRowsOutput[19]) );
  INV_X1 SubCellInst_SboxInst_6_U2_U1 ( .A(SubCellInst_SboxInst_6_YY_0_), .ZN(
        ShiftRowsOutput[18]) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U14 ( .A(Fresh[12]), .B(
        SubCellInst_SboxInst_6_Q1), .Z(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U13 ( .A(Fresh[12]), .B(
        new_AGEMA_signal_1490), .Z(SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U10 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND1_U1_U8 ( .A(Fresh[12]), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U7 ( .A1(new_AGEMA_signal_1490), .A2(
        Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q1), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n8), .B(
        SubCellInst_SboxInst_6_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1566) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_n7), .B(
        SubCellInst_SboxInst_6_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T0) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_Q0), .B(SubCellInst_SboxInst_6_T0), .Z(
        SubCellInst_SboxInst_6_Q2) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1489), 
        .B(new_AGEMA_signal_1566), .Z(new_AGEMA_signal_1620) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U14 ( .A(Fresh[13]), .B(
        SubCellInst_SboxInst_6_Q4), .Z(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U13 ( .A(Fresh[13]), .B(
        new_AGEMA_signal_1491), .Z(SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U10 ( .A1(Ciphertext_s1[26]), .A2(
        SubCellInst_SboxInst_6_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_6_n3), 
        .A2(SubCellInst_SboxInst_6_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND3_U1_U8 ( .A(Fresh[13]), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U7 ( .A1(new_AGEMA_signal_1491), .A2(
        Ciphertext_s1[26]), .ZN(SubCellInst_SboxInst_6_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q4), 
        .A2(SubCellInst_SboxInst_6_n3), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n8), .B(
        SubCellInst_SboxInst_6_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1567) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_n7), .B(
        SubCellInst_SboxInst_6_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T2) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[26]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L1), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_Q7) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1568), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1621) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_2_), .B(SubCellInst_SboxInst_6_T0), .Z(
        SubCellInst_SboxInst_6_L3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1205), 
        .B(new_AGEMA_signal_1566), .Z(new_AGEMA_signal_1622) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L3), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1622), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1736) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_XX_1_), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1203), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1684) );
  INV_X1 SubCellInst_SboxInst_7_U3_U1 ( .A(SubCellInst_SboxInst_7_YY_1_), .ZN(
        ShiftRowsOutput[23]) );
  INV_X1 SubCellInst_SboxInst_7_U2_U1 ( .A(SubCellInst_SboxInst_7_YY_0_), .ZN(
        ShiftRowsOutput[22]) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U14 ( .A(Fresh[14]), .B(
        SubCellInst_SboxInst_7_Q1), .Z(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U13 ( .A(Fresh[14]), .B(
        new_AGEMA_signal_1496), .Z(SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U10 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND1_U1_U8 ( .A(Fresh[14]), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U7 ( .A1(new_AGEMA_signal_1496), .A2(
        Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q1), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n8), .B(
        SubCellInst_SboxInst_7_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1569) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_n7), .B(
        SubCellInst_SboxInst_7_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T0) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_Q0), .B(SubCellInst_SboxInst_7_T0), .Z(
        SubCellInst_SboxInst_7_Q2) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1495), 
        .B(new_AGEMA_signal_1569), .Z(new_AGEMA_signal_1624) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U14 ( .A(Fresh[15]), .B(
        SubCellInst_SboxInst_7_Q4), .Z(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U13 ( .A(Fresh[15]), .B(
        new_AGEMA_signal_1497), .Z(SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U10 ( .A1(Ciphertext_s1[30]), .A2(
        SubCellInst_SboxInst_7_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_7_n3), 
        .A2(SubCellInst_SboxInst_7_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND3_U1_U8 ( .A(Fresh[15]), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U7 ( .A1(new_AGEMA_signal_1497), .A2(
        Ciphertext_s1[30]), .ZN(SubCellInst_SboxInst_7_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q4), 
        .A2(SubCellInst_SboxInst_7_n3), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n8), .B(
        SubCellInst_SboxInst_7_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1570) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_n7), .B(
        SubCellInst_SboxInst_7_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T2) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[30]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L1), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_Q7) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1571), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1625) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_2_), .B(SubCellInst_SboxInst_7_T0), .Z(
        SubCellInst_SboxInst_7_L3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1211), 
        .B(new_AGEMA_signal_1569), .Z(new_AGEMA_signal_1626) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L3), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1626), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1738) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_XX_1_), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1209), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1688) );
  INV_X1 SubCellInst_SboxInst_8_U3_U1 ( .A(SubCellInst_SboxInst_8_YY_1_), .ZN(
        AddRoundConstantOutput[35]) );
  INV_X1 SubCellInst_SboxInst_8_U2_U1 ( .A(SubCellInst_SboxInst_8_YY_0_), .ZN(
        AddRoundConstantOutput[34]) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U14 ( .A(Fresh[16]), .B(
        SubCellInst_SboxInst_8_Q1), .Z(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U13 ( .A(Fresh[16]), .B(
        new_AGEMA_signal_1502), .Z(SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U10 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND1_U1_U8 ( .A(Fresh[16]), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U7 ( .A1(new_AGEMA_signal_1502), .A2(
        Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q1), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n8), .B(
        SubCellInst_SboxInst_8_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1572) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_n7), .B(
        SubCellInst_SboxInst_8_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T0) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_Q0), .B(SubCellInst_SboxInst_8_T0), .Z(
        SubCellInst_SboxInst_8_Q2) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1501), 
        .B(new_AGEMA_signal_1572), .Z(new_AGEMA_signal_1628) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U14 ( .A(Fresh[17]), .B(
        SubCellInst_SboxInst_8_Q4), .Z(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U13 ( .A(Fresh[17]), .B(
        new_AGEMA_signal_1503), .Z(SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U10 ( .A1(Ciphertext_s1[34]), .A2(
        SubCellInst_SboxInst_8_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_8_n3), 
        .A2(SubCellInst_SboxInst_8_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND3_U1_U8 ( .A(Fresh[17]), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U7 ( .A1(new_AGEMA_signal_1503), .A2(
        Ciphertext_s1[34]), .ZN(SubCellInst_SboxInst_8_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q4), 
        .A2(SubCellInst_SboxInst_8_n3), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n8), .B(
        SubCellInst_SboxInst_8_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1573) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_n7), .B(
        SubCellInst_SboxInst_8_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T2) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[34]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L1), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_Q7) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1574), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1629) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_2_), .B(SubCellInst_SboxInst_8_T0), .Z(
        SubCellInst_SboxInst_8_L3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1217), 
        .B(new_AGEMA_signal_1572), .Z(new_AGEMA_signal_1630) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L3), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1630), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1740) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_XX_1_), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1215), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1692) );
  INV_X1 SubCellInst_SboxInst_9_U3_U1 ( .A(SubCellInst_SboxInst_9_YY_1_), .ZN(
        AddRoundConstantOutput[39]) );
  INV_X1 SubCellInst_SboxInst_9_U2_U1 ( .A(SubCellInst_SboxInst_9_YY_0_), .ZN(
        AddRoundConstantOutput[38]) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U14 ( .A(Fresh[18]), .B(
        SubCellInst_SboxInst_9_Q1), .Z(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U13 ( .A(Fresh[18]), .B(
        new_AGEMA_signal_1508), .Z(SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U10 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND1_U1_U8 ( .A(Fresh[18]), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U7 ( .A1(new_AGEMA_signal_1508), .A2(
        Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q1), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n8), .B(
        SubCellInst_SboxInst_9_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1575) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_n7), .B(
        SubCellInst_SboxInst_9_AND1_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T0) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_Q0), .B(SubCellInst_SboxInst_9_T0), .Z(
        SubCellInst_SboxInst_9_Q2) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1507), 
        .B(new_AGEMA_signal_1575), .Z(new_AGEMA_signal_1632) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U14 ( .A(Fresh[19]), .B(
        SubCellInst_SboxInst_9_Q4), .Z(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U13 ( .A(Fresh[19]), .B(
        new_AGEMA_signal_1509), .Z(SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U10 ( .A1(Ciphertext_s1[38]), .A2(
        SubCellInst_SboxInst_9_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_9_n3), 
        .A2(SubCellInst_SboxInst_9_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND3_U1_U8 ( .A(Fresh[19]), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U7 ( .A1(new_AGEMA_signal_1509), .A2(
        Ciphertext_s1[38]), .ZN(SubCellInst_SboxInst_9_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q4), 
        .A2(SubCellInst_SboxInst_9_n3), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n8), .B(
        SubCellInst_SboxInst_9_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1576) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_n7), .B(
        SubCellInst_SboxInst_9_AND3_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T2) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[38]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L1), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_Q7) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1577), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1633) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_2_), .B(SubCellInst_SboxInst_9_T0), .Z(
        SubCellInst_SboxInst_9_L3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1223), 
        .B(new_AGEMA_signal_1575), .Z(new_AGEMA_signal_1634) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L3), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1634), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1742) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_XX_1_), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1221), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1696) );
  INV_X1 SubCellInst_SboxInst_10_U3_U1 ( .A(SubCellInst_SboxInst_10_YY_1_), 
        .ZN(AddRoundConstantOutput[43]) );
  INV_X1 SubCellInst_SboxInst_10_U2_U1 ( .A(SubCellInst_SboxInst_10_YY_0_), 
        .ZN(AddRoundConstantOutput[42]) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U14 ( .A(Fresh[20]), .B(
        SubCellInst_SboxInst_10_Q1), .Z(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U13 ( .A(Fresh[20]), .B(
        new_AGEMA_signal_1514), .Z(SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U10 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_10_n3), 
        .A2(SubCellInst_SboxInst_10_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND1_U1_U8 ( .A(Fresh[20]), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U7 ( .A1(new_AGEMA_signal_1514), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q1), 
        .A2(SubCellInst_SboxInst_10_n3), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n8), .B(
        SubCellInst_SboxInst_10_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1578)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_n7), .B(
        SubCellInst_SboxInst_10_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T0) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_Q0), .B(SubCellInst_SboxInst_10_T0), .Z(
        SubCellInst_SboxInst_10_Q2) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1513), 
        .B(new_AGEMA_signal_1578), .Z(new_AGEMA_signal_1636) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U14 ( .A(Fresh[21]), .B(
        SubCellInst_SboxInst_10_Q4), .Z(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U13 ( .A(Fresh[21]), .B(
        new_AGEMA_signal_1515), .Z(SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U10 ( .A1(Ciphertext_s1[42]), .A2(
        SubCellInst_SboxInst_10_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_10_n3), 
        .A2(SubCellInst_SboxInst_10_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND3_U1_U8 ( .A(Fresh[21]), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U7 ( .A1(new_AGEMA_signal_1515), 
        .A2(Ciphertext_s1[42]), .ZN(SubCellInst_SboxInst_10_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q4), 
        .A2(SubCellInst_SboxInst_10_n3), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n8), .B(
        SubCellInst_SboxInst_10_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1579)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_n7), .B(
        SubCellInst_SboxInst_10_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T2) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[42]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L1), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_Q7) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1580), 
        .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1637) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_2_), .B(SubCellInst_SboxInst_10_T0), .Z(
        SubCellInst_SboxInst_10_L3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1229), .B(new_AGEMA_signal_1578), .Z(new_AGEMA_signal_1638) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L3), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1638), .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1744) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_XX_1_), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1227), .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1700) );
  INV_X1 SubCellInst_SboxInst_11_U3_U1 ( .A(SubCellInst_SboxInst_11_YY_1_), 
        .ZN(SubCellOutput_47) );
  INV_X1 SubCellInst_SboxInst_11_U2_U1 ( .A(SubCellInst_SboxInst_11_YY_0_), 
        .ZN(SubCellOutput_46) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U14 ( .A(Fresh[22]), .B(
        SubCellInst_SboxInst_11_Q1), .Z(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U13 ( .A(Fresh[22]), .B(
        new_AGEMA_signal_1520), .Z(SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U10 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_11_n3), 
        .A2(SubCellInst_SboxInst_11_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND1_U1_U8 ( .A(Fresh[22]), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U7 ( .A1(new_AGEMA_signal_1520), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q1), 
        .A2(SubCellInst_SboxInst_11_n3), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n8), .B(
        SubCellInst_SboxInst_11_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1581)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_n7), .B(
        SubCellInst_SboxInst_11_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T0) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_Q0), .B(SubCellInst_SboxInst_11_T0), .Z(
        SubCellInst_SboxInst_11_Q2) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1519), 
        .B(new_AGEMA_signal_1581), .Z(new_AGEMA_signal_1640) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U14 ( .A(Fresh[23]), .B(
        SubCellInst_SboxInst_11_Q4), .Z(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U13 ( .A(Fresh[23]), .B(
        new_AGEMA_signal_1521), .Z(SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U10 ( .A1(Ciphertext_s1[46]), .A2(
        SubCellInst_SboxInst_11_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_11_n3), 
        .A2(SubCellInst_SboxInst_11_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND3_U1_U8 ( .A(Fresh[23]), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U7 ( .A1(new_AGEMA_signal_1521), 
        .A2(Ciphertext_s1[46]), .ZN(SubCellInst_SboxInst_11_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q4), 
        .A2(SubCellInst_SboxInst_11_n3), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n8), .B(
        SubCellInst_SboxInst_11_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1582)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_n7), .B(
        SubCellInst_SboxInst_11_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T2) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[46]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L1), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_Q7) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1583), 
        .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1641) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_2_), .B(SubCellInst_SboxInst_11_T0), .Z(
        SubCellInst_SboxInst_11_L3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1235), .B(new_AGEMA_signal_1581), .Z(new_AGEMA_signal_1642) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L3), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1642), .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1746) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_XX_1_), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1233), .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1704) );
  INV_X1 SubCellInst_SboxInst_12_U3_U1 ( .A(SubCellInst_SboxInst_12_YY_1_), 
        .ZN(AddRoundConstantOutput[51]) );
  INV_X1 SubCellInst_SboxInst_12_U2_U1 ( .A(SubCellInst_SboxInst_12_YY_0_), 
        .ZN(AddRoundConstantOutput[50]) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U14 ( .A(Fresh[24]), .B(
        SubCellInst_SboxInst_12_Q1), .Z(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U13 ( .A(Fresh[24]), .B(
        new_AGEMA_signal_1526), .Z(SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U10 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_12_n3), 
        .A2(SubCellInst_SboxInst_12_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND1_U1_U8 ( .A(Fresh[24]), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U7 ( .A1(new_AGEMA_signal_1526), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q1), 
        .A2(SubCellInst_SboxInst_12_n3), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n8), .B(
        SubCellInst_SboxInst_12_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1584)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_n7), .B(
        SubCellInst_SboxInst_12_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T0) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_Q0), .B(SubCellInst_SboxInst_12_T0), .Z(
        SubCellInst_SboxInst_12_Q2) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1525), 
        .B(new_AGEMA_signal_1584), .Z(new_AGEMA_signal_1644) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U14 ( .A(Fresh[25]), .B(
        SubCellInst_SboxInst_12_Q4), .Z(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U13 ( .A(Fresh[25]), .B(
        new_AGEMA_signal_1527), .Z(SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U10 ( .A1(Ciphertext_s1[50]), .A2(
        SubCellInst_SboxInst_12_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_12_n3), 
        .A2(SubCellInst_SboxInst_12_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND3_U1_U8 ( .A(Fresh[25]), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U7 ( .A1(new_AGEMA_signal_1527), 
        .A2(Ciphertext_s1[50]), .ZN(SubCellInst_SboxInst_12_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q4), 
        .A2(SubCellInst_SboxInst_12_n3), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n8), .B(
        SubCellInst_SboxInst_12_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1585)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_n7), .B(
        SubCellInst_SboxInst_12_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T2) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[50]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L1), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_Q7) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1586), 
        .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1645) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_2_), .B(SubCellInst_SboxInst_12_T0), .Z(
        SubCellInst_SboxInst_12_L3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1241), .B(new_AGEMA_signal_1584), .Z(new_AGEMA_signal_1646) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L3), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1646), .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1748) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_XX_1_), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1239), .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1708) );
  INV_X1 SubCellInst_SboxInst_13_U3_U1 ( .A(SubCellInst_SboxInst_13_YY_1_), 
        .ZN(AddRoundConstantOutput[55]) );
  INV_X1 SubCellInst_SboxInst_13_U2_U1 ( .A(SubCellInst_SboxInst_13_YY_0_), 
        .ZN(AddRoundConstantOutput[54]) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U14 ( .A(Fresh[26]), .B(
        SubCellInst_SboxInst_13_Q1), .Z(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U13 ( .A(Fresh[26]), .B(
        new_AGEMA_signal_1532), .Z(SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U10 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_13_n3), 
        .A2(SubCellInst_SboxInst_13_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND1_U1_U8 ( .A(Fresh[26]), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U7 ( .A1(new_AGEMA_signal_1532), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q1), 
        .A2(SubCellInst_SboxInst_13_n3), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n8), .B(
        SubCellInst_SboxInst_13_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1587)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_n7), .B(
        SubCellInst_SboxInst_13_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T0) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_Q0), .B(SubCellInst_SboxInst_13_T0), .Z(
        SubCellInst_SboxInst_13_Q2) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1531), 
        .B(new_AGEMA_signal_1587), .Z(new_AGEMA_signal_1648) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U14 ( .A(Fresh[27]), .B(
        SubCellInst_SboxInst_13_Q4), .Z(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U13 ( .A(Fresh[27]), .B(
        new_AGEMA_signal_1533), .Z(SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U10 ( .A1(Ciphertext_s1[54]), .A2(
        SubCellInst_SboxInst_13_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_13_n3), 
        .A2(SubCellInst_SboxInst_13_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND3_U1_U8 ( .A(Fresh[27]), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U7 ( .A1(new_AGEMA_signal_1533), 
        .A2(Ciphertext_s1[54]), .ZN(SubCellInst_SboxInst_13_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q4), 
        .A2(SubCellInst_SboxInst_13_n3), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n8), .B(
        SubCellInst_SboxInst_13_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1588)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_n7), .B(
        SubCellInst_SboxInst_13_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T2) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[54]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L1), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_Q7) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1589), 
        .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1649) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_2_), .B(SubCellInst_SboxInst_13_T0), .Z(
        SubCellInst_SboxInst_13_L3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1247), .B(new_AGEMA_signal_1587), .Z(new_AGEMA_signal_1650) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L3), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1650), .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1750) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_XX_1_), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1245), .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1712) );
  INV_X1 SubCellInst_SboxInst_14_U3_U1 ( .A(SubCellInst_SboxInst_14_YY_1_), 
        .ZN(AddRoundConstantOutput[59]) );
  INV_X1 SubCellInst_SboxInst_14_U2_U1 ( .A(SubCellInst_SboxInst_14_YY_0_), 
        .ZN(AddRoundConstantOutput[58]) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U14 ( .A(Fresh[28]), .B(
        SubCellInst_SboxInst_14_Q1), .Z(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U13 ( .A(Fresh[28]), .B(
        new_AGEMA_signal_1538), .Z(SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U10 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_14_n3), 
        .A2(SubCellInst_SboxInst_14_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND1_U1_U8 ( .A(Fresh[28]), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U7 ( .A1(new_AGEMA_signal_1538), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q1), 
        .A2(SubCellInst_SboxInst_14_n3), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n8), .B(
        SubCellInst_SboxInst_14_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1590)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_n7), .B(
        SubCellInst_SboxInst_14_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T0) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_Q0), .B(SubCellInst_SboxInst_14_T0), .Z(
        SubCellInst_SboxInst_14_Q2) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1537), 
        .B(new_AGEMA_signal_1590), .Z(new_AGEMA_signal_1652) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U14 ( .A(Fresh[29]), .B(
        SubCellInst_SboxInst_14_Q4), .Z(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U13 ( .A(Fresh[29]), .B(
        new_AGEMA_signal_1539), .Z(SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U10 ( .A1(Ciphertext_s1[58]), .A2(
        SubCellInst_SboxInst_14_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_14_n3), 
        .A2(SubCellInst_SboxInst_14_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND3_U1_U8 ( .A(Fresh[29]), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U7 ( .A1(new_AGEMA_signal_1539), 
        .A2(Ciphertext_s1[58]), .ZN(SubCellInst_SboxInst_14_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q4), 
        .A2(SubCellInst_SboxInst_14_n3), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n8), .B(
        SubCellInst_SboxInst_14_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1591)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_n7), .B(
        SubCellInst_SboxInst_14_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T2) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[58]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L1), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_Q7) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1592), 
        .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1653) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_2_), .B(SubCellInst_SboxInst_14_T0), .Z(
        SubCellInst_SboxInst_14_L3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1253), .B(new_AGEMA_signal_1590), .Z(new_AGEMA_signal_1654) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L3), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1654), .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1752) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_XX_1_), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1251), .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1716) );
  INV_X1 SubCellInst_SboxInst_15_U3_U1 ( .A(SubCellInst_SboxInst_15_YY_1_), 
        .ZN(SubCellOutput[63]) );
  INV_X1 SubCellInst_SboxInst_15_U2_U1 ( .A(SubCellInst_SboxInst_15_YY_0_), 
        .ZN(SubCellOutput[62]) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U14 ( .A(Fresh[30]), .B(
        SubCellInst_SboxInst_15_Q1), .Z(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U13 ( .A(Fresh[30]), .B(
        new_AGEMA_signal_1544), .Z(SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U10 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U9 ( .A1(SubCellInst_SboxInst_15_n3), 
        .A2(SubCellInst_SboxInst_15_AND1_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND1_U1_U8 ( .A(Fresh[30]), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U7 ( .A1(new_AGEMA_signal_1544), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND1_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND1_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q1), 
        .A2(SubCellInst_SboxInst_15_n3), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n8), .B(
        SubCellInst_SboxInst_15_AND1_U1_z_1__1_), .ZN(new_AGEMA_signal_1593)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_n7), .B(
        SubCellInst_SboxInst_15_AND1_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T0) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND1_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND1_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND1_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND1_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND1_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_Q0), .B(SubCellInst_SboxInst_15_T0), .Z(
        SubCellInst_SboxInst_15_Q2) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR2_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1543), 
        .B(new_AGEMA_signal_1593), .Z(new_AGEMA_signal_1656) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U14 ( .A(Fresh[31]), .B(
        SubCellInst_SboxInst_15_Q4), .Z(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U13 ( .A(Fresh[31]), .B(
        new_AGEMA_signal_1545), .Z(SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U10 ( .A1(Ciphertext_s1[62]), .A2(
        SubCellInst_SboxInst_15_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U9 ( .A1(SubCellInst_SboxInst_15_n3), 
        .A2(SubCellInst_SboxInst_15_AND3_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND3_U1_U8 ( .A(Fresh[31]), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U7 ( .A1(new_AGEMA_signal_1545), 
        .A2(Ciphertext_s1[62]), .ZN(SubCellInst_SboxInst_15_AND3_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND3_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q4), 
        .A2(SubCellInst_SboxInst_15_n3), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n8), .B(
        SubCellInst_SboxInst_15_AND3_U1_z_1__1_), .ZN(new_AGEMA_signal_1594)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_n7), .B(
        SubCellInst_SboxInst_15_AND3_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T2) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND3_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND3_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_n3), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[62]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND3_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND3_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND3_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L1), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_Q7) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR7_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1595), 
        .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1657) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_2_), .B(SubCellInst_SboxInst_15_T0), .Z(
        SubCellInst_SboxInst_15_L3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR11_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1259), .B(new_AGEMA_signal_1593), .Z(new_AGEMA_signal_1658) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L3), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_1_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1658), .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1754) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_XX_1_), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_YY_0_) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1257), .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1720) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_2_n1), .B(FSMUpdate[3]), .ZN(
        AddRoundConstantOutput[62]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1756), .B(1'b0), .Z(new_AGEMA_signal_1800) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[62]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1720), .Z(new_AGEMA_signal_1756) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_3_n1), .B(FSMUpdate[4]), .ZN(
        AddRoundConstantOutput[63]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1801), .B(1'b0), .Z(new_AGEMA_signal_1843) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[63]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1754), .Z(new_AGEMA_signal_1801) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_2_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[46]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1757), .B(1'b0), .Z(new_AGEMA_signal_1802) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_46), .ZN(AddConstXOR_AddConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1704), .Z(new_AGEMA_signal_1757) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_3_n1), .B(1'b0), .ZN(
        AddRoundConstantOutput[47]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1803), .B(1'b0), .Z(new_AGEMA_signal_1845) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_47), .ZN(AddConstXOR_AddConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1746), .Z(new_AGEMA_signal_1803) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_2_n1), .B(
        TweakeyGeneration_key_Feedback[2]), .ZN(ShiftRowsOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1758), .B(new_AGEMA_signal_1266), .Z(
        new_AGEMA_signal_1804) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[34]), .ZN(AddRoundTweakeyXOR_XORInst_0_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1692), .Z(new_AGEMA_signal_1758) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_3_n1), .B(
        TweakeyGeneration_key_Feedback[3]), .ZN(ShiftRowsOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1805), .B(new_AGEMA_signal_1269), .Z(
        new_AGEMA_signal_1847) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[35]), .ZN(AddRoundTweakeyXOR_XORInst_0_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1740), .Z(new_AGEMA_signal_1805) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_2_n1), .B(
        TweakeyGeneration_key_Feedback[6]), .ZN(ShiftRowsOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1759), .B(new_AGEMA_signal_1278), .Z(
        new_AGEMA_signal_1806) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[38]), .ZN(AddRoundTweakeyXOR_XORInst_1_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1696), .Z(new_AGEMA_signal_1759) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_3_n1), .B(
        TweakeyGeneration_key_Feedback[7]), .ZN(ShiftRowsOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1807), .B(new_AGEMA_signal_1281), .Z(
        new_AGEMA_signal_1849) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[39]), .ZN(AddRoundTweakeyXOR_XORInst_1_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1742), .Z(new_AGEMA_signal_1807) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_2_n1), .B(
        TweakeyGeneration_key_Feedback[10]), .ZN(ShiftRowsOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1760), .B(new_AGEMA_signal_1290), .Z(
        new_AGEMA_signal_1808) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[42]), .ZN(AddRoundTweakeyXOR_XORInst_2_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1700), .Z(new_AGEMA_signal_1760) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_3_n1), .B(
        TweakeyGeneration_key_Feedback[11]), .ZN(ShiftRowsOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1809), .B(new_AGEMA_signal_1293), .Z(
        new_AGEMA_signal_1851) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[43]), .ZN(AddRoundTweakeyXOR_XORInst_2_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1744), .Z(new_AGEMA_signal_1809) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_2_n1), .B(
        TweakeyGeneration_key_Feedback[14]), .ZN(ShiftRowsOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1852), .B(new_AGEMA_signal_1302), .Z(
        new_AGEMA_signal_1890) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[46]), .ZN(AddRoundTweakeyXOR_XORInst_3_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1802), .Z(new_AGEMA_signal_1852) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_3_n1), .B(
        TweakeyGeneration_key_Feedback[15]), .ZN(ShiftRowsOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1891), .B(new_AGEMA_signal_1305), .Z(
        new_AGEMA_signal_1953) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[47]), .ZN(AddRoundTweakeyXOR_XORInst_3_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1845), .Z(new_AGEMA_signal_1891) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_2_n1), .B(
        TweakeyGeneration_key_Feedback[18]), .ZN(MCOutput[34]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1761), .B(new_AGEMA_signal_1314), .Z(
        new_AGEMA_signal_1810) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[50]), .ZN(AddRoundTweakeyXOR_XORInst_4_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1708), .Z(new_AGEMA_signal_1761) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_3_n1), .B(
        TweakeyGeneration_key_Feedback[19]), .ZN(MCOutput[35]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1811), .B(new_AGEMA_signal_1317), .Z(
        new_AGEMA_signal_1854) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[51]), .ZN(AddRoundTweakeyXOR_XORInst_4_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1748), .Z(new_AGEMA_signal_1811) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_2_n1), .B(
        TweakeyGeneration_key_Feedback[22]), .ZN(MCOutput[38]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1762), .B(new_AGEMA_signal_1326), .Z(
        new_AGEMA_signal_1812) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[54]), .ZN(AddRoundTweakeyXOR_XORInst_5_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1712), .Z(new_AGEMA_signal_1762) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_3_n1), .B(
        TweakeyGeneration_key_Feedback[23]), .ZN(MCOutput[39]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1813), .B(new_AGEMA_signal_1329), .Z(
        new_AGEMA_signal_1856) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[55]), .ZN(AddRoundTweakeyXOR_XORInst_5_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1750), .Z(new_AGEMA_signal_1813) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_2_n1), .B(
        TweakeyGeneration_key_Feedback[26]), .ZN(MCOutput[42]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1763), .B(new_AGEMA_signal_1338), .Z(
        new_AGEMA_signal_1814) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[58]), .ZN(AddRoundTweakeyXOR_XORInst_6_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1716), .Z(new_AGEMA_signal_1763) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_3_n1), .B(
        TweakeyGeneration_key_Feedback[27]), .ZN(MCOutput[43]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1815), .B(new_AGEMA_signal_1341), .Z(
        new_AGEMA_signal_1858) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[59]), .ZN(AddRoundTweakeyXOR_XORInst_6_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1752), .Z(new_AGEMA_signal_1815) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_2_n1), .B(
        TweakeyGeneration_key_Feedback[30]), .ZN(MCOutput[46]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1859), .B(new_AGEMA_signal_1350), .Z(
        new_AGEMA_signal_1898) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[62]), .ZN(AddRoundTweakeyXOR_XORInst_7_2_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1800), .Z(new_AGEMA_signal_1859) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_3_n1), .B(
        TweakeyGeneration_key_Feedback[31]), .ZN(MCOutput[47]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1899), .B(new_AGEMA_signal_1353), .Z(
        new_AGEMA_signal_1958) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[63]), .ZN(AddRoundTweakeyXOR_XORInst_7_3_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1843), .Z(new_AGEMA_signal_1899) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_2_n2), 
        .B(MCInst_MCR0_XORInst_0_2_n1), .ZN(MCOutput[50]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1861), .B(
        new_AGEMA_signal_1764), .Z(new_AGEMA_signal_1901) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[18]), .B(
        ShiftRowsOutput[2]), .ZN(MCInst_MCR0_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1684), .B(
        new_AGEMA_signal_1672), .Z(new_AGEMA_signal_1764) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .Z(MCInst_MCR0_XORInst_0_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1810), .Z(new_AGEMA_signal_1861) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_3_n2), 
        .B(MCInst_MCR0_XORInst_0_3_n1), .ZN(MCOutput[51]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1902), .B(
        new_AGEMA_signal_1816), .Z(new_AGEMA_signal_1960) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[19]), .B(
        ShiftRowsOutput[3]), .ZN(MCInst_MCR0_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1736), .B(
        new_AGEMA_signal_1730), .Z(new_AGEMA_signal_1816) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .Z(MCInst_MCR0_XORInst_0_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1854), .Z(new_AGEMA_signal_1902) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_2_n2), 
        .B(MCInst_MCR0_XORInst_1_2_n1), .ZN(MCOutput[54]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1863), .B(
        new_AGEMA_signal_1765), .Z(new_AGEMA_signal_1903) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[22]), .B(
        ShiftRowsOutput[6]), .ZN(MCInst_MCR0_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1688), .B(
        new_AGEMA_signal_1660), .Z(new_AGEMA_signal_1765) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .Z(MCInst_MCR0_XORInst_1_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1812), .Z(new_AGEMA_signal_1863) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_3_n2), 
        .B(MCInst_MCR0_XORInst_1_3_n1), .ZN(MCOutput[55]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1904), .B(
        new_AGEMA_signal_1817), .Z(new_AGEMA_signal_1963) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[23]), .B(
        ShiftRowsOutput[7]), .ZN(MCInst_MCR0_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1738), .B(
        new_AGEMA_signal_1724), .Z(new_AGEMA_signal_1817) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .Z(MCInst_MCR0_XORInst_1_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1856), .Z(new_AGEMA_signal_1904) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_2_n2), 
        .B(MCInst_MCR0_XORInst_2_2_n1), .ZN(MCOutput[58]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1865), .B(
        new_AGEMA_signal_1766), .Z(new_AGEMA_signal_1906) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[26]), .B(
        ShiftRowsOutput[10]), .ZN(MCInst_MCR0_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1676), .B(
        new_AGEMA_signal_1664), .Z(new_AGEMA_signal_1766) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .Z(MCInst_MCR0_XORInst_2_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1814), .Z(new_AGEMA_signal_1865) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_3_n2), 
        .B(MCInst_MCR0_XORInst_2_3_n1), .ZN(MCOutput[59]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1907), .B(
        new_AGEMA_signal_1818), .Z(new_AGEMA_signal_1965) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[27]), .B(
        ShiftRowsOutput[11]), .ZN(MCInst_MCR0_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1732), .B(
        new_AGEMA_signal_1726), .Z(new_AGEMA_signal_1818) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .Z(MCInst_MCR0_XORInst_2_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1858), .Z(new_AGEMA_signal_1907) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_2_n2), 
        .B(MCInst_MCR0_XORInst_3_2_n1), .ZN(MCOutput[62]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1966), .B(
        new_AGEMA_signal_1767), .Z(new_AGEMA_signal_2017) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins0_U1 ( .A(ShiftRowsOutput[30]), .B(
        ShiftRowsOutput[14]), .ZN(MCInst_MCR0_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1680), .B(
        new_AGEMA_signal_1668), .Z(new_AGEMA_signal_1767) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .Z(MCInst_MCR0_XORInst_3_2_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1898), .Z(new_AGEMA_signal_1966) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_3_n2), 
        .B(MCInst_MCR0_XORInst_3_3_n1), .ZN(MCOutput[63]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2018), .B(
        new_AGEMA_signal_1819), .Z(new_AGEMA_signal_2067) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins0_U1 ( .A(ShiftRowsOutput[31]), .B(
        ShiftRowsOutput[15]), .ZN(MCInst_MCR0_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1734), .B(
        new_AGEMA_signal_1728), .Z(new_AGEMA_signal_1819) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .Z(MCInst_MCR0_XORInst_3_3_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2018) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[18]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1867), .B(
        new_AGEMA_signal_1684), .Z(new_AGEMA_signal_1909) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[34]), .ZN(MCInst_MCR2_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1806), .Z(new_AGEMA_signal_1867) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[19]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1910), .B(
        new_AGEMA_signal_1736), .Z(new_AGEMA_signal_1968) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[35]), .ZN(MCInst_MCR2_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1849), .Z(new_AGEMA_signal_1910) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[22]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1868), .B(
        new_AGEMA_signal_1688), .Z(new_AGEMA_signal_1911) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[38]), .ZN(MCInst_MCR2_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1808), .Z(new_AGEMA_signal_1868) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[23]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1912), .B(
        new_AGEMA_signal_1738), .Z(new_AGEMA_signal_1970) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[39]), .ZN(MCInst_MCR2_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1851), .Z(new_AGEMA_signal_1912) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[26]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1971), .B(
        new_AGEMA_signal_1676), .Z(new_AGEMA_signal_2023) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[42]), .ZN(MCInst_MCR2_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1890), .Z(new_AGEMA_signal_1971) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[27]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2024), .B(
        new_AGEMA_signal_1732), .Z(new_AGEMA_signal_2071) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[43]), .ZN(MCInst_MCR2_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1953), .Z(new_AGEMA_signal_2024) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[30]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1869), .B(
        new_AGEMA_signal_1680), .Z(new_AGEMA_signal_1913) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[46]), .ZN(MCInst_MCR2_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1804), .Z(new_AGEMA_signal_1869) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[31]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1914), .B(
        new_AGEMA_signal_1734), .Z(new_AGEMA_signal_1973) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[47]), .ZN(MCInst_MCR2_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1847), .Z(new_AGEMA_signal_1914) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_2_n1), 
        .B(ShiftRowsOutput[18]), .ZN(MCOutput[2]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1870), .B(
        new_AGEMA_signal_1684), .Z(new_AGEMA_signal_1915) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[34]), 
        .ZN(MCInst_MCR3_XORInst_0_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1810), .Z(new_AGEMA_signal_1870) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_3_n1), 
        .B(ShiftRowsOutput[19]), .ZN(MCOutput[3]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1916), .B(
        new_AGEMA_signal_1736), .Z(new_AGEMA_signal_1975) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[35]), 
        .ZN(MCInst_MCR3_XORInst_0_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1854), .Z(new_AGEMA_signal_1916) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_2_n1), 
        .B(ShiftRowsOutput[22]), .ZN(MCOutput[6]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1871), .B(
        new_AGEMA_signal_1688), .Z(new_AGEMA_signal_1917) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[38]), 
        .ZN(MCInst_MCR3_XORInst_1_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1812), .Z(new_AGEMA_signal_1871) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_3_n1), 
        .B(ShiftRowsOutput[23]), .ZN(MCOutput[7]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1918), .B(
        new_AGEMA_signal_1738), .Z(new_AGEMA_signal_1977) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[39]), 
        .ZN(MCInst_MCR3_XORInst_1_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1856), .Z(new_AGEMA_signal_1918) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_2_n1), 
        .B(ShiftRowsOutput[26]), .ZN(MCOutput[10]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1872), .B(
        new_AGEMA_signal_1676), .Z(new_AGEMA_signal_1919) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[42]), 
        .ZN(MCInst_MCR3_XORInst_2_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1814), .Z(new_AGEMA_signal_1872) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_3_n1), 
        .B(ShiftRowsOutput[27]), .ZN(MCOutput[11]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1920), .B(
        new_AGEMA_signal_1732), .Z(new_AGEMA_signal_1979) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[43]), 
        .ZN(MCInst_MCR3_XORInst_2_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1858), .Z(new_AGEMA_signal_1920) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_2_n1), 
        .B(ShiftRowsOutput[30]), .ZN(MCOutput[14]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1980), .B(
        new_AGEMA_signal_1680), .Z(new_AGEMA_signal_2033) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[46]), 
        .ZN(MCInst_MCR3_XORInst_3_2_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_2_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1898), .Z(new_AGEMA_signal_1980) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_3_n1), 
        .B(ShiftRowsOutput[31]), .ZN(MCOutput[15]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2034), .B(
        new_AGEMA_signal_1734), .Z(new_AGEMA_signal_2077) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[47]), 
        .ZN(MCInst_MCR3_XORInst_3_3_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_3_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1958), .Z(new_AGEMA_signal_2034) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_0_U1 ( .A(MCOutput[0]), .B(
        Plaintext_s0[0]), .S(rst), .Z(StateRegInput[0]) );
  MUX2_X1 PlaintextMUX_MUXInst_0_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2027), .B(
        Plaintext_s1[0]), .S(rst), .Z(new_AGEMA_signal_2036) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_0_U1 ( .A(MCOutput[1]), .B(
        Plaintext_s0[1]), .S(rst), .Z(StateRegInput[1]) );
  MUX2_X1 PlaintextMUX_MUXInst_1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2073), .B(
        Plaintext_s1[1]), .S(rst), .Z(new_AGEMA_signal_2079) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_0_U1 ( .A(MCOutput[4]), .B(
        Plaintext_s0[4]), .S(rst), .Z(StateRegInput[4]) );
  MUX2_X1 PlaintextMUX_MUXInst_4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2029), .B(
        Plaintext_s1[4]), .S(rst), .Z(new_AGEMA_signal_2038) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_0_U1 ( .A(MCOutput[5]), .B(
        Plaintext_s0[5]), .S(rst), .Z(StateRegInput[5]) );
  MUX2_X1 PlaintextMUX_MUXInst_5_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2074), .B(
        Plaintext_s1[5]), .S(rst), .Z(new_AGEMA_signal_2081) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_0_U1 ( .A(MCOutput[8]), .B(
        Plaintext_s0[8]), .S(rst), .Z(StateRegInput[8]) );
  MUX2_X1 PlaintextMUX_MUXInst_8_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2031), .B(
        Plaintext_s1[8]), .S(rst), .Z(new_AGEMA_signal_2040) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_0_U1 ( .A(MCOutput[9]), .B(
        Plaintext_s0[9]), .S(rst), .Z(StateRegInput[9]) );
  MUX2_X1 PlaintextMUX_MUXInst_9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2075), .B(
        Plaintext_s1[9]), .S(rst), .Z(new_AGEMA_signal_2083) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_0_U1 ( .A(MCOutput[12]), .B(
        Plaintext_s0[12]), .S(rst), .Z(StateRegInput[12]) );
  MUX2_X1 PlaintextMUX_MUXInst_12_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2108), .B(
        Plaintext_s1[12]), .S(rst), .Z(new_AGEMA_signal_2111) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_0_U1 ( .A(MCOutput[13]), .B(
        Plaintext_s0[13]), .S(rst), .Z(StateRegInput[13]) );
  MUX2_X1 PlaintextMUX_MUXInst_13_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2118), .B(
        Plaintext_s1[13]), .S(rst), .Z(new_AGEMA_signal_2120) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_0_U1 ( .A(MCOutput[16]), .B(
        Plaintext_s0[16]), .S(rst), .Z(StateRegInput[16]) );
  MUX2_X1 PlaintextMUX_MUXInst_16_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2019), .B(
        Plaintext_s1[16]), .S(rst), .Z(new_AGEMA_signal_2044) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_0_U1 ( .A(MCOutput[17]), .B(
        Plaintext_s0[17]), .S(rst), .Z(StateRegInput[17]) );
  MUX2_X1 PlaintextMUX_MUXInst_17_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2068), .B(
        Plaintext_s1[17]), .S(rst), .Z(new_AGEMA_signal_2087) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_0_U1 ( .A(MCOutput[20]), .B(
        Plaintext_s0[20]), .S(rst), .Z(StateRegInput[20]) );
  MUX2_X1 PlaintextMUX_MUXInst_20_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2021), .B(
        Plaintext_s1[20]), .S(rst), .Z(new_AGEMA_signal_2046) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_0_U1 ( .A(MCOutput[21]), .B(
        Plaintext_s0[21]), .S(rst), .Z(StateRegInput[21]) );
  MUX2_X1 PlaintextMUX_MUXInst_21_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2069), .B(
        Plaintext_s1[21]), .S(rst), .Z(new_AGEMA_signal_2089) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_0_U1 ( .A(MCOutput[24]), .B(
        Plaintext_s0[24]), .S(rst), .Z(StateRegInput[24]) );
  MUX2_X1 PlaintextMUX_MUXInst_24_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2106), .B(
        Plaintext_s1[24]), .S(rst), .Z(new_AGEMA_signal_2113) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_0_U1 ( .A(MCOutput[25]), .B(
        Plaintext_s0[25]), .S(rst), .Z(StateRegInput[25]) );
  MUX2_X1 PlaintextMUX_MUXInst_25_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2117), .B(
        Plaintext_s1[25]), .S(rst), .Z(new_AGEMA_signal_2122) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_0_U1 ( .A(MCOutput[28]), .B(
        Plaintext_s0[28]), .S(rst), .Z(StateRegInput[28]) );
  MUX2_X1 PlaintextMUX_MUXInst_28_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2025), .B(
        Plaintext_s1[28]), .S(rst), .Z(new_AGEMA_signal_2050) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_0_U1 ( .A(MCOutput[29]), .B(
        Plaintext_s0[29]), .S(rst), .Z(StateRegInput[29]) );
  MUX2_X1 PlaintextMUX_MUXInst_29_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2072), .B(
        Plaintext_s1[29]), .S(rst), .Z(new_AGEMA_signal_2093) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_0_U1 ( .A(MCOutput[32]), .B(
        Plaintext_s0[32]), .S(rst), .Z(StateRegInput[32]) );
  MUX2_X1 PlaintextMUX_MUXInst_32_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1892), .B(
        Plaintext_s1[32]), .S(rst), .Z(new_AGEMA_signal_1934) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_0_U1 ( .A(MCOutput[33]), .B(
        Plaintext_s0[33]), .S(rst), .Z(StateRegInput[33]) );
  MUX2_X1 PlaintextMUX_MUXInst_33_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1954), .B(
        Plaintext_s1[33]), .S(rst), .Z(new_AGEMA_signal_1994) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_0_U1 ( .A(MCOutput[36]), .B(
        Plaintext_s0[36]), .S(rst), .Z(StateRegInput[36]) );
  MUX2_X1 PlaintextMUX_MUXInst_36_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1894), .B(
        Plaintext_s1[36]), .S(rst), .Z(new_AGEMA_signal_1936) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_0_U1 ( .A(MCOutput[37]), .B(
        Plaintext_s0[37]), .S(rst), .Z(StateRegInput[37]) );
  MUX2_X1 PlaintextMUX_MUXInst_37_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1955), .B(
        Plaintext_s1[37]), .S(rst), .Z(new_AGEMA_signal_1996) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_0_U1 ( .A(MCOutput[40]), .B(
        Plaintext_s0[40]), .S(rst), .Z(StateRegInput[40]) );
  MUX2_X1 PlaintextMUX_MUXInst_40_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1896), .B(
        Plaintext_s1[40]), .S(rst), .Z(new_AGEMA_signal_1938) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_0_U1 ( .A(MCOutput[41]), .B(
        Plaintext_s0[41]), .S(rst), .Z(StateRegInput[41]) );
  MUX2_X1 PlaintextMUX_MUXInst_41_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1956), .B(
        Plaintext_s1[41]), .S(rst), .Z(new_AGEMA_signal_1998) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_0_U1 ( .A(MCOutput[44]), .B(
        Plaintext_s0[44]), .S(rst), .Z(StateRegInput[44]) );
  MUX2_X1 PlaintextMUX_MUXInst_44_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2009), .B(
        Plaintext_s1[44]), .S(rst), .Z(new_AGEMA_signal_2052) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_0_U1 ( .A(MCOutput[45]), .B(
        Plaintext_s0[45]), .S(rst), .Z(StateRegInput[45]) );
  MUX2_X1 PlaintextMUX_MUXInst_45_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2062), .B(
        Plaintext_s1[45]), .S(rst), .Z(new_AGEMA_signal_2095) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_0_U1 ( .A(MCOutput[48]), .B(
        Plaintext_s0[48]), .S(rst), .Z(StateRegInput[48]) );
  MUX2_X1 PlaintextMUX_MUXInst_48_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2011), .B(
        Plaintext_s1[48]), .S(rst), .Z(new_AGEMA_signal_2054) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_0_U1 ( .A(MCOutput[49]), .B(
        Plaintext_s0[49]), .S(rst), .Z(StateRegInput[49]) );
  MUX2_X1 PlaintextMUX_MUXInst_49_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2063), .B(
        Plaintext_s1[49]), .S(rst), .Z(new_AGEMA_signal_2097) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_0_U1 ( .A(MCOutput[52]), .B(
        Plaintext_s0[52]), .S(rst), .Z(StateRegInput[52]) );
  MUX2_X1 PlaintextMUX_MUXInst_52_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2013), .B(
        Plaintext_s1[52]), .S(rst), .Z(new_AGEMA_signal_2056) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_0_U1 ( .A(MCOutput[53]), .B(
        Plaintext_s0[53]), .S(rst), .Z(StateRegInput[53]) );
  MUX2_X1 PlaintextMUX_MUXInst_53_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2064), .B(
        Plaintext_s1[53]), .S(rst), .Z(new_AGEMA_signal_2099) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_0_U1 ( .A(MCOutput[56]), .B(
        Plaintext_s0[56]), .S(rst), .Z(StateRegInput[56]) );
  MUX2_X1 PlaintextMUX_MUXInst_56_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2015), .B(
        Plaintext_s1[56]), .S(rst), .Z(new_AGEMA_signal_2058) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_0_U1 ( .A(MCOutput[57]), .B(
        Plaintext_s0[57]), .S(rst), .Z(StateRegInput[57]) );
  MUX2_X1 PlaintextMUX_MUXInst_57_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2065), .B(
        Plaintext_s1[57]), .S(rst), .Z(new_AGEMA_signal_2101) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_0_U1 ( .A(MCOutput[60]), .B(
        Plaintext_s0[60]), .S(rst), .Z(StateRegInput[60]) );
  MUX2_X1 PlaintextMUX_MUXInst_60_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2104), .B(
        Plaintext_s1[60]), .S(rst), .Z(new_AGEMA_signal_2115) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_0_U1 ( .A(MCOutput[61]), .B(
        Plaintext_s0[61]), .S(rst), .Z(StateRegInput[61]) );
  MUX2_X1 PlaintextMUX_MUXInst_61_U1_Ins_1_U1 ( .A(new_AGEMA_signal_2116), .B(
        Plaintext_s1[61]), .S(rst), .Z(new_AGEMA_signal_2124) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U14 ( .A(Fresh[32]), .B(
        SubCellInst_SboxInst_0_Q2), .Z(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U13 ( .A(Fresh[32]), .B(
        new_AGEMA_signal_1596), .Z(SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U10 ( .A1(Ciphertext_s1[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U9 ( .A1(Ciphertext_s0[1]), .A2(
        SubCellInst_SboxInst_0_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND2_U1_U8 ( .A(Fresh[32]), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U7 ( .A1(new_AGEMA_signal_1596), .A2(
        Ciphertext_s1[1]), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q2), 
        .A2(Ciphertext_s0[1]), .ZN(SubCellInst_SboxInst_0_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n8), .B(
        SubCellInst_SboxInst_0_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1661) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_n7), .B(
        SubCellInst_SboxInst_0_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T1) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_T1), .B(SubCellInst_SboxInst_0_T2), .Z(
        SubCellInst_SboxInst_0_L0) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1661), 
        .B(new_AGEMA_signal_1549), .Z(new_AGEMA_signal_1725) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U14 ( .A(Fresh[33]), .B(
        SubCellInst_SboxInst_0_Q7), .Z(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U13 ( .A(Fresh[33]), .B(
        new_AGEMA_signal_1597), .Z(SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U10 ( .A1(new_AGEMA_signal_1456), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_0_Q6), 
        .A2(SubCellInst_SboxInst_0_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_0_AND4_U1_U8 ( .A(Fresh[33]), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U7 ( .A1(new_AGEMA_signal_1597), .A2(
        new_AGEMA_signal_1456), .ZN(SubCellInst_SboxInst_0_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_0_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_0_Q7), 
        .A2(SubCellInst_SboxInst_0_Q6), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n8), .B(
        SubCellInst_SboxInst_0_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1662) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_n7), .B(
        SubCellInst_SboxInst_0_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_0_T3) );
  XNOR2_X1 SubCellInst_SboxInst_0_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_0_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_0_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1456), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_0_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_0_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_L2), .Z(
        SubCellInst_SboxInst_0_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1725), 
        .B(new_AGEMA_signal_1457), .Z(new_AGEMA_signal_1768) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_0_L0), .B(SubCellInst_SboxInst_0_T3), .Z(
        ShiftRowsOutput[4]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1725), 
        .B(new_AGEMA_signal_1662), .Z(new_AGEMA_signal_1769) );
  XNOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_0_YY_1_), .B(SubCellInst_SboxInst_0_YY_3), .ZN(
        ShiftRowsOutput[5]) );
  XOR2_X1 SubCellInst_SboxInst_0_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1724), .B(new_AGEMA_signal_1768), .Z(new_AGEMA_signal_1826) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U14 ( .A(Fresh[34]), .B(
        SubCellInst_SboxInst_1_Q2), .Z(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U13 ( .A(Fresh[34]), .B(
        new_AGEMA_signal_1600), .Z(SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U10 ( .A1(Ciphertext_s1[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U9 ( .A1(Ciphertext_s0[5]), .A2(
        SubCellInst_SboxInst_1_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND2_U1_U8 ( .A(Fresh[34]), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U7 ( .A1(new_AGEMA_signal_1600), .A2(
        Ciphertext_s1[5]), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q2), 
        .A2(Ciphertext_s0[5]), .ZN(SubCellInst_SboxInst_1_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n8), .B(
        SubCellInst_SboxInst_1_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1665) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_n7), .B(
        SubCellInst_SboxInst_1_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T1) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[5]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[5]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_T1), .B(SubCellInst_SboxInst_1_T2), .Z(
        SubCellInst_SboxInst_1_L0) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1665), 
        .B(new_AGEMA_signal_1552), .Z(new_AGEMA_signal_1727) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U14 ( .A(Fresh[35]), .B(
        SubCellInst_SboxInst_1_Q7), .Z(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U13 ( .A(Fresh[35]), .B(
        new_AGEMA_signal_1601), .Z(SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U10 ( .A1(new_AGEMA_signal_1462), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_1_Q6), 
        .A2(SubCellInst_SboxInst_1_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_1_AND4_U1_U8 ( .A(Fresh[35]), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U7 ( .A1(new_AGEMA_signal_1601), .A2(
        new_AGEMA_signal_1462), .ZN(SubCellInst_SboxInst_1_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_1_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_1_Q7), 
        .A2(SubCellInst_SboxInst_1_Q6), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n8), .B(
        SubCellInst_SboxInst_1_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1666) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_n7), .B(
        SubCellInst_SboxInst_1_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_1_T3) );
  XNOR2_X1 SubCellInst_SboxInst_1_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_1_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_1_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1462), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_1_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_1_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_L2), .Z(
        SubCellInst_SboxInst_1_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1727), 
        .B(new_AGEMA_signal_1463), .Z(new_AGEMA_signal_1770) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_1_L0), .B(SubCellInst_SboxInst_1_T3), .Z(
        ShiftRowsOutput[8]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1727), 
        .B(new_AGEMA_signal_1666), .Z(new_AGEMA_signal_1771) );
  XNOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_1_YY_1_), .B(SubCellInst_SboxInst_1_YY_3), .ZN(
        ShiftRowsOutput[9]) );
  XOR2_X1 SubCellInst_SboxInst_1_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1726), .B(new_AGEMA_signal_1770), .Z(new_AGEMA_signal_1827) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U14 ( .A(Fresh[36]), .B(
        SubCellInst_SboxInst_2_Q2), .Z(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U13 ( .A(Fresh[36]), .B(
        new_AGEMA_signal_1604), .Z(SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U10 ( .A1(Ciphertext_s1[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U9 ( .A1(Ciphertext_s0[9]), .A2(
        SubCellInst_SboxInst_2_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND2_U1_U8 ( .A(Fresh[36]), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U7 ( .A1(new_AGEMA_signal_1604), .A2(
        Ciphertext_s1[9]), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q2), 
        .A2(Ciphertext_s0[9]), .ZN(SubCellInst_SboxInst_2_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n8), .B(
        SubCellInst_SboxInst_2_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1669) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_n7), .B(
        SubCellInst_SboxInst_2_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T1) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[9]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[9]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_T1), .B(SubCellInst_SboxInst_2_T2), .Z(
        SubCellInst_SboxInst_2_L0) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1669), 
        .B(new_AGEMA_signal_1555), .Z(new_AGEMA_signal_1729) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U14 ( .A(Fresh[37]), .B(
        SubCellInst_SboxInst_2_Q7), .Z(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U13 ( .A(Fresh[37]), .B(
        new_AGEMA_signal_1605), .Z(SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U10 ( .A1(new_AGEMA_signal_1468), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_2_Q6), 
        .A2(SubCellInst_SboxInst_2_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_2_AND4_U1_U8 ( .A(Fresh[37]), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U7 ( .A1(new_AGEMA_signal_1605), .A2(
        new_AGEMA_signal_1468), .ZN(SubCellInst_SboxInst_2_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_2_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_2_Q7), 
        .A2(SubCellInst_SboxInst_2_Q6), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n8), .B(
        SubCellInst_SboxInst_2_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1670) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_n7), .B(
        SubCellInst_SboxInst_2_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_2_T3) );
  XNOR2_X1 SubCellInst_SboxInst_2_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_2_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_2_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1468), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_2_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_2_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_L2), .Z(
        SubCellInst_SboxInst_2_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1729), 
        .B(new_AGEMA_signal_1469), .Z(new_AGEMA_signal_1772) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_2_L0), .B(SubCellInst_SboxInst_2_T3), .Z(
        ShiftRowsOutput[12]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1729), 
        .B(new_AGEMA_signal_1670), .Z(new_AGEMA_signal_1773) );
  XNOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_2_YY_1_), .B(SubCellInst_SboxInst_2_YY_3), .ZN(
        ShiftRowsOutput[13]) );
  XOR2_X1 SubCellInst_SboxInst_2_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1728), .B(new_AGEMA_signal_1772), .Z(new_AGEMA_signal_1828) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U14 ( .A(Fresh[38]), .B(
        SubCellInst_SboxInst_3_Q2), .Z(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U13 ( .A(Fresh[38]), .B(
        new_AGEMA_signal_1608), .Z(SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U10 ( .A1(Ciphertext_s1[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U9 ( .A1(Ciphertext_s0[13]), .A2(
        SubCellInst_SboxInst_3_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND2_U1_U8 ( .A(Fresh[38]), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U7 ( .A1(new_AGEMA_signal_1608), .A2(
        Ciphertext_s1[13]), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q2), 
        .A2(Ciphertext_s0[13]), .ZN(SubCellInst_SboxInst_3_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n8), .B(
        SubCellInst_SboxInst_3_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1673) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_n7), .B(
        SubCellInst_SboxInst_3_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T1) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[13]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[13]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_T1), .B(SubCellInst_SboxInst_3_T2), .Z(
        SubCellInst_SboxInst_3_L0) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1673), 
        .B(new_AGEMA_signal_1558), .Z(new_AGEMA_signal_1731) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U14 ( .A(Fresh[39]), .B(
        SubCellInst_SboxInst_3_Q7), .Z(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U13 ( .A(Fresh[39]), .B(
        new_AGEMA_signal_1609), .Z(SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U10 ( .A1(new_AGEMA_signal_1474), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_3_Q6), 
        .A2(SubCellInst_SboxInst_3_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_3_AND4_U1_U8 ( .A(Fresh[39]), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U7 ( .A1(new_AGEMA_signal_1609), .A2(
        new_AGEMA_signal_1474), .ZN(SubCellInst_SboxInst_3_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_3_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_3_Q7), 
        .A2(SubCellInst_SboxInst_3_Q6), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n8), .B(
        SubCellInst_SboxInst_3_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1674) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_n7), .B(
        SubCellInst_SboxInst_3_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_3_T3) );
  XNOR2_X1 SubCellInst_SboxInst_3_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_3_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_3_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1474), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_3_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_3_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_L2), .Z(
        SubCellInst_SboxInst_3_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1731), 
        .B(new_AGEMA_signal_1475), .Z(new_AGEMA_signal_1774) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_3_L0), .B(SubCellInst_SboxInst_3_T3), .Z(
        ShiftRowsOutput[0]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1731), 
        .B(new_AGEMA_signal_1674), .Z(new_AGEMA_signal_1775) );
  XNOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_3_YY_1_), .B(SubCellInst_SboxInst_3_YY_3), .ZN(
        ShiftRowsOutput[1]) );
  XOR2_X1 SubCellInst_SboxInst_3_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1730), .B(new_AGEMA_signal_1774), .Z(new_AGEMA_signal_1829) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U14 ( .A(Fresh[40]), .B(
        SubCellInst_SboxInst_4_Q2), .Z(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U13 ( .A(Fresh[40]), .B(
        new_AGEMA_signal_1612), .Z(SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U10 ( .A1(Ciphertext_s1[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U9 ( .A1(Ciphertext_s0[17]), .A2(
        SubCellInst_SboxInst_4_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND2_U1_U8 ( .A(Fresh[40]), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U7 ( .A1(new_AGEMA_signal_1612), .A2(
        Ciphertext_s1[17]), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q2), 
        .A2(Ciphertext_s0[17]), .ZN(SubCellInst_SboxInst_4_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n8), .B(
        SubCellInst_SboxInst_4_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1677) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_n7), .B(
        SubCellInst_SboxInst_4_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T1) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[17]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[17]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_T1), .B(SubCellInst_SboxInst_4_T2), .Z(
        SubCellInst_SboxInst_4_L0) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1677), 
        .B(new_AGEMA_signal_1561), .Z(new_AGEMA_signal_1733) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U14 ( .A(Fresh[41]), .B(
        SubCellInst_SboxInst_4_Q7), .Z(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U13 ( .A(Fresh[41]), .B(
        new_AGEMA_signal_1613), .Z(SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U10 ( .A1(new_AGEMA_signal_1480), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_4_Q6), 
        .A2(SubCellInst_SboxInst_4_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_4_AND4_U1_U8 ( .A(Fresh[41]), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U7 ( .A1(new_AGEMA_signal_1613), .A2(
        new_AGEMA_signal_1480), .ZN(SubCellInst_SboxInst_4_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_4_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_4_Q7), 
        .A2(SubCellInst_SboxInst_4_Q6), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n8), .B(
        SubCellInst_SboxInst_4_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1678) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_n7), .B(
        SubCellInst_SboxInst_4_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_4_T3) );
  XNOR2_X1 SubCellInst_SboxInst_4_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_4_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_4_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1480), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_4_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_4_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_L2), .Z(
        SubCellInst_SboxInst_4_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1733), 
        .B(new_AGEMA_signal_1481), .Z(new_AGEMA_signal_1776) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_4_L0), .B(SubCellInst_SboxInst_4_T3), .Z(
        ShiftRowsOutput[24]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1733), 
        .B(new_AGEMA_signal_1678), .Z(new_AGEMA_signal_1777) );
  XNOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_4_YY_1_), .B(SubCellInst_SboxInst_4_YY_3), .ZN(
        ShiftRowsOutput[25]) );
  XOR2_X1 SubCellInst_SboxInst_4_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1732), .B(new_AGEMA_signal_1776), .Z(new_AGEMA_signal_1830) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U14 ( .A(Fresh[42]), .B(
        SubCellInst_SboxInst_5_Q2), .Z(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U13 ( .A(Fresh[42]), .B(
        new_AGEMA_signal_1616), .Z(SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U10 ( .A1(Ciphertext_s1[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U9 ( .A1(Ciphertext_s0[21]), .A2(
        SubCellInst_SboxInst_5_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND2_U1_U8 ( .A(Fresh[42]), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U7 ( .A1(new_AGEMA_signal_1616), .A2(
        Ciphertext_s1[21]), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q2), 
        .A2(Ciphertext_s0[21]), .ZN(SubCellInst_SboxInst_5_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n8), .B(
        SubCellInst_SboxInst_5_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1681) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_n7), .B(
        SubCellInst_SboxInst_5_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T1) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[21]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[21]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_T1), .B(SubCellInst_SboxInst_5_T2), .Z(
        SubCellInst_SboxInst_5_L0) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1681), 
        .B(new_AGEMA_signal_1564), .Z(new_AGEMA_signal_1735) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U14 ( .A(Fresh[43]), .B(
        SubCellInst_SboxInst_5_Q7), .Z(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U13 ( .A(Fresh[43]), .B(
        new_AGEMA_signal_1617), .Z(SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U10 ( .A1(new_AGEMA_signal_1486), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_5_Q6), 
        .A2(SubCellInst_SboxInst_5_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_5_AND4_U1_U8 ( .A(Fresh[43]), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U7 ( .A1(new_AGEMA_signal_1617), .A2(
        new_AGEMA_signal_1486), .ZN(SubCellInst_SboxInst_5_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_5_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_5_Q7), 
        .A2(SubCellInst_SboxInst_5_Q6), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n8), .B(
        SubCellInst_SboxInst_5_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1682) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_n7), .B(
        SubCellInst_SboxInst_5_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_5_T3) );
  XNOR2_X1 SubCellInst_SboxInst_5_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_5_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_5_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1486), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_5_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_5_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_L2), .Z(
        SubCellInst_SboxInst_5_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1735), 
        .B(new_AGEMA_signal_1487), .Z(new_AGEMA_signal_1778) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_5_L0), .B(SubCellInst_SboxInst_5_T3), .Z(
        ShiftRowsOutput[28]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1735), 
        .B(new_AGEMA_signal_1682), .Z(new_AGEMA_signal_1779) );
  XNOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_5_YY_1_), .B(SubCellInst_SboxInst_5_YY_3), .ZN(
        ShiftRowsOutput[29]) );
  XOR2_X1 SubCellInst_SboxInst_5_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1734), .B(new_AGEMA_signal_1778), .Z(new_AGEMA_signal_1831) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U14 ( .A(Fresh[44]), .B(
        SubCellInst_SboxInst_6_Q2), .Z(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U13 ( .A(Fresh[44]), .B(
        new_AGEMA_signal_1620), .Z(SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U10 ( .A1(Ciphertext_s1[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U9 ( .A1(Ciphertext_s0[25]), .A2(
        SubCellInst_SboxInst_6_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND2_U1_U8 ( .A(Fresh[44]), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U7 ( .A1(new_AGEMA_signal_1620), .A2(
        Ciphertext_s1[25]), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q2), 
        .A2(Ciphertext_s0[25]), .ZN(SubCellInst_SboxInst_6_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n8), .B(
        SubCellInst_SboxInst_6_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1685) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_n7), .B(
        SubCellInst_SboxInst_6_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T1) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[25]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[25]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_T1), .B(SubCellInst_SboxInst_6_T2), .Z(
        SubCellInst_SboxInst_6_L0) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1685), 
        .B(new_AGEMA_signal_1567), .Z(new_AGEMA_signal_1737) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U14 ( .A(Fresh[45]), .B(
        SubCellInst_SboxInst_6_Q7), .Z(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U13 ( .A(Fresh[45]), .B(
        new_AGEMA_signal_1621), .Z(SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U10 ( .A1(new_AGEMA_signal_1492), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_6_Q6), 
        .A2(SubCellInst_SboxInst_6_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_6_AND4_U1_U8 ( .A(Fresh[45]), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U7 ( .A1(new_AGEMA_signal_1621), .A2(
        new_AGEMA_signal_1492), .ZN(SubCellInst_SboxInst_6_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_6_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_6_Q7), 
        .A2(SubCellInst_SboxInst_6_Q6), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n8), .B(
        SubCellInst_SboxInst_6_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1686) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_n7), .B(
        SubCellInst_SboxInst_6_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_6_T3) );
  XNOR2_X1 SubCellInst_SboxInst_6_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_6_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_6_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1492), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_6_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_6_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_L2), .Z(
        SubCellInst_SboxInst_6_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1737), 
        .B(new_AGEMA_signal_1493), .Z(new_AGEMA_signal_1780) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_6_L0), .B(SubCellInst_SboxInst_6_T3), .Z(
        ShiftRowsOutput[16]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1737), 
        .B(new_AGEMA_signal_1686), .Z(new_AGEMA_signal_1781) );
  XNOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_6_YY_1_), .B(SubCellInst_SboxInst_6_YY_3), .ZN(
        ShiftRowsOutput[17]) );
  XOR2_X1 SubCellInst_SboxInst_6_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1736), .B(new_AGEMA_signal_1780), .Z(new_AGEMA_signal_1832) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U14 ( .A(Fresh[46]), .B(
        SubCellInst_SboxInst_7_Q2), .Z(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U13 ( .A(Fresh[46]), .B(
        new_AGEMA_signal_1624), .Z(SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U10 ( .A1(Ciphertext_s1[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U9 ( .A1(Ciphertext_s0[29]), .A2(
        SubCellInst_SboxInst_7_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND2_U1_U8 ( .A(Fresh[46]), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U7 ( .A1(new_AGEMA_signal_1624), .A2(
        Ciphertext_s1[29]), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q2), 
        .A2(Ciphertext_s0[29]), .ZN(SubCellInst_SboxInst_7_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n8), .B(
        SubCellInst_SboxInst_7_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1689) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_n7), .B(
        SubCellInst_SboxInst_7_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T1) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[29]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[29]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_T1), .B(SubCellInst_SboxInst_7_T2), .Z(
        SubCellInst_SboxInst_7_L0) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1689), 
        .B(new_AGEMA_signal_1570), .Z(new_AGEMA_signal_1739) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U14 ( .A(Fresh[47]), .B(
        SubCellInst_SboxInst_7_Q7), .Z(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U13 ( .A(Fresh[47]), .B(
        new_AGEMA_signal_1625), .Z(SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U10 ( .A1(new_AGEMA_signal_1498), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_7_Q6), 
        .A2(SubCellInst_SboxInst_7_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_7_AND4_U1_U8 ( .A(Fresh[47]), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U7 ( .A1(new_AGEMA_signal_1625), .A2(
        new_AGEMA_signal_1498), .ZN(SubCellInst_SboxInst_7_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_7_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_7_Q7), 
        .A2(SubCellInst_SboxInst_7_Q6), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n8), .B(
        SubCellInst_SboxInst_7_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1690) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_n7), .B(
        SubCellInst_SboxInst_7_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_7_T3) );
  XNOR2_X1 SubCellInst_SboxInst_7_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_7_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_7_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1498), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_7_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_7_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_L2), .Z(
        SubCellInst_SboxInst_7_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1739), 
        .B(new_AGEMA_signal_1499), .Z(new_AGEMA_signal_1782) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_7_L0), .B(SubCellInst_SboxInst_7_T3), .Z(
        ShiftRowsOutput[20]) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1739), 
        .B(new_AGEMA_signal_1690), .Z(new_AGEMA_signal_1783) );
  XNOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_7_YY_1_), .B(SubCellInst_SboxInst_7_YY_3), .ZN(
        SubCellOutput_29) );
  XOR2_X1 SubCellInst_SboxInst_7_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1738), .B(new_AGEMA_signal_1782), .Z(new_AGEMA_signal_1879) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U14 ( .A(Fresh[48]), .B(
        SubCellInst_SboxInst_8_Q2), .Z(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U13 ( .A(Fresh[48]), .B(
        new_AGEMA_signal_1628), .Z(SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U10 ( .A1(Ciphertext_s1[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U9 ( .A1(Ciphertext_s0[33]), .A2(
        SubCellInst_SboxInst_8_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND2_U1_U8 ( .A(Fresh[48]), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U7 ( .A1(new_AGEMA_signal_1628), .A2(
        Ciphertext_s1[33]), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q2), 
        .A2(Ciphertext_s0[33]), .ZN(SubCellInst_SboxInst_8_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n8), .B(
        SubCellInst_SboxInst_8_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1693) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_n7), .B(
        SubCellInst_SboxInst_8_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T1) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[33]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[33]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_T1), .B(SubCellInst_SboxInst_8_T2), .Z(
        SubCellInst_SboxInst_8_L0) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1693), 
        .B(new_AGEMA_signal_1573), .Z(new_AGEMA_signal_1741) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U14 ( .A(Fresh[49]), .B(
        SubCellInst_SboxInst_8_Q7), .Z(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U13 ( .A(Fresh[49]), .B(
        new_AGEMA_signal_1629), .Z(SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U10 ( .A1(new_AGEMA_signal_1504), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_8_Q6), 
        .A2(SubCellInst_SboxInst_8_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_8_AND4_U1_U8 ( .A(Fresh[49]), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U7 ( .A1(new_AGEMA_signal_1629), .A2(
        new_AGEMA_signal_1504), .ZN(SubCellInst_SboxInst_8_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_8_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_8_Q7), 
        .A2(SubCellInst_SboxInst_8_Q6), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n8), .B(
        SubCellInst_SboxInst_8_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1694) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_n7), .B(
        SubCellInst_SboxInst_8_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_8_T3) );
  XNOR2_X1 SubCellInst_SboxInst_8_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_8_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_8_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1504), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_8_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_8_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_L2), .Z(
        SubCellInst_SboxInst_8_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1741), 
        .B(new_AGEMA_signal_1505), .Z(new_AGEMA_signal_1784) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_8_L0), .B(SubCellInst_SboxInst_8_T3), .Z(
        AddRoundConstantOutput[32]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1741), 
        .B(new_AGEMA_signal_1694), .Z(new_AGEMA_signal_1785) );
  XNOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_8_YY_1_), .B(SubCellInst_SboxInst_8_YY_3), .ZN(
        AddRoundConstantOutput[33]) );
  XOR2_X1 SubCellInst_SboxInst_8_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1740), .B(new_AGEMA_signal_1784), .Z(new_AGEMA_signal_1834) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U14 ( .A(Fresh[50]), .B(
        SubCellInst_SboxInst_9_Q2), .Z(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U13 ( .A(Fresh[50]), .B(
        new_AGEMA_signal_1632), .Z(SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U10 ( .A1(Ciphertext_s1[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U9 ( .A1(Ciphertext_s0[37]), .A2(
        SubCellInst_SboxInst_9_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND2_U1_U8 ( .A(Fresh[50]), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U7 ( .A1(new_AGEMA_signal_1632), .A2(
        Ciphertext_s1[37]), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q2), 
        .A2(Ciphertext_s0[37]), .ZN(SubCellInst_SboxInst_9_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n8), .B(
        SubCellInst_SboxInst_9_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1697) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_n7), .B(
        SubCellInst_SboxInst_9_AND2_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T1) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[37]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[37]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_T1), .B(SubCellInst_SboxInst_9_T2), .Z(
        SubCellInst_SboxInst_9_L0) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1697), 
        .B(new_AGEMA_signal_1576), .Z(new_AGEMA_signal_1743) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U14 ( .A(Fresh[51]), .B(
        SubCellInst_SboxInst_9_Q7), .Z(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U13 ( .A(Fresh[51]), .B(
        new_AGEMA_signal_1633), .Z(SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U10 ( .A1(new_AGEMA_signal_1510), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_9_Q6), 
        .A2(SubCellInst_SboxInst_9_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_9_AND4_U1_U8 ( .A(Fresh[51]), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U7 ( .A1(new_AGEMA_signal_1633), .A2(
        new_AGEMA_signal_1510), .ZN(SubCellInst_SboxInst_9_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_9_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_9_Q7), 
        .A2(SubCellInst_SboxInst_9_Q6), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n8), .B(
        SubCellInst_SboxInst_9_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1698) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_n7), .B(
        SubCellInst_SboxInst_9_AND4_U1_z_0__0_), .ZN(SubCellInst_SboxInst_9_T3) );
  XNOR2_X1 SubCellInst_SboxInst_9_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_9_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_9_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1510), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_9_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_9_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_L2), .Z(
        SubCellInst_SboxInst_9_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1743), 
        .B(new_AGEMA_signal_1511), .Z(new_AGEMA_signal_1786) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_9_L0), .B(SubCellInst_SboxInst_9_T3), .Z(
        AddRoundConstantOutput[36]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1743), 
        .B(new_AGEMA_signal_1698), .Z(new_AGEMA_signal_1787) );
  XNOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_9_YY_1_), .B(SubCellInst_SboxInst_9_YY_3), .ZN(
        AddRoundConstantOutput[37]) );
  XOR2_X1 SubCellInst_SboxInst_9_XOR_o1_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1742), .B(new_AGEMA_signal_1786), .Z(new_AGEMA_signal_1835) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U14 ( .A(Fresh[52]), .B(
        SubCellInst_SboxInst_10_Q2), .Z(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U13 ( .A(Fresh[52]), .B(
        new_AGEMA_signal_1636), .Z(SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U10 ( .A1(Ciphertext_s1[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U9 ( .A1(Ciphertext_s0[41]), .A2(
        SubCellInst_SboxInst_10_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND2_U1_U8 ( .A(Fresh[52]), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U7 ( .A1(new_AGEMA_signal_1636), 
        .A2(Ciphertext_s1[41]), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q2), 
        .A2(Ciphertext_s0[41]), .ZN(SubCellInst_SboxInst_10_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n8), .B(
        SubCellInst_SboxInst_10_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1701)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_n7), .B(
        SubCellInst_SboxInst_10_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T1) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[41]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[41]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_T1), .B(SubCellInst_SboxInst_10_T2), .Z(
        SubCellInst_SboxInst_10_L0) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1701), 
        .B(new_AGEMA_signal_1579), .Z(new_AGEMA_signal_1745) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U14 ( .A(Fresh[53]), .B(
        SubCellInst_SboxInst_10_Q7), .Z(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U13 ( .A(Fresh[53]), .B(
        new_AGEMA_signal_1637), .Z(SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U10 ( .A1(new_AGEMA_signal_1516), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_10_Q6), 
        .A2(SubCellInst_SboxInst_10_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_10_AND4_U1_U8 ( .A(Fresh[53]), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U7 ( .A1(new_AGEMA_signal_1637), 
        .A2(new_AGEMA_signal_1516), .ZN(SubCellInst_SboxInst_10_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_10_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_10_Q7), 
        .A2(SubCellInst_SboxInst_10_Q6), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n8), .B(
        SubCellInst_SboxInst_10_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1702)
         );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_n7), .B(
        SubCellInst_SboxInst_10_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_10_T3) );
  XNOR2_X1 SubCellInst_SboxInst_10_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_10_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1516), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_10_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_10_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_10_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_L2), .Z(
        SubCellInst_SboxInst_10_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1745), 
        .B(new_AGEMA_signal_1517), .Z(new_AGEMA_signal_1788) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_10_L0), .B(SubCellInst_SboxInst_10_T3), .Z(
        AddRoundConstantOutput[40]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1745), .B(new_AGEMA_signal_1702), .Z(new_AGEMA_signal_1789) );
  XNOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_10_YY_1_), .B(SubCellInst_SboxInst_10_YY_3), .ZN(
        AddRoundConstantOutput[41]) );
  XOR2_X1 SubCellInst_SboxInst_10_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1744), .B(new_AGEMA_signal_1788), .Z(
        new_AGEMA_signal_1836) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U14 ( .A(Fresh[54]), .B(
        SubCellInst_SboxInst_11_Q2), .Z(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U13 ( .A(Fresh[54]), .B(
        new_AGEMA_signal_1640), .Z(SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U10 ( .A1(Ciphertext_s1[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U9 ( .A1(Ciphertext_s0[45]), .A2(
        SubCellInst_SboxInst_11_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND2_U1_U8 ( .A(Fresh[54]), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U7 ( .A1(new_AGEMA_signal_1640), 
        .A2(Ciphertext_s1[45]), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q2), 
        .A2(Ciphertext_s0[45]), .ZN(SubCellInst_SboxInst_11_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n8), .B(
        SubCellInst_SboxInst_11_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1705)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_n7), .B(
        SubCellInst_SboxInst_11_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T1) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[45]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[45]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_T1), .B(SubCellInst_SboxInst_11_T2), .Z(
        SubCellInst_SboxInst_11_L0) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1705), 
        .B(new_AGEMA_signal_1582), .Z(new_AGEMA_signal_1747) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U14 ( .A(Fresh[55]), .B(
        SubCellInst_SboxInst_11_Q7), .Z(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U13 ( .A(Fresh[55]), .B(
        new_AGEMA_signal_1641), .Z(SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U10 ( .A1(new_AGEMA_signal_1522), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_11_Q6), 
        .A2(SubCellInst_SboxInst_11_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_11_AND4_U1_U8 ( .A(Fresh[55]), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U7 ( .A1(new_AGEMA_signal_1641), 
        .A2(new_AGEMA_signal_1522), .ZN(SubCellInst_SboxInst_11_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_11_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_11_Q7), 
        .A2(SubCellInst_SboxInst_11_Q6), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n8), .B(
        SubCellInst_SboxInst_11_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1706)
         );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_n7), .B(
        SubCellInst_SboxInst_11_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_11_T3) );
  XNOR2_X1 SubCellInst_SboxInst_11_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_11_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1522), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_11_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_11_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_11_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_L2), .Z(
        SubCellInst_SboxInst_11_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1747), 
        .B(new_AGEMA_signal_1523), .Z(new_AGEMA_signal_1790) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_11_L0), .B(SubCellInst_SboxInst_11_T3), .Z(
        SubCellOutput_44) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1747), .B(new_AGEMA_signal_1706), .Z(new_AGEMA_signal_1791) );
  XNOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_11_YY_1_), .B(SubCellInst_SboxInst_11_YY_3), .ZN(
        SubCellOutput_45) );
  XOR2_X1 SubCellInst_SboxInst_11_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1746), .B(new_AGEMA_signal_1790), .Z(
        new_AGEMA_signal_1837) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U14 ( .A(Fresh[56]), .B(
        SubCellInst_SboxInst_12_Q2), .Z(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U13 ( .A(Fresh[56]), .B(
        new_AGEMA_signal_1644), .Z(SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U10 ( .A1(Ciphertext_s1[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U9 ( .A1(Ciphertext_s0[49]), .A2(
        SubCellInst_SboxInst_12_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND2_U1_U8 ( .A(Fresh[56]), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U7 ( .A1(new_AGEMA_signal_1644), 
        .A2(Ciphertext_s1[49]), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q2), 
        .A2(Ciphertext_s0[49]), .ZN(SubCellInst_SboxInst_12_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n8), .B(
        SubCellInst_SboxInst_12_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1709)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_n7), .B(
        SubCellInst_SboxInst_12_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T1) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[49]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[49]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_T1), .B(SubCellInst_SboxInst_12_T2), .Z(
        SubCellInst_SboxInst_12_L0) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1709), 
        .B(new_AGEMA_signal_1585), .Z(new_AGEMA_signal_1749) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U14 ( .A(Fresh[57]), .B(
        SubCellInst_SboxInst_12_Q7), .Z(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U13 ( .A(Fresh[57]), .B(
        new_AGEMA_signal_1645), .Z(SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U10 ( .A1(new_AGEMA_signal_1528), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_12_Q6), 
        .A2(SubCellInst_SboxInst_12_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_12_AND4_U1_U8 ( .A(Fresh[57]), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U7 ( .A1(new_AGEMA_signal_1645), 
        .A2(new_AGEMA_signal_1528), .ZN(SubCellInst_SboxInst_12_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_12_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_12_Q7), 
        .A2(SubCellInst_SboxInst_12_Q6), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n8), .B(
        SubCellInst_SboxInst_12_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1710)
         );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_n7), .B(
        SubCellInst_SboxInst_12_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_12_T3) );
  XNOR2_X1 SubCellInst_SboxInst_12_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_12_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1528), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_12_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_12_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_12_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_L2), .Z(
        SubCellInst_SboxInst_12_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1749), 
        .B(new_AGEMA_signal_1529), .Z(new_AGEMA_signal_1792) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_12_L0), .B(SubCellInst_SboxInst_12_T3), .Z(
        AddRoundConstantOutput[48]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1749), .B(new_AGEMA_signal_1710), .Z(new_AGEMA_signal_1793) );
  XNOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_12_YY_1_), .B(SubCellInst_SboxInst_12_YY_3), .ZN(
        AddRoundConstantOutput[49]) );
  XOR2_X1 SubCellInst_SboxInst_12_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1748), .B(new_AGEMA_signal_1792), .Z(
        new_AGEMA_signal_1838) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U14 ( .A(Fresh[58]), .B(
        SubCellInst_SboxInst_13_Q2), .Z(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U13 ( .A(Fresh[58]), .B(
        new_AGEMA_signal_1648), .Z(SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U10 ( .A1(Ciphertext_s1[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U9 ( .A1(Ciphertext_s0[53]), .A2(
        SubCellInst_SboxInst_13_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND2_U1_U8 ( .A(Fresh[58]), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U7 ( .A1(new_AGEMA_signal_1648), 
        .A2(Ciphertext_s1[53]), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q2), 
        .A2(Ciphertext_s0[53]), .ZN(SubCellInst_SboxInst_13_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n8), .B(
        SubCellInst_SboxInst_13_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1713)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_n7), .B(
        SubCellInst_SboxInst_13_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T1) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[53]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[53]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_T1), .B(SubCellInst_SboxInst_13_T2), .Z(
        SubCellInst_SboxInst_13_L0) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1713), 
        .B(new_AGEMA_signal_1588), .Z(new_AGEMA_signal_1751) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U14 ( .A(Fresh[59]), .B(
        SubCellInst_SboxInst_13_Q7), .Z(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U13 ( .A(Fresh[59]), .B(
        new_AGEMA_signal_1649), .Z(SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U10 ( .A1(new_AGEMA_signal_1534), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_13_Q6), 
        .A2(SubCellInst_SboxInst_13_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_13_AND4_U1_U8 ( .A(Fresh[59]), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U7 ( .A1(new_AGEMA_signal_1649), 
        .A2(new_AGEMA_signal_1534), .ZN(SubCellInst_SboxInst_13_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_13_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_13_Q7), 
        .A2(SubCellInst_SboxInst_13_Q6), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n8), .B(
        SubCellInst_SboxInst_13_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1714)
         );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_n7), .B(
        SubCellInst_SboxInst_13_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_13_T3) );
  XNOR2_X1 SubCellInst_SboxInst_13_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_13_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1534), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_13_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_13_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_13_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_L2), .Z(
        SubCellInst_SboxInst_13_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1751), 
        .B(new_AGEMA_signal_1535), .Z(new_AGEMA_signal_1794) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_13_L0), .B(SubCellInst_SboxInst_13_T3), .Z(
        AddRoundConstantOutput[52]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1751), .B(new_AGEMA_signal_1714), .Z(new_AGEMA_signal_1795) );
  XNOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_13_YY_1_), .B(SubCellInst_SboxInst_13_YY_3), .ZN(
        AddRoundConstantOutput[53]) );
  XOR2_X1 SubCellInst_SboxInst_13_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1750), .B(new_AGEMA_signal_1794), .Z(
        new_AGEMA_signal_1839) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U14 ( .A(Fresh[60]), .B(
        SubCellInst_SboxInst_14_Q2), .Z(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U13 ( .A(Fresh[60]), .B(
        new_AGEMA_signal_1652), .Z(SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U10 ( .A1(Ciphertext_s1[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U9 ( .A1(Ciphertext_s0[57]), .A2(
        SubCellInst_SboxInst_14_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND2_U1_U8 ( .A(Fresh[60]), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U7 ( .A1(new_AGEMA_signal_1652), 
        .A2(Ciphertext_s1[57]), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q2), 
        .A2(Ciphertext_s0[57]), .ZN(SubCellInst_SboxInst_14_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n8), .B(
        SubCellInst_SboxInst_14_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1717)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_n7), .B(
        SubCellInst_SboxInst_14_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T1) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[57]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[57]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_T1), .B(SubCellInst_SboxInst_14_T2), .Z(
        SubCellInst_SboxInst_14_L0) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1717), 
        .B(new_AGEMA_signal_1591), .Z(new_AGEMA_signal_1753) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U14 ( .A(Fresh[61]), .B(
        SubCellInst_SboxInst_14_Q7), .Z(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U13 ( .A(Fresh[61]), .B(
        new_AGEMA_signal_1653), .Z(SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U10 ( .A1(new_AGEMA_signal_1540), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_14_Q6), 
        .A2(SubCellInst_SboxInst_14_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_14_AND4_U1_U8 ( .A(Fresh[61]), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U7 ( .A1(new_AGEMA_signal_1653), 
        .A2(new_AGEMA_signal_1540), .ZN(SubCellInst_SboxInst_14_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_14_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_14_Q7), 
        .A2(SubCellInst_SboxInst_14_Q6), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n8), .B(
        SubCellInst_SboxInst_14_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1718)
         );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_n7), .B(
        SubCellInst_SboxInst_14_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_14_T3) );
  XNOR2_X1 SubCellInst_SboxInst_14_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_14_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1540), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_14_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_14_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_14_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_L2), .Z(
        SubCellInst_SboxInst_14_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1753), 
        .B(new_AGEMA_signal_1541), .Z(new_AGEMA_signal_1796) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_14_L0), .B(SubCellInst_SboxInst_14_T3), .Z(
        AddRoundConstantOutput[56]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1753), .B(new_AGEMA_signal_1718), .Z(new_AGEMA_signal_1797) );
  XNOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_14_YY_1_), .B(SubCellInst_SboxInst_14_YY_3), .ZN(
        AddRoundConstantOutput[57]) );
  XOR2_X1 SubCellInst_SboxInst_14_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1752), .B(new_AGEMA_signal_1796), .Z(
        new_AGEMA_signal_1840) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U14 ( .A(Fresh[62]), .B(
        SubCellInst_SboxInst_15_Q2), .Z(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U13 ( .A(Fresh[62]), .B(
        new_AGEMA_signal_1656), .Z(SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U10 ( .A1(Ciphertext_s1[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U9 ( .A1(Ciphertext_s0[61]), .A2(
        SubCellInst_SboxInst_15_AND2_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND2_U1_U8 ( .A(Fresh[62]), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U7 ( .A1(new_AGEMA_signal_1656), 
        .A2(Ciphertext_s1[61]), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND2_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q2), 
        .A2(Ciphertext_s0[61]), .ZN(SubCellInst_SboxInst_15_AND2_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n8), .B(
        SubCellInst_SboxInst_15_AND2_U1_z_1__1_), .ZN(new_AGEMA_signal_1721)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_n7), .B(
        SubCellInst_SboxInst_15_AND2_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T1) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND2_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND2_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_0_s_current_state_reg ( .D(
        Ciphertext_s0[61]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_a_i_1_s_current_state_reg ( .D(
        Ciphertext_s1[61]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND2_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND2_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND2_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_T1), .B(SubCellInst_SboxInst_15_T2), .Z(
        SubCellInst_SboxInst_15_L0) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR4_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1721), 
        .B(new_AGEMA_signal_1594), .Z(new_AGEMA_signal_1755) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U14 ( .A(Fresh[63]), .B(
        SubCellInst_SboxInst_15_Q7), .Z(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_) );
  XOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U13 ( .A(Fresh[63]), .B(
        new_AGEMA_signal_1657), .Z(SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_)
         );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U12 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[1]), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U11 ( .A1(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[0]), .A2(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U10 ( .A1(new_AGEMA_signal_1546), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_) );
  NOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U9 ( .A1(SubCellInst_SboxInst_15_Q6), 
        .A2(SubCellInst_SboxInst_15_AND4_U1_n9), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_) );
  INV_X1 SubCellInst_SboxInst_15_AND4_U1_U8 ( .A(Fresh[63]), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n9) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U7 ( .A1(new_AGEMA_signal_1657), 
        .A2(new_AGEMA_signal_1546), .ZN(SubCellInst_SboxInst_15_AND4_U1_mul[1]) );
  AND2_X1 SubCellInst_SboxInst_15_AND4_U1_U6 ( .A1(SubCellInst_SboxInst_15_Q7), 
        .A2(SubCellInst_SboxInst_15_Q6), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_mul[0]) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U5 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n8), .B(
        SubCellInst_SboxInst_15_AND4_U1_z_1__1_), .ZN(new_AGEMA_signal_1722)
         );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U4 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n8) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U3 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_n7), .B(
        SubCellInst_SboxInst_15_AND4_U1_z_0__0_), .ZN(
        SubCellInst_SboxInst_15_T3) );
  XNOR2_X1 SubCellInst_SboxInst_15_AND4_U1_U2 ( .A(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .B(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .ZN(
        SubCellInst_SboxInst_15_AND4_U1_n7) );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[0]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z_0__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_Q6), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[0]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_0_1_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_0_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_0__1_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s1_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_mul_pipe_s2_1_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_mul_s1_out[1]), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_z_1__1_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_a_i_1_s_current_state_reg ( .D(
        new_AGEMA_signal_1546), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_a_reg[1]), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_s_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_s_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_s_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_0_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_1_reg_1_0_s_current_state_reg ( .D(
        SubCellInst_SboxInst_15_AND4_U1_p_1_in_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_1_out_1__0_), .QN() );
  DFF_X1 SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_1_0_s_current_state_reg ( 
        .D(SubCellInst_SboxInst_15_AND4_U1_p_0_out_1__0_), .CK(clk), .Q(
        SubCellInst_SboxInst_15_AND4_U1_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_L2), .Z(
        SubCellInst_SboxInst_15_YY_3) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR9_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1755), 
        .B(new_AGEMA_signal_1547), .Z(new_AGEMA_signal_1798) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_0_U1 ( .A(
        SubCellInst_SboxInst_15_L0), .B(SubCellInst_SboxInst_15_T3), .Z(
        SubCellOutput[60]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR10_U1_Ins_1_U1 ( .A(new_AGEMA_signal_1755), .B(new_AGEMA_signal_1722), .Z(new_AGEMA_signal_1799) );
  XNOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins0_U1 ( .A(
        SubCellInst_SboxInst_15_YY_1_), .B(SubCellInst_SboxInst_15_YY_3), .ZN(
        SubCellOutput[61]) );
  XOR2_X1 SubCellInst_SboxInst_15_XOR_o1_U1_Ins_1_U1 ( .A(
        new_AGEMA_signal_1754), .B(new_AGEMA_signal_1798), .Z(
        new_AGEMA_signal_1841) );
  INV_X1 AddConstXOR_U2_U1 ( .A(SubCellOutput_29), .ZN(ShiftRowsOutput[21]) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_0_n1), .B(FSMUpdate[1]), .ZN(
        AddRoundConstantOutput[60]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1842), .B(1'b0), .Z(new_AGEMA_signal_1880) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[60]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1799), .Z(new_AGEMA_signal_1842) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_0_1_n1), .B(FSM_1), .ZN(
        AddRoundConstantOutput[61]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1881), .B(1'b0), .Z(new_AGEMA_signal_1947) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput[61]), .ZN(AddConstXOR_AddConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1841), .Z(new_AGEMA_signal_1881) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_0_n1), .B(FSM[4]), .ZN(
        AddRoundConstantOutput[44]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1844), .B(1'b0), .Z(new_AGEMA_signal_1882) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_44), .ZN(AddConstXOR_AddConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1791), .Z(new_AGEMA_signal_1844) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddConstXOR_AddConstXOR_XORInst_1_1_n1), .B(FSM[5]), .ZN(
        AddRoundConstantOutput[45]) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1883), .B(1'b0), .Z(new_AGEMA_signal_1948) );
  XNOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        SubCellOutput_45), .ZN(AddConstXOR_AddConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddConstXOR_AddConstXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1837), .Z(new_AGEMA_signal_1883) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_0_n1), .B(
        TweakeyGeneration_key_Feedback[0]), .ZN(ShiftRowsOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1846), .B(new_AGEMA_signal_1260), .Z(
        new_AGEMA_signal_1884) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[32]), .ZN(AddRoundTweakeyXOR_XORInst_0_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1785), .Z(new_AGEMA_signal_1846) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_0_1_n1), .B(
        TweakeyGeneration_key_Feedback[1]), .ZN(ShiftRowsOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1885), .B(new_AGEMA_signal_1263), .Z(
        new_AGEMA_signal_1949) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[33]), .ZN(AddRoundTweakeyXOR_XORInst_0_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1834), .Z(new_AGEMA_signal_1885) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_0_n1), .B(
        TweakeyGeneration_key_Feedback[4]), .ZN(ShiftRowsOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1848), .B(new_AGEMA_signal_1272), .Z(
        new_AGEMA_signal_1886) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[36]), .ZN(AddRoundTweakeyXOR_XORInst_1_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1787), .Z(new_AGEMA_signal_1848) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_1_1_n1), .B(
        TweakeyGeneration_key_Feedback[5]), .ZN(ShiftRowsOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1887), .B(new_AGEMA_signal_1275), .Z(
        new_AGEMA_signal_1950) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[37]), .ZN(AddRoundTweakeyXOR_XORInst_1_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1835), .Z(new_AGEMA_signal_1887) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_0_n1), .B(
        TweakeyGeneration_key_Feedback[8]), .ZN(ShiftRowsOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1850), .B(new_AGEMA_signal_1284), .Z(
        new_AGEMA_signal_1888) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[40]), .ZN(AddRoundTweakeyXOR_XORInst_2_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1789), .Z(new_AGEMA_signal_1850) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_2_1_n1), .B(
        TweakeyGeneration_key_Feedback[9]), .ZN(ShiftRowsOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1889), .B(new_AGEMA_signal_1287), .Z(
        new_AGEMA_signal_1951) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[41]), .ZN(AddRoundTweakeyXOR_XORInst_2_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1836), .Z(new_AGEMA_signal_1889) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_0_n1), .B(
        TweakeyGeneration_key_Feedback[12]), .ZN(ShiftRowsOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1952), .B(new_AGEMA_signal_1296), .Z(
        new_AGEMA_signal_2007) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[44]), .ZN(AddRoundTweakeyXOR_XORInst_3_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1882), .Z(new_AGEMA_signal_1952) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_3_1_n1), .B(
        TweakeyGeneration_key_Feedback[13]), .ZN(ShiftRowsOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2008), .B(new_AGEMA_signal_1299), .Z(
        new_AGEMA_signal_2061) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[45]), .ZN(AddRoundTweakeyXOR_XORInst_3_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1948), .Z(new_AGEMA_signal_2008) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_0_n1), .B(
        TweakeyGeneration_key_Feedback[16]), .ZN(MCOutput[32]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1853), .B(new_AGEMA_signal_1308), .Z(
        new_AGEMA_signal_1892) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[48]), .ZN(AddRoundTweakeyXOR_XORInst_4_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1793), .Z(new_AGEMA_signal_1853) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_4_1_n1), .B(
        TweakeyGeneration_key_Feedback[17]), .ZN(MCOutput[33]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1893), .B(new_AGEMA_signal_1311), .Z(
        new_AGEMA_signal_1954) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[49]), .ZN(AddRoundTweakeyXOR_XORInst_4_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_4_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1838), .Z(new_AGEMA_signal_1893) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_0_n1), .B(
        TweakeyGeneration_key_Feedback[20]), .ZN(MCOutput[36]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1855), .B(new_AGEMA_signal_1320), .Z(
        new_AGEMA_signal_1894) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[52]), .ZN(AddRoundTweakeyXOR_XORInst_5_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1795), .Z(new_AGEMA_signal_1855) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_5_1_n1), .B(
        TweakeyGeneration_key_Feedback[21]), .ZN(MCOutput[37]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1895), .B(new_AGEMA_signal_1323), .Z(
        new_AGEMA_signal_1955) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[53]), .ZN(AddRoundTweakeyXOR_XORInst_5_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_5_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1839), .Z(new_AGEMA_signal_1895) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_0_n1), .B(
        TweakeyGeneration_key_Feedback[24]), .ZN(MCOutput[40]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1857), .B(new_AGEMA_signal_1332), .Z(
        new_AGEMA_signal_1896) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[56]), .ZN(AddRoundTweakeyXOR_XORInst_6_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1797), .Z(new_AGEMA_signal_1857) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_6_1_n1), .B(
        TweakeyGeneration_key_Feedback[25]), .ZN(MCOutput[41]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1897), .B(new_AGEMA_signal_1335), .Z(
        new_AGEMA_signal_1956) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[57]), .ZN(AddRoundTweakeyXOR_XORInst_6_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_6_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1840), .Z(new_AGEMA_signal_1897) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_0_n1), .B(
        TweakeyGeneration_key_Feedback[28]), .ZN(MCOutput[44]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_1957), .B(new_AGEMA_signal_1344), .Z(
        new_AGEMA_signal_2009) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[60]), .ZN(AddRoundTweakeyXOR_XORInst_7_0_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1880), .Z(new_AGEMA_signal_1957) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins0_U1 ( .A(
        AddRoundTweakeyXOR_XORInst_7_1_n1), .B(
        TweakeyGeneration_key_Feedback[29]), .ZN(MCOutput[45]) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U2_Ins_1_U1 ( .A(
        new_AGEMA_signal_2010), .B(new_AGEMA_signal_1347), .Z(
        new_AGEMA_signal_2062) );
  XNOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins0_U1 ( .A(1'b0), .B(
        AddRoundConstantOutput[61]), .ZN(AddRoundTweakeyXOR_XORInst_7_1_n1) );
  XOR2_X1 AddRoundTweakeyXOR_XORInst_7_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1947), .Z(new_AGEMA_signal_2010) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_0_n2), 
        .B(MCInst_MCR0_XORInst_0_0_n1), .ZN(MCOutput[48]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1959), .B(
        new_AGEMA_signal_1860), .Z(new_AGEMA_signal_2011) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[16]), .B(
        ShiftRowsOutput[0]), .ZN(MCInst_MCR0_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1781), .B(
        new_AGEMA_signal_1775), .Z(new_AGEMA_signal_1860) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .Z(MCInst_MCR0_XORInst_0_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1892), .Z(new_AGEMA_signal_1959) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_0_1_n2), 
        .B(MCInst_MCR0_XORInst_0_1_n1), .ZN(MCOutput[49]) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2012), .B(
        new_AGEMA_signal_1900), .Z(new_AGEMA_signal_2063) );
  XNOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[17]), .B(
        ShiftRowsOutput[1]), .ZN(MCInst_MCR0_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1832), .B(
        new_AGEMA_signal_1829), .Z(new_AGEMA_signal_1900) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .Z(MCInst_MCR0_XORInst_0_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1954), .Z(new_AGEMA_signal_2012) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_0_n2), 
        .B(MCInst_MCR0_XORInst_1_0_n1), .ZN(MCOutput[52]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1961), .B(
        new_AGEMA_signal_1862), .Z(new_AGEMA_signal_2013) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[20]), .B(
        ShiftRowsOutput[4]), .ZN(MCInst_MCR0_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1783), .B(
        new_AGEMA_signal_1769), .Z(new_AGEMA_signal_1862) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .Z(MCInst_MCR0_XORInst_1_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1894), .Z(new_AGEMA_signal_1961) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_1_1_n2), 
        .B(MCInst_MCR0_XORInst_1_1_n1), .ZN(MCOutput[53]) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2014), .B(
        new_AGEMA_signal_1962), .Z(new_AGEMA_signal_2064) );
  XNOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[21]), .B(
        ShiftRowsOutput[5]), .ZN(MCInst_MCR0_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1879), .B(
        new_AGEMA_signal_1826), .Z(new_AGEMA_signal_1962) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .Z(MCInst_MCR0_XORInst_1_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1955), .Z(new_AGEMA_signal_2014) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_0_n2), 
        .B(MCInst_MCR0_XORInst_2_0_n1), .ZN(MCOutput[56]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_1964), .B(
        new_AGEMA_signal_1864), .Z(new_AGEMA_signal_2015) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[24]), .B(
        ShiftRowsOutput[8]), .ZN(MCInst_MCR0_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1777), .B(
        new_AGEMA_signal_1771), .Z(new_AGEMA_signal_1864) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .Z(MCInst_MCR0_XORInst_2_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1896), .Z(new_AGEMA_signal_1964) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_2_1_n2), 
        .B(MCInst_MCR0_XORInst_2_1_n1), .ZN(MCOutput[57]) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2016), .B(
        new_AGEMA_signal_1905), .Z(new_AGEMA_signal_2065) );
  XNOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[25]), .B(
        ShiftRowsOutput[9]), .ZN(MCInst_MCR0_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1830), .B(
        new_AGEMA_signal_1827), .Z(new_AGEMA_signal_1905) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .Z(MCInst_MCR0_XORInst_2_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2016) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_0_n2), 
        .B(MCInst_MCR0_XORInst_3_0_n1), .ZN(MCOutput[60]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2066), .B(
        new_AGEMA_signal_1866), .Z(new_AGEMA_signal_2104) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins0_U1 ( .A(ShiftRowsOutput[28]), .B(
        ShiftRowsOutput[12]), .ZN(MCInst_MCR0_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1779), .B(
        new_AGEMA_signal_1773), .Z(new_AGEMA_signal_1866) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .Z(MCInst_MCR0_XORInst_3_0_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2009), .Z(new_AGEMA_signal_2066) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins0_U1 ( .A(MCInst_MCR0_XORInst_3_1_n2), 
        .B(MCInst_MCR0_XORInst_3_1_n1), .ZN(MCOutput[61]) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U3_Ins_1_U1 ( .A(new_AGEMA_signal_2105), .B(
        new_AGEMA_signal_1908), .Z(new_AGEMA_signal_2116) );
  XNOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins0_U1 ( .A(ShiftRowsOutput[29]), .B(
        ShiftRowsOutput[13]), .ZN(MCInst_MCR0_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1831), .B(
        new_AGEMA_signal_1828), .Z(new_AGEMA_signal_1908) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .Z(MCInst_MCR0_XORInst_3_1_n2) );
  XOR2_X1 MCInst_MCR0_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2062), .Z(new_AGEMA_signal_2105) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[16]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1967), .B(
        new_AGEMA_signal_1781), .Z(new_AGEMA_signal_2019) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[32]), .ZN(MCInst_MCR2_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1886), .Z(new_AGEMA_signal_1967) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[17]) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2020), .B(
        new_AGEMA_signal_1832), .Z(new_AGEMA_signal_2068) );
  XNOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[33]), .ZN(MCInst_MCR2_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1950), .Z(new_AGEMA_signal_2020) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[20]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1969), .B(
        new_AGEMA_signal_1783), .Z(new_AGEMA_signal_2021) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[36]), .ZN(MCInst_MCR2_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1888), .Z(new_AGEMA_signal_1969) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[21]) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2022), .B(
        new_AGEMA_signal_1879), .Z(new_AGEMA_signal_2069) );
  XNOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[37]), .ZN(MCInst_MCR2_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1951), .Z(new_AGEMA_signal_2022) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[24]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2070), .B(
        new_AGEMA_signal_1777), .Z(new_AGEMA_signal_2106) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[40]), .ZN(MCInst_MCR2_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2007), .Z(new_AGEMA_signal_2070) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[25]) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2107), .B(
        new_AGEMA_signal_1830), .Z(new_AGEMA_signal_2117) );
  XNOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[41]), .ZN(MCInst_MCR2_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2061), .Z(new_AGEMA_signal_2107) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[28]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1972), .B(
        new_AGEMA_signal_1779), .Z(new_AGEMA_signal_2025) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[44]), .ZN(MCInst_MCR2_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1884), .Z(new_AGEMA_signal_1972) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR2_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[29]) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2026), .B(
        new_AGEMA_signal_1831), .Z(new_AGEMA_signal_2072) );
  XNOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(
        ShiftRowsOutput[45]), .ZN(MCInst_MCR2_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR2_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1949), .Z(new_AGEMA_signal_2026) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_0_n1), 
        .B(ShiftRowsOutput[16]), .ZN(MCOutput[0]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1974), .B(
        new_AGEMA_signal_1781), .Z(new_AGEMA_signal_2027) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[32]), 
        .ZN(MCInst_MCR3_XORInst_0_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1892), .Z(new_AGEMA_signal_1974) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_0_1_n1), 
        .B(ShiftRowsOutput[17]), .ZN(MCOutput[1]) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2028), .B(
        new_AGEMA_signal_1832), .Z(new_AGEMA_signal_2073) );
  XNOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[33]), 
        .ZN(MCInst_MCR3_XORInst_0_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_0_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1954), .Z(new_AGEMA_signal_2028) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_0_n1), 
        .B(ShiftRowsOutput[20]), .ZN(MCOutput[4]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1976), .B(
        new_AGEMA_signal_1783), .Z(new_AGEMA_signal_2029) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[36]), 
        .ZN(MCInst_MCR3_XORInst_1_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1894), .Z(new_AGEMA_signal_1976) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_1_1_n1), 
        .B(ShiftRowsOutput[21]), .ZN(MCOutput[5]) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2030), .B(
        new_AGEMA_signal_1879), .Z(new_AGEMA_signal_2074) );
  XNOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[37]), 
        .ZN(MCInst_MCR3_XORInst_1_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_1_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1955), .Z(new_AGEMA_signal_2030) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_0_n1), 
        .B(ShiftRowsOutput[24]), .ZN(MCOutput[8]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_1978), .B(
        new_AGEMA_signal_1777), .Z(new_AGEMA_signal_2031) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[40]), 
        .ZN(MCInst_MCR3_XORInst_2_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1896), .Z(new_AGEMA_signal_1978) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_2_1_n1), 
        .B(ShiftRowsOutput[25]), .ZN(MCOutput[9]) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2032), .B(
        new_AGEMA_signal_1830), .Z(new_AGEMA_signal_2075) );
  XNOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[41]), 
        .ZN(MCInst_MCR3_XORInst_2_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_2_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_1956), .Z(new_AGEMA_signal_2032) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_0_n1), 
        .B(ShiftRowsOutput[28]), .ZN(MCOutput[12]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2076), .B(
        new_AGEMA_signal_1779), .Z(new_AGEMA_signal_2108) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[44]), 
        .ZN(MCInst_MCR3_XORInst_3_0_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_0_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2009), .Z(new_AGEMA_signal_2076) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins0_U1 ( .A(MCInst_MCR3_XORInst_3_1_n1), 
        .B(ShiftRowsOutput[29]), .ZN(MCOutput[13]) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U2_Ins_1_U1 ( .A(new_AGEMA_signal_2109), .B(
        new_AGEMA_signal_1831), .Z(new_AGEMA_signal_2118) );
  XNOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins0_U1 ( .A(1'b0), .B(MCOutput[45]), 
        .ZN(MCInst_MCR3_XORInst_3_1_n1) );
  XOR2_X1 MCInst_MCR3_XORInst_3_1_U1_Ins_1_U1 ( .A(1'b0), .B(
        new_AGEMA_signal_2062), .Z(new_AGEMA_signal_2109) );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[63]), .CK(clk_gated), .Q(Ciphertext_s0[63]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2103), .CK(clk_gated), .Q(Ciphertext_s1[63]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[62]), .CK(clk_gated), .Q(Ciphertext_s0[62]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2060), .CK(clk_gated), .Q(Ciphertext_s1[62]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[61]), .CK(clk_gated), .Q(Ciphertext_s0[61]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2124), .CK(clk_gated), .Q(Ciphertext_s1[61]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[60]), .CK(clk_gated), .Q(Ciphertext_s0[60]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2115), .CK(clk_gated), .Q(Ciphertext_s1[60]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[59]), .CK(clk_gated), .Q(Ciphertext_s0[59]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2006), .CK(clk_gated), .Q(Ciphertext_s1[59]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[58]), .CK(clk_gated), .Q(Ciphertext_s0[58]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1946), .CK(clk_gated), .Q(Ciphertext_s1[58]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[57]), .CK(clk_gated), .Q(Ciphertext_s0[57]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2101), .CK(clk_gated), .Q(Ciphertext_s1[57]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[56]), .CK(clk_gated), .Q(Ciphertext_s0[56]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2058), .CK(clk_gated), .Q(Ciphertext_s1[56]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[55]), .CK(clk_gated), .Q(Ciphertext_s0[55]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2004), .CK(clk_gated), .Q(Ciphertext_s1[55]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[54]), .CK(clk_gated), .Q(Ciphertext_s0[54]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1944), .CK(clk_gated), .Q(Ciphertext_s1[54]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[53]), .CK(clk_gated), .Q(Ciphertext_s0[53]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2099), .CK(clk_gated), .Q(Ciphertext_s1[53]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[52]), .CK(clk_gated), .Q(Ciphertext_s0[52]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2056), .CK(clk_gated), .Q(Ciphertext_s1[52]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[51]), .CK(clk_gated), .Q(Ciphertext_s0[51]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2002), .CK(clk_gated), .Q(Ciphertext_s1[51]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[50]), .CK(clk_gated), .Q(Ciphertext_s0[50]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1942), .CK(clk_gated), .Q(Ciphertext_s1[50]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[49]), .CK(clk_gated), .Q(Ciphertext_s0[49]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2097), .CK(clk_gated), .Q(Ciphertext_s1[49]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[48]), .CK(clk_gated), .Q(Ciphertext_s0[48]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2054), .CK(clk_gated), .Q(Ciphertext_s1[48]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[47]), .CK(clk_gated), .Q(Ciphertext_s0[47]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2000), .CK(clk_gated), .Q(Ciphertext_s1[47]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[46]), .CK(clk_gated), .Q(Ciphertext_s0[46]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1940), .CK(clk_gated), .Q(Ciphertext_s1[46]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[45]), .CK(clk_gated), .Q(Ciphertext_s0[45]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2095), .CK(clk_gated), .Q(Ciphertext_s1[45]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[44]), .CK(clk_gated), .Q(Ciphertext_s0[44]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2052), .CK(clk_gated), .Q(Ciphertext_s1[44]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[43]), .CK(clk_gated), .Q(Ciphertext_s0[43]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1878), .CK(clk_gated), .Q(Ciphertext_s1[43]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[42]), .CK(clk_gated), .Q(Ciphertext_s0[42]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1825), .CK(clk_gated), .Q(Ciphertext_s1[42]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[41]), .CK(clk_gated), .Q(Ciphertext_s0[41]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1998), .CK(clk_gated), .Q(Ciphertext_s1[41]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[40]), .CK(clk_gated), .Q(Ciphertext_s0[40]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1938), .CK(clk_gated), .Q(Ciphertext_s1[40]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[39]), .CK(clk_gated), .Q(Ciphertext_s0[39]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1876), .CK(clk_gated), .Q(Ciphertext_s1[39]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[38]), .CK(clk_gated), .Q(Ciphertext_s0[38]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1823), .CK(clk_gated), .Q(Ciphertext_s1[38]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[37]), .CK(clk_gated), .Q(Ciphertext_s0[37]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1996), .CK(clk_gated), .Q(Ciphertext_s1[37]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[36]), .CK(clk_gated), .Q(Ciphertext_s0[36]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1936), .CK(clk_gated), .Q(Ciphertext_s1[36]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[35]), .CK(clk_gated), .Q(Ciphertext_s0[35]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1874), .CK(clk_gated), .Q(Ciphertext_s1[35]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[34]), .CK(clk_gated), .Q(Ciphertext_s0[34]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1821), .CK(clk_gated), .Q(Ciphertext_s1[34]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[33]), .CK(clk_gated), .Q(Ciphertext_s0[33]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1994), .CK(clk_gated), .Q(Ciphertext_s1[33]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[32]), .CK(clk_gated), .Q(Ciphertext_s0[32]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1934), .CK(clk_gated), .Q(Ciphertext_s1[32]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[31]), .CK(clk_gated), .Q(Ciphertext_s0[31]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1992), .CK(clk_gated), .Q(Ciphertext_s1[31]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[30]), .CK(clk_gated), .Q(Ciphertext_s0[30]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1932), .CK(clk_gated), .Q(Ciphertext_s1[30]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[29]), .CK(clk_gated), .Q(Ciphertext_s0[29]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2093), .CK(clk_gated), .Q(Ciphertext_s1[29]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[28]), .CK(clk_gated), .Q(Ciphertext_s0[28]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2050), .CK(clk_gated), .Q(Ciphertext_s1[28]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[27]), .CK(clk_gated), .Q(Ciphertext_s0[27]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2091), .CK(clk_gated), .Q(Ciphertext_s1[27]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[26]), .CK(clk_gated), .Q(Ciphertext_s0[26]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2048), .CK(clk_gated), .Q(Ciphertext_s1[26]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[25]), .CK(clk_gated), .Q(Ciphertext_s0[25]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2122), .CK(clk_gated), .Q(Ciphertext_s1[25]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[24]), .CK(clk_gated), .Q(Ciphertext_s0[24]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2113), .CK(clk_gated), .Q(Ciphertext_s1[24]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[23]), .CK(clk_gated), .Q(Ciphertext_s0[23]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1990), .CK(clk_gated), .Q(Ciphertext_s1[23]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[22]), .CK(clk_gated), .Q(Ciphertext_s0[22]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1930), .CK(clk_gated), .Q(Ciphertext_s1[22]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[21]), .CK(clk_gated), .Q(Ciphertext_s0[21]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2089), .CK(clk_gated), .Q(Ciphertext_s1[21]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[20]), .CK(clk_gated), .Q(Ciphertext_s0[20]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2046), .CK(clk_gated), .Q(Ciphertext_s1[20]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[19]), .CK(clk_gated), .Q(Ciphertext_s0[19]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1988), .CK(clk_gated), .Q(Ciphertext_s1[19]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[18]), .CK(clk_gated), .Q(Ciphertext_s0[18]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1928), .CK(clk_gated), .Q(Ciphertext_s1[18]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[17]), .CK(clk_gated), .Q(Ciphertext_s0[17]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2087), .CK(clk_gated), .Q(Ciphertext_s1[17]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[16]), .CK(clk_gated), .Q(Ciphertext_s0[16]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2044), .CK(clk_gated), .Q(Ciphertext_s1[16]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[15]), .CK(clk_gated), .Q(Ciphertext_s0[15]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2085), .CK(clk_gated), .Q(Ciphertext_s1[15]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[14]), .CK(clk_gated), .Q(Ciphertext_s0[14]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2042), .CK(clk_gated), .Q(Ciphertext_s1[14]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[13]), .CK(clk_gated), .Q(Ciphertext_s0[13]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2120), .CK(clk_gated), .Q(Ciphertext_s1[13]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[12]), .CK(clk_gated), .Q(Ciphertext_s0[12]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2111), .CK(clk_gated), .Q(Ciphertext_s1[12]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[11]), .CK(clk_gated), .Q(Ciphertext_s0[11]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1986), .CK(clk_gated), .Q(Ciphertext_s1[11]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[10]), .CK(clk_gated), .Q(Ciphertext_s0[10]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1926), .CK(clk_gated), .Q(Ciphertext_s1[10]), 
        .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[9]), .CK(clk_gated), .Q(Ciphertext_s0[9]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2083), .CK(clk_gated), .Q(Ciphertext_s1[9]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[8]), .CK(clk_gated), .Q(Ciphertext_s0[8]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2040), .CK(clk_gated), .Q(Ciphertext_s1[8]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[7]), .CK(clk_gated), .Q(Ciphertext_s0[7]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1984), .CK(clk_gated), .Q(Ciphertext_s1[7]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[6]), .CK(clk_gated), .Q(Ciphertext_s0[6]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1924), .CK(clk_gated), .Q(Ciphertext_s1[6]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[5]), .CK(clk_gated), .Q(Ciphertext_s0[5]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2081), .CK(clk_gated), .Q(Ciphertext_s1[5]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[4]), .CK(clk_gated), .Q(Ciphertext_s0[4]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2038), .CK(clk_gated), .Q(Ciphertext_s1[4]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[3]), .CK(clk_gated), .Q(Ciphertext_s0[3]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1982), .CK(clk_gated), .Q(Ciphertext_s1[3]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[2]), .CK(clk_gated), .Q(Ciphertext_s0[2]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1922), .CK(clk_gated), .Q(Ciphertext_s1[2]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[1]), .CK(clk_gated), .Q(Ciphertext_s0[1]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2079), .CK(clk_gated), .Q(Ciphertext_s1[1]), .QN()
         );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(StateRegInput[0]), .CK(clk_gated), .Q(Ciphertext_s0[0]), .QN() );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_2036), .CK(clk_gated), .Q(Ciphertext_s1[0]), .QN()
         );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[63]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[31]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1451), .CK(clk_gated), .Q(new_AGEMA_signal_1353), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[62]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[30]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1448), .CK(clk_gated), .Q(new_AGEMA_signal_1350), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[61]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[29]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1445), .CK(clk_gated), .Q(new_AGEMA_signal_1347), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[60]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[28]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1442), .CK(clk_gated), .Q(new_AGEMA_signal_1344), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[59]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[27]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1439), .CK(clk_gated), .Q(new_AGEMA_signal_1341), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[58]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[26]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1436), .CK(clk_gated), .Q(new_AGEMA_signal_1338), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[57]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[25]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1433), .CK(clk_gated), .Q(new_AGEMA_signal_1335), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[56]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[24]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1430), .CK(clk_gated), .Q(new_AGEMA_signal_1332), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[55]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[23]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1427), .CK(clk_gated), .Q(new_AGEMA_signal_1329), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[54]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[22]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1424), .CK(clk_gated), .Q(new_AGEMA_signal_1326), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[53]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[21]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1421), .CK(clk_gated), .Q(new_AGEMA_signal_1323), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[52]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[20]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1418), .CK(clk_gated), .Q(new_AGEMA_signal_1320), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[51]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[19]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1415), .CK(clk_gated), .Q(new_AGEMA_signal_1317), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[50]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[18]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1412), .CK(clk_gated), .Q(new_AGEMA_signal_1314), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[49]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[17]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1409), .CK(clk_gated), .Q(new_AGEMA_signal_1311), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[48]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[16]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1406), .CK(clk_gated), .Q(new_AGEMA_signal_1308), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[47]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[15]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1403), .CK(clk_gated), .Q(new_AGEMA_signal_1305), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[46]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[14]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1400), .CK(clk_gated), .Q(new_AGEMA_signal_1302), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[45]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[13]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1397), .CK(clk_gated), .Q(new_AGEMA_signal_1299), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[44]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[12]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1394), .CK(clk_gated), .Q(new_AGEMA_signal_1296), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[43]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[11]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1391), .CK(clk_gated), .Q(new_AGEMA_signal_1293), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[42]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[10]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1388), .CK(clk_gated), .Q(new_AGEMA_signal_1290), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[41]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[9]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1385), .CK(clk_gated), .Q(new_AGEMA_signal_1287), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[40]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[8]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1382), .CK(clk_gated), .Q(new_AGEMA_signal_1284), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[39]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[7]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1379), .CK(clk_gated), .Q(new_AGEMA_signal_1281), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[38]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[6]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1376), .CK(clk_gated), .Q(new_AGEMA_signal_1278), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[37]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[5]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1373), .CK(clk_gated), .Q(new_AGEMA_signal_1275), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[36]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[4]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1370), .CK(clk_gated), .Q(new_AGEMA_signal_1272), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[35]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[3]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1367), .CK(clk_gated), .Q(new_AGEMA_signal_1269), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[34]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[2]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1364), .CK(clk_gated), .Q(new_AGEMA_signal_1266), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[33]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[1]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1361), .CK(clk_gated), .Q(new_AGEMA_signal_1263), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[32]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[0]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1358), .CK(clk_gated), .Q(new_AGEMA_signal_1260), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[31]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[55]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1355), .CK(clk_gated), .Q(new_AGEMA_signal_1425), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[30]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[54]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1352), .CK(clk_gated), .Q(new_AGEMA_signal_1422), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[29]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[53]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1349), .CK(clk_gated), .Q(new_AGEMA_signal_1419), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[28]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[52]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1346), .CK(clk_gated), .Q(new_AGEMA_signal_1416), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[27]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[63]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1343), .CK(clk_gated), .Q(new_AGEMA_signal_1449), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[26]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[62]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1340), .CK(clk_gated), .Q(new_AGEMA_signal_1446), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[25]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[61]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1337), .CK(clk_gated), .Q(new_AGEMA_signal_1443), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[24]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[60]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1334), .CK(clk_gated), .Q(new_AGEMA_signal_1440), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[23]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[47]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1331), .CK(clk_gated), .Q(new_AGEMA_signal_1401), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[22]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[46]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1328), .CK(clk_gated), .Q(new_AGEMA_signal_1398), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[21]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[45]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1325), .CK(clk_gated), .Q(new_AGEMA_signal_1395), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[20]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[44]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1322), .CK(clk_gated), .Q(new_AGEMA_signal_1392), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[19]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[35]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1319), .CK(clk_gated), .Q(new_AGEMA_signal_1365), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[18]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[34]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1316), .CK(clk_gated), .Q(new_AGEMA_signal_1362), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[17]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[33]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1313), .CK(clk_gated), .Q(new_AGEMA_signal_1359), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[16]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[32]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1310), .CK(clk_gated), .Q(new_AGEMA_signal_1356), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[15]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[39]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1307), .CK(clk_gated), .Q(new_AGEMA_signal_1377), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[14]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[38]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1304), .CK(clk_gated), .Q(new_AGEMA_signal_1374), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[13]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[37]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1301), .CK(clk_gated), .Q(new_AGEMA_signal_1371), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[12]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[36]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1298), .CK(clk_gated), .Q(new_AGEMA_signal_1368), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[11]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[51]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1295), .CK(clk_gated), .Q(new_AGEMA_signal_1413), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[10]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[50]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1292), .CK(clk_gated), .Q(new_AGEMA_signal_1410), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[9]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[49]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1289), .CK(clk_gated), .Q(new_AGEMA_signal_1407), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[8]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[48]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1286), .CK(clk_gated), .Q(new_AGEMA_signal_1404), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[7]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[43]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1283), .CK(clk_gated), .Q(new_AGEMA_signal_1389), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[6]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[42]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1280), .CK(clk_gated), .Q(new_AGEMA_signal_1386), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[5]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[41]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1277), .CK(clk_gated), .Q(new_AGEMA_signal_1383), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[4]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[40]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1274), .CK(clk_gated), .Q(new_AGEMA_signal_1380), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[3]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[59]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1271), .CK(clk_gated), .Q(new_AGEMA_signal_1437), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[2]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[58]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1268), .CK(clk_gated), .Q(new_AGEMA_signal_1434), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[1]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[57]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1265), .CK(clk_gated), .Q(new_AGEMA_signal_1431), 
        .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_0_s_current_state_reg ( 
        .D(TweakeyGeneration_StateRegInput[0]), .CK(clk_gated), .Q(
        TweakeyGeneration_key_Feedback[56]), .QN() );
  DFF_X1 TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF_s_reg_1_s_current_state_reg ( 
        .D(new_AGEMA_signal_1262), .CK(clk_gated), .Q(new_AGEMA_signal_1428), 
        .QN() );
endmodule

