
module PRESENT ( clk, reset, data_in, key, data_out, done );
  (* AGEMA = "secure" *) input [63:0] data_in;
  (* AGEMA = "secure" *) input [79:0] key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input reset;

  output [63:0] data_out;
  output done;
  
  wire   selSbox, ctrlData_0_, intDone, fsm_n15, fsm_n14, fsm_n13, fsm_n12,
         fsm_n11, fsm_n10, fsm_n9, fsm_n8, fsm_n7, fsm_n6, fsm_n4, fsm_n2,
         fsm_n5, fsm_n20, fsm_ps_state_0_, fsm_ps_state_1_, fsm_n21, fsm_n3,
         fsm_rst_countSerial, fsm_en_countRound, fsm_cnt_rnd_n33,
         fsm_cnt_rnd_n32, fsm_cnt_rnd_n31, fsm_cnt_rnd_n30, fsm_cnt_rnd_n29,
         fsm_cnt_rnd_n28, fsm_cnt_rnd_n27, fsm_cnt_rnd_n26, fsm_cnt_rnd_n23,
         fsm_cnt_rnd_n22, fsm_cnt_rnd_n21, fsm_cnt_rnd_n20, fsm_cnt_rnd_n19,
         fsm_cnt_rnd_n17, fsm_cnt_rnd_n15, fsm_cnt_rnd_n13, fsm_cnt_rnd_n12,
         fsm_cnt_rnd_n11, fsm_cnt_rnd_n10, fsm_cnt_rnd_n9, fsm_cnt_rnd_n8,
         fsm_cnt_rnd_n7, fsm_cnt_rnd_n6, fsm_cnt_rnd_n5, fsm_cnt_rnd_n3,
         fsm_cnt_rnd_n24, fsm_cnt_rnd_n41, fsm_cnt_rnd_n25, fsm_cnt_rnd_n1,
         fsm_cnt_rnd_n18, fsm_cnt_rnd_n16, fsm_cnt_rnd_n14,
         fsm_cnt_rnd_count_reg_reg_4__QN, fsm_cnt_ser_n10, fsm_cnt_ser_n9,
         fsm_cnt_ser_n8, fsm_cnt_ser_n7, fsm_cnt_ser_n6, fsm_cnt_ser_n5,
         fsm_cnt_ser_n4, fsm_cnt_ser_n2, fsm_cnt_ser_n20, fsm_cnt_ser_n28,
         fsm_cnt_ser_n26, fsm_cnt_ser_n3, fsm_cnt_ser_n1,
         fsm_cnt_ser_count_reg_reg_2__QN, fsm_cnt_ser_count_reg_reg_0__QN,
         fsm_cnt_ser_count_reg_reg_3__QN, stateFF_state_n7, stateFF_state_n6,
         stateFF_state_n5, stateFF_state_gff_1_s_current_state_reg_0__QN,
         stateFF_state_gff_1_s_current_state_reg_2__QN,
         stateFF_state_gff_1_s_current_state_reg_1__QN,
         stateFF_state_gff_1_s_current_state_reg_3__QN,
         stateFF_state_gff_2_s_current_state_reg_3__QN,
         stateFF_state_gff_2_s_current_state_reg_2__QN,
         stateFF_state_gff_2_s_current_state_reg_1__QN,
         stateFF_state_gff_2_s_current_state_reg_0__QN,
         stateFF_state_gff_3_s_current_state_reg_3__QN,
         stateFF_state_gff_3_s_current_state_reg_2__QN,
         stateFF_state_gff_3_s_current_state_reg_1__QN,
         stateFF_state_gff_3_s_current_state_reg_0__QN,
         stateFF_state_gff_4_s_current_state_reg_3__QN,
         stateFF_state_gff_4_s_current_state_reg_2__QN,
         stateFF_state_gff_4_s_current_state_reg_1__QN,
         stateFF_state_gff_4_s_current_state_reg_0__QN,
         stateFF_state_gff_5_s_current_state_reg_3__QN,
         stateFF_state_gff_5_s_current_state_reg_2__QN,
         stateFF_state_gff_5_s_current_state_reg_1__QN,
         stateFF_state_gff_5_s_current_state_reg_0__QN,
         stateFF_state_gff_6_s_current_state_reg_3__QN,
         stateFF_state_gff_6_s_current_state_reg_2__QN,
         stateFF_state_gff_6_s_current_state_reg_1__QN,
         stateFF_state_gff_6_s_current_state_reg_0__QN,
         stateFF_state_gff_7_s_current_state_reg_3__QN,
         stateFF_state_gff_7_s_current_state_reg_2__QN,
         stateFF_state_gff_7_s_current_state_reg_1__QN,
         stateFF_state_gff_7_s_current_state_reg_0__QN,
         stateFF_state_gff_8_s_current_state_reg_3__QN,
         stateFF_state_gff_8_s_current_state_reg_2__QN,
         stateFF_state_gff_8_s_current_state_reg_1__QN,
         stateFF_state_gff_8_s_current_state_reg_0__QN,
         stateFF_state_gff_9_s_current_state_reg_3__QN,
         stateFF_state_gff_9_s_current_state_reg_2__QN,
         stateFF_state_gff_9_s_current_state_reg_1__QN,
         stateFF_state_gff_9_s_current_state_reg_0__QN,
         stateFF_state_gff_10_s_current_state_reg_3__QN,
         stateFF_state_gff_10_s_current_state_reg_2__QN,
         stateFF_state_gff_10_s_current_state_reg_1__QN,
         stateFF_state_gff_10_s_current_state_reg_0__QN,
         stateFF_state_gff_11_s_current_state_reg_3__QN,
         stateFF_state_gff_11_s_current_state_reg_2__QN,
         stateFF_state_gff_11_s_current_state_reg_1__QN,
         stateFF_state_gff_11_s_current_state_reg_0__QN,
         stateFF_state_gff_12_s_current_state_reg_3__QN,
         stateFF_state_gff_12_s_current_state_reg_2__QN,
         stateFF_state_gff_12_s_current_state_reg_1__QN,
         stateFF_state_gff_12_s_current_state_reg_0__QN,
         stateFF_state_gff_13_s_current_state_reg_3__QN,
         stateFF_state_gff_13_s_current_state_reg_2__QN,
         stateFF_state_gff_13_s_current_state_reg_1__QN,
         stateFF_state_gff_13_s_current_state_reg_0__QN,
         stateFF_state_gff_14_s_current_state_reg_3__QN,
         stateFF_state_gff_14_s_current_state_reg_2__QN,
         stateFF_state_gff_14_s_current_state_reg_1__QN,
         stateFF_state_gff_14_s_current_state_reg_0__QN,
         stateFF_state_gff_15_s_current_state_reg_3__QN,
         stateFF_state_gff_15_s_current_state_reg_2__QN,
         stateFF_state_gff_15_s_current_state_reg_1__QN,
         stateFF_state_gff_15_s_current_state_reg_0__QN,
         stateFF_state_gff_16_s_current_state_reg_3__QN,
         stateFF_state_gff_16_s_current_state_reg_2__QN,
         stateFF_state_gff_16_s_current_state_reg_1__QN,
         stateFF_state_gff_16_s_current_state_reg_0__QN, keyFF_keystate_n8,
         keyFF_keystate_n7, keyFF_keystate_n6,
         keyFF_keystate_gff_1_s_current_state_reg_3__QN,
         keyFF_keystate_gff_1_s_current_state_reg_2__QN,
         keyFF_keystate_gff_1_s_current_state_reg_1__QN,
         keyFF_keystate_gff_1_s_current_state_reg_0__QN,
         keyFF_keystate_gff_2_s_current_state_reg_3__QN,
         keyFF_keystate_gff_2_s_current_state_reg_2__QN,
         keyFF_keystate_gff_2_s_current_state_reg_1__QN,
         keyFF_keystate_gff_2_s_current_state_reg_0__QN,
         keyFF_keystate_gff_3_s_current_state_reg_3__QN,
         keyFF_keystate_gff_3_s_current_state_reg_2__QN,
         keyFF_keystate_gff_3_s_current_state_reg_1__QN,
         keyFF_keystate_gff_3_s_current_state_reg_0__QN,
         keyFF_keystate_gff_4_s_current_state_reg_3__QN,
         keyFF_keystate_gff_4_s_current_state_reg_2__QN,
         keyFF_keystate_gff_4_s_current_state_reg_1__QN,
         keyFF_keystate_gff_4_s_current_state_reg_0__QN,
         keyFF_keystate_gff_5_s_current_state_reg_3__QN,
         keyFF_keystate_gff_5_s_current_state_reg_2__QN,
         keyFF_keystate_gff_5_s_current_state_reg_1__QN,
         keyFF_keystate_gff_5_s_current_state_reg_0__QN,
         keyFF_keystate_gff_6_s_current_state_reg_3__QN,
         keyFF_keystate_gff_6_s_current_state_reg_2__QN,
         keyFF_keystate_gff_6_s_current_state_reg_1__QN,
         keyFF_keystate_gff_6_s_current_state_reg_0__QN,
         keyFF_keystate_gff_7_s_current_state_reg_3__QN,
         keyFF_keystate_gff_7_s_current_state_reg_2__QN,
         keyFF_keystate_gff_7_s_current_state_reg_1__QN,
         keyFF_keystate_gff_7_s_current_state_reg_0__QN,
         keyFF_keystate_gff_8_s_current_state_reg_3__QN,
         keyFF_keystate_gff_8_s_current_state_reg_2__QN,
         keyFF_keystate_gff_8_s_current_state_reg_1__QN,
         keyFF_keystate_gff_8_s_current_state_reg_0__QN,
         keyFF_keystate_gff_9_s_current_state_reg_3__QN,
         keyFF_keystate_gff_9_s_current_state_reg_2__QN,
         keyFF_keystate_gff_9_s_current_state_reg_1__QN,
         keyFF_keystate_gff_9_s_current_state_reg_0__QN,
         keyFF_keystate_gff_10_s_current_state_reg_3__QN,
         keyFF_keystate_gff_10_s_current_state_reg_2__QN,
         keyFF_keystate_gff_10_s_current_state_reg_1__QN,
         keyFF_keystate_gff_10_s_current_state_reg_0__QN,
         keyFF_keystate_gff_11_s_current_state_reg_3__QN,
         keyFF_keystate_gff_11_s_current_state_reg_2__QN,
         keyFF_keystate_gff_11_s_current_state_reg_1__QN,
         keyFF_keystate_gff_11_s_current_state_reg_0__QN,
         keyFF_keystate_gff_12_s_current_state_reg_3__QN,
         keyFF_keystate_gff_12_s_current_state_reg_2__QN,
         keyFF_keystate_gff_12_s_current_state_reg_1__QN,
         keyFF_keystate_gff_12_s_current_state_reg_0__QN,
         keyFF_keystate_gff_13_s_current_state_reg_3__QN,
         keyFF_keystate_gff_13_s_current_state_reg_2__QN,
         keyFF_keystate_gff_13_s_current_state_reg_1__QN,
         keyFF_keystate_gff_13_s_current_state_reg_0__QN,
         keyFF_keystate_gff_14_s_current_state_reg_3__QN,
         keyFF_keystate_gff_14_s_current_state_reg_2__QN,
         keyFF_keystate_gff_14_s_current_state_reg_1__QN,
         keyFF_keystate_gff_14_s_current_state_reg_0__QN,
         keyFF_keystate_gff_15_s_current_state_reg_3__QN,
         keyFF_keystate_gff_15_s_current_state_reg_2__QN,
         keyFF_keystate_gff_15_s_current_state_reg_1__QN,
         keyFF_keystate_gff_15_s_current_state_reg_0__QN,
         keyFF_keystate_gff_16_s_current_state_reg_3__QN,
         keyFF_keystate_gff_16_s_current_state_reg_2__QN,
         keyFF_keystate_gff_16_s_current_state_reg_1__QN,
         keyFF_keystate_gff_16_s_current_state_reg_0__QN,
         keyFF_keystate_gff_17_s_current_state_reg_3__QN,
         keyFF_keystate_gff_17_s_current_state_reg_2__QN,
         keyFF_keystate_gff_17_s_current_state_reg_1__QN,
         keyFF_keystate_gff_17_s_current_state_reg_0__QN,
         keyFF_keystate_gff_18_s_current_state_reg_3__QN,
         keyFF_keystate_gff_18_s_current_state_reg_2__QN,
         keyFF_keystate_gff_18_s_current_state_reg_1__QN,
         keyFF_keystate_gff_18_s_current_state_reg_0__QN,
         keyFF_keystate_gff_19_s_current_state_reg_3__QN,
         keyFF_keystate_gff_19_s_current_state_reg_2__QN,
         keyFF_keystate_gff_19_s_current_state_reg_1__QN,
         keyFF_keystate_gff_19_s_current_state_reg_0__QN,
         keyFF_keystate_gff_20_s_current_state_reg_3__QN,
         keyFF_keystate_gff_20_s_current_state_reg_2__QN,
         keyFF_keystate_gff_20_s_current_state_reg_1__QN,
         keyFF_keystate_gff_20_s_current_state_reg_0__QN, sboxInst_n3,
         sboxInst_n2, sboxInst_n1, sboxInst_L8, sboxInst_L7, sboxInst_T3,
         sboxInst_T1, sboxInst_Q7, sboxInst_Q6, sboxInst_L5, sboxInst_T2,
         sboxInst_L4, sboxInst_Q3, sboxInst_L3, sboxInst_Q2, sboxInst_T0,
         sboxInst_L2, sboxInst_L1, sboxInst_L0;
  wire   [4:0] counter;
  wire   [3:0] serialIn;
  wire   [3:0] sboxOut;
  wire   [3:0] roundkey;
  wire   [3:1] keyRegKS;
  wire   [3:0] sboxIn;
  wire   [3:0] stateXORroundkey;
  wire   [3:0] fsm_countSerial;
  wire   [63:0] stateFF_inputPar;
  wire   [3:0] stateFF_state_gff_1_s_next_state;
  wire   [3:0] stateFF_state_gff_2_s_next_state;
  wire   [3:0] stateFF_state_gff_3_s_next_state;
  wire   [3:0] stateFF_state_gff_4_s_next_state;
  wire   [3:0] stateFF_state_gff_5_s_next_state;
  wire   [3:0] stateFF_state_gff_6_s_next_state;
  wire   [3:0] stateFF_state_gff_7_s_next_state;
  wire   [3:0] stateFF_state_gff_8_s_next_state;
  wire   [3:0] stateFF_state_gff_9_s_next_state;
  wire   [3:0] stateFF_state_gff_10_s_next_state;
  wire   [3:0] stateFF_state_gff_11_s_next_state;
  wire   [3:0] stateFF_state_gff_12_s_next_state;
  wire   [3:0] stateFF_state_gff_13_s_next_state;
  wire   [3:0] stateFF_state_gff_14_s_next_state;
  wire   [3:0] stateFF_state_gff_15_s_next_state;
  wire   [3:0] stateFF_state_gff_16_s_next_state;
  wire   [4:0] keyFF_counterAdd;
  wire   [75:3] keyFF_outputPar;
  wire   [79:0] keyFF_inputPar;
  wire   [3:0] keyFF_keystate_gff_1_s_next_state;
  wire   [3:0] keyFF_keystate_gff_2_s_next_state;
  wire   [3:0] keyFF_keystate_gff_3_s_next_state;
  wire   [3:0] keyFF_keystate_gff_4_s_next_state;
  wire   [3:0] keyFF_keystate_gff_5_s_next_state;
  wire   [3:0] keyFF_keystate_gff_6_s_next_state;
  wire   [3:0] keyFF_keystate_gff_7_s_next_state;
  wire   [3:0] keyFF_keystate_gff_8_s_next_state;
  wire   [3:0] keyFF_keystate_gff_9_s_next_state;
  wire   [3:0] keyFF_keystate_gff_10_s_next_state;
  wire   [3:0] keyFF_keystate_gff_11_s_next_state;
  wire   [3:0] keyFF_keystate_gff_12_s_next_state;
  wire   [3:0] keyFF_keystate_gff_13_s_next_state;
  wire   [3:0] keyFF_keystate_gff_14_s_next_state;
  wire   [3:0] keyFF_keystate_gff_15_s_next_state;
  wire   [3:0] keyFF_keystate_gff_16_s_next_state;
  wire   [3:0] keyFF_keystate_gff_17_s_next_state;
  wire   [3:0] keyFF_keystate_gff_18_s_next_state;
  wire   [3:0] keyFF_keystate_gff_19_s_next_state;
  wire   [3:0] keyFF_keystate_gff_20_s_next_state;

  XOR2_X1 U9 ( .A(roundkey[0]), .B(data_out[60]), .Z(stateXORroundkey[0]) );
  XOR2_X1 U10 ( .A(roundkey[1]), .B(data_out[61]), .Z(stateXORroundkey[1]) );
  XOR2_X1 U11 ( .A(roundkey[2]), .B(data_out[62]), .Z(stateXORroundkey[2]) );
  XOR2_X1 U12 ( .A(roundkey[3]), .B(data_out[63]), .Z(stateXORroundkey[3]) );
  NOR2_X1 fsm_U20 ( .A1(reset), .A2(fsm_n15), .ZN(fsm_n21) );
  NOR2_X1 fsm_U19 ( .A1(fsm_n14), .A2(done), .ZN(fsm_n15) );
  NOR2_X1 fsm_U18 ( .A1(reset), .A2(fsm_n13), .ZN(fsm_n20) );
  NOR2_X1 fsm_U17 ( .A1(fsm_ps_state_1_), .A2(fsm_n12), .ZN(fsm_n13) );
  NOR2_X1 fsm_U16 ( .A1(fsm_n11), .A2(fsm_n10), .ZN(fsm_n12) );
  NAND2_X1 fsm_U15 ( .A1(counter[3]), .A2(counter[1]), .ZN(fsm_n10) );
  OR2_X1 fsm_U14 ( .A1(fsm_n9), .A2(fsm_n8), .ZN(fsm_n11) );
  NAND2_X1 fsm_U13 ( .A1(counter[0]), .A2(counter[4]), .ZN(fsm_n8) );
  NAND2_X1 fsm_U12 ( .A1(counter[2]), .A2(fsm_ps_state_0_), .ZN(fsm_n9) );
  NOR2_X1 fsm_U11 ( .A1(fsm_n3), .A2(fsm_n5), .ZN(done) );
  AND2_X1 fsm_U10 ( .A1(fsm_n14), .A2(fsm_n5), .ZN(fsm_en_countRound) );
  AND2_X1 fsm_U9 ( .A1(fsm_countSerial[2]), .A2(fsm_n7), .ZN(fsm_n14) );
  NOR2_X1 fsm_U8 ( .A1(fsm_n6), .A2(fsm_n4), .ZN(fsm_n7) );
  NAND2_X1 fsm_U7 ( .A1(fsm_countSerial[1]), .A2(fsm_countSerial[0]), .ZN(
        fsm_n4) );
  NAND2_X1 fsm_U6 ( .A1(fsm_n3), .A2(fsm_countSerial[3]), .ZN(fsm_n6) );
  NOR2_X1 fsm_U5 ( .A1(fsm_ps_state_0_), .A2(fsm_n5), .ZN(intDone) );
  NOR2_X1 fsm_U4 ( .A1(fsm_ps_state_1_), .A2(fsm_n3), .ZN(selSbox) );
  NOR2_X1 fsm_U3 ( .A1(reset), .A2(selSbox), .ZN(fsm_rst_countSerial) );
  INV_X1 fsm_U2 ( .A(reset), .ZN(fsm_n2) );
  INV_X1 fsm_U1 ( .A(fsm_rst_countSerial), .ZN(ctrlData_0_) );
  NAND2_X1 fsm_cnt_rnd_U28 ( .A1(fsm_cnt_rnd_n33), .A2(fsm_cnt_rnd_n32), .ZN(
        fsm_cnt_rnd_n41) );
  NAND2_X1 fsm_cnt_rnd_U27 ( .A1(fsm_cnt_rnd_n31), .A2(counter[1]), .ZN(
        fsm_cnt_rnd_n32) );
  NAND2_X1 fsm_cnt_rnd_U26 ( .A1(fsm_cnt_rnd_n30), .A2(fsm_cnt_rnd_n24), .ZN(
        fsm_cnt_rnd_n33) );
  NAND2_X1 fsm_cnt_rnd_U25 ( .A1(fsm_cnt_rnd_n29), .A2(counter[0]), .ZN(
        fsm_cnt_rnd_n30) );
  NAND2_X1 fsm_cnt_rnd_U24 ( .A1(fsm_cnt_rnd_n28), .A2(fsm_cnt_rnd_n27), .ZN(
        fsm_cnt_rnd_n18) );
  NAND2_X1 fsm_cnt_rnd_U23 ( .A1(fsm_cnt_rnd_n26), .A2(counter[0]), .ZN(
        fsm_cnt_rnd_n27) );
  MUX2_X1 fsm_cnt_rnd_U22 ( .A(fsm_cnt_rnd_n23), .B(fsm_cnt_rnd_n22), .S(
        fsm_cnt_rnd_n5), .Z(fsm_cnt_rnd_n16) );
  NAND2_X1 fsm_cnt_rnd_U21 ( .A1(fsm_cnt_rnd_n31), .A2(fsm_cnt_rnd_n21), .ZN(
        fsm_cnt_rnd_n23) );
  NAND2_X1 fsm_cnt_rnd_U20 ( .A1(fsm_cnt_rnd_n29), .A2(fsm_cnt_rnd_n24), .ZN(
        fsm_cnt_rnd_n21) );
  NOR2_X1 fsm_cnt_rnd_U19 ( .A1(fsm_cnt_rnd_n20), .A2(fsm_cnt_rnd_n26), .ZN(
        fsm_cnt_rnd_n31) );
  NOR2_X1 fsm_cnt_rnd_U18 ( .A1(fsm_en_countRound), .A2(fsm_cnt_rnd_n6), .ZN(
        fsm_cnt_rnd_n26) );
  INV_X1 fsm_cnt_rnd_U17 ( .A(fsm_cnt_rnd_n28), .ZN(fsm_cnt_rnd_n20) );
  NAND2_X1 fsm_cnt_rnd_U16 ( .A1(fsm_cnt_rnd_n29), .A2(fsm_cnt_rnd_n3), .ZN(
        fsm_cnt_rnd_n28) );
  MUX2_X1 fsm_cnt_rnd_U15 ( .A(fsm_cnt_rnd_n19), .B(fsm_cnt_rnd_n17), .S(
        counter[4]), .Z(fsm_cnt_rnd_n14) );
  NAND2_X1 fsm_cnt_rnd_U14 ( .A1(fsm_cnt_rnd_n15), .A2(fsm_cnt_rnd_n13), .ZN(
        fsm_cnt_rnd_n17) );
  NAND2_X1 fsm_cnt_rnd_U13 ( .A1(fsm_cnt_rnd_n29), .A2(fsm_cnt_rnd_n25), .ZN(
        fsm_cnt_rnd_n15) );
  INV_X1 fsm_cnt_rnd_U12 ( .A(fsm_cnt_rnd_n12), .ZN(fsm_cnt_rnd_n29) );
  NOR2_X1 fsm_cnt_rnd_U11 ( .A1(fsm_cnt_rnd_n25), .A2(fsm_cnt_rnd_n11), .ZN(
        fsm_cnt_rnd_n19) );
  INV_X1 fsm_cnt_rnd_U10 ( .A(fsm_cnt_rnd_n10), .ZN(fsm_cnt_rnd_n1) );
  MUX2_X1 fsm_cnt_rnd_U9 ( .A(fsm_cnt_rnd_n13), .B(fsm_cnt_rnd_n11), .S(
        fsm_cnt_rnd_n25), .Z(fsm_cnt_rnd_n10) );
  NAND2_X1 fsm_cnt_rnd_U8 ( .A1(counter[2]), .A2(fsm_cnt_rnd_n22), .ZN(
        fsm_cnt_rnd_n11) );
  NOR2_X1 fsm_cnt_rnd_U7 ( .A1(fsm_cnt_rnd_n12), .A2(fsm_cnt_rnd_n9), .ZN(
        fsm_cnt_rnd_n22) );
  NAND2_X1 fsm_cnt_rnd_U6 ( .A1(fsm_en_countRound), .A2(fsm_n2), .ZN(
        fsm_cnt_rnd_n12) );
  NAND2_X1 fsm_cnt_rnd_U5 ( .A1(fsm_n2), .A2(fsm_cnt_rnd_n8), .ZN(
        fsm_cnt_rnd_n13) );
  NAND2_X1 fsm_cnt_rnd_U4 ( .A1(fsm_en_countRound), .A2(fsm_cnt_rnd_n7), .ZN(
        fsm_cnt_rnd_n8) );
  NOR2_X1 fsm_cnt_rnd_U3 ( .A1(fsm_cnt_rnd_n5), .A2(fsm_cnt_rnd_n9), .ZN(
        fsm_cnt_rnd_n7) );
  OR2_X1 fsm_cnt_rnd_U2 ( .A1(fsm_cnt_rnd_n24), .A2(fsm_cnt_rnd_n3), .ZN(
        fsm_cnt_rnd_n9) );
  INV_X1 fsm_cnt_rnd_U1 ( .A(fsm_n2), .ZN(fsm_cnt_rnd_n6) );
  INV_X1 fsm_cnt_rnd_count_reg_reg_4__U1 ( .A(counter[4]), .ZN(
        fsm_cnt_rnd_count_reg_reg_4__QN) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_4__FF_FF ( .D(fsm_cnt_rnd_n14), .CK(clk), 
        .Q(counter[4]), .QN() );
  INV_X1 fsm_cnt_rnd_count_reg_reg_2__U1 ( .A(counter[2]), .ZN(fsm_cnt_rnd_n5)
         );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_2__FF_FF ( .D(fsm_cnt_rnd_n16), .CK(clk), 
        .Q(counter[2]), .QN() );
  INV_X1 fsm_cnt_rnd_count_reg_reg_0__U1 ( .A(counter[0]), .ZN(fsm_cnt_rnd_n3)
         );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_0__FF_FF ( .D(fsm_cnt_rnd_n18), .CK(clk), 
        .Q(counter[0]), .QN() );
  INV_X1 fsm_cnt_rnd_count_reg_reg_3__U1 ( .A(counter[3]), .ZN(fsm_cnt_rnd_n25) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_3__FF_FF ( .D(fsm_cnt_rnd_n1), .CK(clk), 
        .Q(counter[3]), .QN() );
  INV_X1 fsm_cnt_rnd_count_reg_reg_1__U1 ( .A(fsm_cnt_rnd_n24), .ZN(counter[1]) );
  DFF_X1 fsm_cnt_rnd_count_reg_reg_1__FF_FF ( .D(fsm_cnt_rnd_n41), .CK(clk), 
        .Q(fsm_cnt_rnd_n24), .QN() );
  NOR2_X1 fsm_cnt_ser_U12 ( .A1(fsm_cnt_ser_n10), .A2(fsm_cnt_ser_n9), .ZN(
        fsm_cnt_ser_n3) );
  XNOR2_X1 fsm_cnt_ser_U11 ( .A(fsm_n3), .B(fsm_countSerial[0]), .ZN(
        fsm_cnt_ser_n10) );
  NOR2_X1 fsm_cnt_ser_U10 ( .A1(fsm_cnt_ser_n9), .A2(fsm_cnt_ser_n8), .ZN(
        fsm_cnt_ser_n28) );
  XOR2_X1 fsm_cnt_ser_U9 ( .A(fsm_countSerial[1]), .B(fsm_cnt_ser_n7), .Z(
        fsm_cnt_ser_n8) );
  NOR2_X1 fsm_cnt_ser_U8 ( .A1(fsm_cnt_ser_n9), .A2(fsm_cnt_ser_n6), .ZN(
        fsm_cnt_ser_n26) );
  XOR2_X1 fsm_cnt_ser_U7 ( .A(fsm_countSerial[3]), .B(fsm_cnt_ser_n5), .Z(
        fsm_cnt_ser_n6) );
  NAND2_X1 fsm_cnt_ser_U6 ( .A1(fsm_cnt_ser_n4), .A2(fsm_countSerial[2]), .ZN(
        fsm_cnt_ser_n5) );
  NOR2_X1 fsm_cnt_ser_U5 ( .A1(fsm_cnt_ser_n2), .A2(fsm_cnt_ser_n9), .ZN(
        fsm_cnt_ser_n1) );
  INV_X1 fsm_cnt_ser_U4 ( .A(fsm_rst_countSerial), .ZN(fsm_cnt_ser_n9) );
  XNOR2_X1 fsm_cnt_ser_U3 ( .A(fsm_cnt_ser_n4), .B(fsm_countSerial[2]), .ZN(
        fsm_cnt_ser_n2) );
  NOR2_X1 fsm_cnt_ser_U2 ( .A1(fsm_cnt_ser_n20), .A2(fsm_cnt_ser_n7), .ZN(
        fsm_cnt_ser_n4) );
  NAND2_X1 fsm_cnt_ser_U1 ( .A1(fsm_n3), .A2(fsm_countSerial[0]), .ZN(
        fsm_cnt_ser_n7) );
  INV_X1 fsm_cnt_ser_count_reg_reg_2__U1 ( .A(fsm_countSerial[2]), .ZN(
        fsm_cnt_ser_count_reg_reg_2__QN) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_2__FF_FF ( .D(fsm_cnt_ser_n1), .CK(clk), 
        .Q(fsm_countSerial[2]), .QN() );
  INV_X1 fsm_cnt_ser_count_reg_reg_0__U1 ( .A(fsm_countSerial[0]), .ZN(
        fsm_cnt_ser_count_reg_reg_0__QN) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_0__FF_FF ( .D(fsm_cnt_ser_n3), .CK(clk), 
        .Q(fsm_countSerial[0]), .QN() );
  INV_X1 fsm_cnt_ser_count_reg_reg_3__U1 ( .A(fsm_countSerial[3]), .ZN(
        fsm_cnt_ser_count_reg_reg_3__QN) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_3__FF_FF ( .D(fsm_cnt_ser_n26), .CK(clk), 
        .Q(fsm_countSerial[3]), .QN() );
  INV_X1 fsm_cnt_ser_count_reg_reg_1__U1 ( .A(fsm_countSerial[1]), .ZN(
        fsm_cnt_ser_n20) );
  DFF_X1 fsm_cnt_ser_count_reg_reg_1__FF_FF ( .D(fsm_cnt_ser_n28), .CK(clk), 
        .Q(fsm_countSerial[1]), .QN() );
  INV_X1 fsm_ps_state_reg_0__U1 ( .A(fsm_ps_state_0_), .ZN(fsm_n3) );
  DFF_X1 fsm_ps_state_reg_0__FF_FF ( .D(fsm_n21), .CK(clk), .Q(fsm_ps_state_0_), .QN() );
  INV_X1 fsm_ps_state_reg_1__U1 ( .A(fsm_ps_state_1_), .ZN(fsm_n5) );
  DFF_X1 fsm_ps_state_reg_1__FF_FF ( .D(fsm_n20), .CK(clk), .Q(fsm_ps_state_1_), .QN() );
  INV_X2 stateFF_state_U3 ( .A(stateFF_state_n7), .ZN(stateFF_state_n6) );
  INV_X2 stateFF_state_U2 ( .A(stateFF_state_n7), .ZN(stateFF_state_n5) );
  INV_X1 stateFF_state_U1 ( .A(ctrlData_0_), .ZN(stateFF_state_n7) );
  MUX2_X1 stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1 ( .A(serialIn[0]), .B(
        stateFF_inputPar[0]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_1_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1 ( .A(serialIn[1]), .B(
        stateFF_inputPar[1]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_1_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1 ( .A(serialIn[2]), .B(
        stateFF_inputPar[2]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_1_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1 ( .A(serialIn[3]), .B(
        stateFF_inputPar[3]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_1_s_next_state[3]) );
  INV_X1 stateFF_state_gff_1_s_current_state_reg_0__U1 ( .A(data_out[0]), .ZN(
        stateFF_state_gff_1_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_1_s_next_state[0]), .CK(clk), .Q(data_out[0]), .QN()
         );
  INV_X1 stateFF_state_gff_1_s_current_state_reg_2__U1 ( .A(data_out[2]), .ZN(
        stateFF_state_gff_1_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_1_s_next_state[2]), .CK(clk), .Q(data_out[2]), .QN()
         );
  INV_X1 stateFF_state_gff_1_s_current_state_reg_1__U1 ( .A(data_out[1]), .ZN(
        stateFF_state_gff_1_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_1_s_next_state[1]), .CK(clk), .Q(data_out[1]), .QN()
         );
  INV_X1 stateFF_state_gff_1_s_current_state_reg_3__U1 ( .A(data_out[3]), .ZN(
        stateFF_state_gff_1_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_1_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_1_s_next_state[3]), .CK(clk), .Q(data_out[3]), .QN()
         );
  INV_X1 stateFF_state_gff_2_s_current_state_reg_3__U1 ( .A(data_out[7]), .ZN(
        stateFF_state_gff_2_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_2_s_next_state[3]), .CK(clk), .Q(data_out[7]), .QN()
         );
  INV_X1 stateFF_state_gff_2_s_current_state_reg_2__U1 ( .A(data_out[6]), .ZN(
        stateFF_state_gff_2_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_2_s_next_state[2]), .CK(clk), .Q(data_out[6]), .QN()
         );
  INV_X1 stateFF_state_gff_2_s_current_state_reg_1__U1 ( .A(data_out[5]), .ZN(
        stateFF_state_gff_2_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_2_s_next_state[1]), .CK(clk), .Q(data_out[5]), .QN()
         );
  INV_X1 stateFF_state_gff_2_s_current_state_reg_0__U1 ( .A(data_out[4]), .ZN(
        stateFF_state_gff_2_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_2_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_2_s_next_state[0]), .CK(clk), .Q(data_out[4]), .QN()
         );
  MUX2_X1 stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1 ( .A(data_out[0]), .B(
        stateFF_inputPar[4]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_2_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1 ( .A(data_out[1]), .B(
        stateFF_inputPar[5]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_2_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1 ( .A(data_out[2]), .B(
        stateFF_inputPar[6]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_2_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1 ( .A(data_out[3]), .B(
        stateFF_inputPar[7]), .S(ctrlData_0_), .Z(
        stateFF_state_gff_2_s_next_state[3]) );
  INV_X1 stateFF_state_gff_3_s_current_state_reg_3__U1 ( .A(data_out[11]), 
        .ZN(stateFF_state_gff_3_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_3_s_next_state[3]), .CK(clk), .Q(data_out[11]), 
        .QN() );
  INV_X1 stateFF_state_gff_3_s_current_state_reg_2__U1 ( .A(data_out[10]), 
        .ZN(stateFF_state_gff_3_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_3_s_next_state[2]), .CK(clk), .Q(data_out[10]), 
        .QN() );
  INV_X1 stateFF_state_gff_3_s_current_state_reg_1__U1 ( .A(data_out[9]), .ZN(
        stateFF_state_gff_3_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_3_s_next_state[1]), .CK(clk), .Q(data_out[9]), .QN()
         );
  INV_X1 stateFF_state_gff_3_s_current_state_reg_0__U1 ( .A(data_out[8]), .ZN(
        stateFF_state_gff_3_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_3_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_3_s_next_state[0]), .CK(clk), .Q(data_out[8]), .QN()
         );
  MUX2_X1 stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1 ( .A(data_out[4]), .B(
        stateFF_inputPar[8]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_3_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1 ( .A(data_out[5]), .B(
        stateFF_inputPar[9]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_3_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1 ( .A(data_out[6]), .B(
        stateFF_inputPar[10]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_3_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1 ( .A(data_out[7]), .B(
        stateFF_inputPar[11]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_3_s_next_state[3]) );
  INV_X1 stateFF_state_gff_4_s_current_state_reg_3__U1 ( .A(data_out[15]), 
        .ZN(stateFF_state_gff_4_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_4_s_next_state[3]), .CK(clk), .Q(data_out[15]), 
        .QN() );
  INV_X1 stateFF_state_gff_4_s_current_state_reg_2__U1 ( .A(data_out[14]), 
        .ZN(stateFF_state_gff_4_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_4_s_next_state[2]), .CK(clk), .Q(data_out[14]), 
        .QN() );
  INV_X1 stateFF_state_gff_4_s_current_state_reg_1__U1 ( .A(data_out[13]), 
        .ZN(stateFF_state_gff_4_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_4_s_next_state[1]), .CK(clk), .Q(data_out[13]), 
        .QN() );
  INV_X1 stateFF_state_gff_4_s_current_state_reg_0__U1 ( .A(data_out[12]), 
        .ZN(stateFF_state_gff_4_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_4_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_4_s_next_state[0]), .CK(clk), .Q(data_out[12]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1 ( .A(data_out[8]), .B(
        stateFF_inputPar[12]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_4_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1 ( .A(data_out[9]), .B(
        stateFF_inputPar[13]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_4_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1 ( .A(data_out[10]), .B(
        stateFF_inputPar[14]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_4_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1 ( .A(data_out[11]), .B(
        stateFF_inputPar[15]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_4_s_next_state[3]) );
  INV_X1 stateFF_state_gff_5_s_current_state_reg_3__U1 ( .A(data_out[19]), 
        .ZN(stateFF_state_gff_5_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_5_s_next_state[3]), .CK(clk), .Q(data_out[19]), 
        .QN() );
  INV_X1 stateFF_state_gff_5_s_current_state_reg_2__U1 ( .A(data_out[18]), 
        .ZN(stateFF_state_gff_5_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_5_s_next_state[2]), .CK(clk), .Q(data_out[18]), 
        .QN() );
  INV_X1 stateFF_state_gff_5_s_current_state_reg_1__U1 ( .A(data_out[17]), 
        .ZN(stateFF_state_gff_5_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_5_s_next_state[1]), .CK(clk), .Q(data_out[17]), 
        .QN() );
  INV_X1 stateFF_state_gff_5_s_current_state_reg_0__U1 ( .A(data_out[16]), 
        .ZN(stateFF_state_gff_5_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_5_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_5_s_next_state[0]), .CK(clk), .Q(data_out[16]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1 ( .A(data_out[12]), .B(
        stateFF_inputPar[16]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_5_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1 ( .A(data_out[13]), .B(
        stateFF_inputPar[17]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_5_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1 ( .A(data_out[14]), .B(
        stateFF_inputPar[18]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_5_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1 ( .A(data_out[15]), .B(
        stateFF_inputPar[19]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_5_s_next_state[3]) );
  INV_X1 stateFF_state_gff_6_s_current_state_reg_3__U1 ( .A(data_out[23]), 
        .ZN(stateFF_state_gff_6_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_6_s_next_state[3]), .CK(clk), .Q(data_out[23]), 
        .QN() );
  INV_X1 stateFF_state_gff_6_s_current_state_reg_2__U1 ( .A(data_out[22]), 
        .ZN(stateFF_state_gff_6_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_6_s_next_state[2]), .CK(clk), .Q(data_out[22]), 
        .QN() );
  INV_X1 stateFF_state_gff_6_s_current_state_reg_1__U1 ( .A(data_out[21]), 
        .ZN(stateFF_state_gff_6_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_6_s_next_state[1]), .CK(clk), .Q(data_out[21]), 
        .QN() );
  INV_X1 stateFF_state_gff_6_s_current_state_reg_0__U1 ( .A(data_out[20]), 
        .ZN(stateFF_state_gff_6_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_6_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_6_s_next_state[0]), .CK(clk), .Q(data_out[20]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1 ( .A(data_out[16]), .B(
        stateFF_inputPar[20]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_6_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1 ( .A(data_out[17]), .B(
        stateFF_inputPar[21]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_6_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1 ( .A(data_out[18]), .B(
        stateFF_inputPar[22]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_6_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1 ( .A(data_out[19]), .B(
        stateFF_inputPar[23]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_6_s_next_state[3]) );
  INV_X1 stateFF_state_gff_7_s_current_state_reg_3__U1 ( .A(data_out[27]), 
        .ZN(stateFF_state_gff_7_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_7_s_next_state[3]), .CK(clk), .Q(data_out[27]), 
        .QN() );
  INV_X1 stateFF_state_gff_7_s_current_state_reg_2__U1 ( .A(data_out[26]), 
        .ZN(stateFF_state_gff_7_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_7_s_next_state[2]), .CK(clk), .Q(data_out[26]), 
        .QN() );
  INV_X1 stateFF_state_gff_7_s_current_state_reg_1__U1 ( .A(data_out[25]), 
        .ZN(stateFF_state_gff_7_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_7_s_next_state[1]), .CK(clk), .Q(data_out[25]), 
        .QN() );
  INV_X1 stateFF_state_gff_7_s_current_state_reg_0__U1 ( .A(data_out[24]), 
        .ZN(stateFF_state_gff_7_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_7_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_7_s_next_state[0]), .CK(clk), .Q(data_out[24]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1 ( .A(data_out[20]), .B(
        stateFF_inputPar[24]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_7_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1 ( .A(data_out[21]), .B(
        stateFF_inputPar[25]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_7_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1 ( .A(data_out[22]), .B(
        stateFF_inputPar[26]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_7_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1 ( .A(data_out[23]), .B(
        stateFF_inputPar[27]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_7_s_next_state[3]) );
  INV_X1 stateFF_state_gff_8_s_current_state_reg_3__U1 ( .A(data_out[31]), 
        .ZN(stateFF_state_gff_8_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_8_s_next_state[3]), .CK(clk), .Q(data_out[31]), 
        .QN() );
  INV_X1 stateFF_state_gff_8_s_current_state_reg_2__U1 ( .A(data_out[30]), 
        .ZN(stateFF_state_gff_8_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_8_s_next_state[2]), .CK(clk), .Q(data_out[30]), 
        .QN() );
  INV_X1 stateFF_state_gff_8_s_current_state_reg_1__U1 ( .A(data_out[29]), 
        .ZN(stateFF_state_gff_8_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_8_s_next_state[1]), .CK(clk), .Q(data_out[29]), 
        .QN() );
  INV_X1 stateFF_state_gff_8_s_current_state_reg_0__U1 ( .A(data_out[28]), 
        .ZN(stateFF_state_gff_8_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_8_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_8_s_next_state[0]), .CK(clk), .Q(data_out[28]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1 ( .A(data_out[24]), .B(
        stateFF_inputPar[28]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_8_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1 ( .A(data_out[25]), .B(
        stateFF_inputPar[29]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_8_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1 ( .A(data_out[26]), .B(
        stateFF_inputPar[30]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_8_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1 ( .A(data_out[27]), .B(
        stateFF_inputPar[31]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_8_s_next_state[3]) );
  INV_X1 stateFF_state_gff_9_s_current_state_reg_3__U1 ( .A(data_out[35]), 
        .ZN(stateFF_state_gff_9_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_9_s_next_state[3]), .CK(clk), .Q(data_out[35]), 
        .QN() );
  INV_X1 stateFF_state_gff_9_s_current_state_reg_2__U1 ( .A(data_out[34]), 
        .ZN(stateFF_state_gff_9_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_9_s_next_state[2]), .CK(clk), .Q(data_out[34]), 
        .QN() );
  INV_X1 stateFF_state_gff_9_s_current_state_reg_1__U1 ( .A(data_out[33]), 
        .ZN(stateFF_state_gff_9_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_9_s_next_state[1]), .CK(clk), .Q(data_out[33]), 
        .QN() );
  INV_X1 stateFF_state_gff_9_s_current_state_reg_0__U1 ( .A(data_out[32]), 
        .ZN(stateFF_state_gff_9_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_9_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_9_s_next_state[0]), .CK(clk), .Q(data_out[32]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1 ( .A(data_out[28]), .B(
        stateFF_inputPar[32]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_9_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1 ( .A(data_out[29]), .B(
        stateFF_inputPar[33]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_9_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1 ( .A(data_out[30]), .B(
        stateFF_inputPar[34]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_9_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1 ( .A(data_out[31]), .B(
        stateFF_inputPar[35]), .S(stateFF_state_n6), .Z(
        stateFF_state_gff_9_s_next_state[3]) );
  INV_X1 stateFF_state_gff_10_s_current_state_reg_3__U1 ( .A(data_out[39]), 
        .ZN(stateFF_state_gff_10_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_10_s_next_state[3]), .CK(clk), .Q(data_out[39]), 
        .QN() );
  INV_X1 stateFF_state_gff_10_s_current_state_reg_2__U1 ( .A(data_out[38]), 
        .ZN(stateFF_state_gff_10_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_10_s_next_state[2]), .CK(clk), .Q(data_out[38]), 
        .QN() );
  INV_X1 stateFF_state_gff_10_s_current_state_reg_1__U1 ( .A(data_out[37]), 
        .ZN(stateFF_state_gff_10_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_10_s_next_state[1]), .CK(clk), .Q(data_out[37]), 
        .QN() );
  INV_X1 stateFF_state_gff_10_s_current_state_reg_0__U1 ( .A(data_out[36]), 
        .ZN(stateFF_state_gff_10_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_10_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_10_s_next_state[0]), .CK(clk), .Q(data_out[36]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1 ( .A(data_out[32]), .B(
        stateFF_inputPar[36]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_10_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1 ( .A(data_out[33]), .B(
        stateFF_inputPar[37]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_10_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1 ( .A(data_out[34]), .B(
        stateFF_inputPar[38]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_10_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1 ( .A(data_out[35]), .B(
        stateFF_inputPar[39]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_10_s_next_state[3]) );
  INV_X1 stateFF_state_gff_11_s_current_state_reg_3__U1 ( .A(data_out[43]), 
        .ZN(stateFF_state_gff_11_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_11_s_next_state[3]), .CK(clk), .Q(data_out[43]), 
        .QN() );
  INV_X1 stateFF_state_gff_11_s_current_state_reg_2__U1 ( .A(data_out[42]), 
        .ZN(stateFF_state_gff_11_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_11_s_next_state[2]), .CK(clk), .Q(data_out[42]), 
        .QN() );
  INV_X1 stateFF_state_gff_11_s_current_state_reg_1__U1 ( .A(data_out[41]), 
        .ZN(stateFF_state_gff_11_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_11_s_next_state[1]), .CK(clk), .Q(data_out[41]), 
        .QN() );
  INV_X1 stateFF_state_gff_11_s_current_state_reg_0__U1 ( .A(data_out[40]), 
        .ZN(stateFF_state_gff_11_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_11_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_11_s_next_state[0]), .CK(clk), .Q(data_out[40]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1 ( .A(data_out[36]), .B(
        stateFF_inputPar[40]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_11_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1 ( .A(data_out[37]), .B(
        stateFF_inputPar[41]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_11_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1 ( .A(data_out[38]), .B(
        stateFF_inputPar[42]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_11_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1 ( .A(data_out[39]), .B(
        stateFF_inputPar[43]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_11_s_next_state[3]) );
  INV_X1 stateFF_state_gff_12_s_current_state_reg_3__U1 ( .A(data_out[47]), 
        .ZN(stateFF_state_gff_12_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_12_s_next_state[3]), .CK(clk), .Q(data_out[47]), 
        .QN() );
  INV_X1 stateFF_state_gff_12_s_current_state_reg_2__U1 ( .A(data_out[46]), 
        .ZN(stateFF_state_gff_12_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_12_s_next_state[2]), .CK(clk), .Q(data_out[46]), 
        .QN() );
  INV_X1 stateFF_state_gff_12_s_current_state_reg_1__U1 ( .A(data_out[45]), 
        .ZN(stateFF_state_gff_12_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_12_s_next_state[1]), .CK(clk), .Q(data_out[45]), 
        .QN() );
  INV_X1 stateFF_state_gff_12_s_current_state_reg_0__U1 ( .A(data_out[44]), 
        .ZN(stateFF_state_gff_12_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_12_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_12_s_next_state[0]), .CK(clk), .Q(data_out[44]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1 ( .A(data_out[40]), .B(
        stateFF_inputPar[44]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_12_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1 ( .A(data_out[41]), .B(
        stateFF_inputPar[45]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_12_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1 ( .A(data_out[42]), .B(
        stateFF_inputPar[46]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_12_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1 ( .A(data_out[43]), .B(
        stateFF_inputPar[47]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_12_s_next_state[3]) );
  INV_X1 stateFF_state_gff_13_s_current_state_reg_3__U1 ( .A(data_out[51]), 
        .ZN(stateFF_state_gff_13_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_13_s_next_state[3]), .CK(clk), .Q(data_out[51]), 
        .QN() );
  INV_X1 stateFF_state_gff_13_s_current_state_reg_2__U1 ( .A(data_out[50]), 
        .ZN(stateFF_state_gff_13_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_13_s_next_state[2]), .CK(clk), .Q(data_out[50]), 
        .QN() );
  INV_X1 stateFF_state_gff_13_s_current_state_reg_1__U1 ( .A(data_out[49]), 
        .ZN(stateFF_state_gff_13_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_13_s_next_state[1]), .CK(clk), .Q(data_out[49]), 
        .QN() );
  INV_X1 stateFF_state_gff_13_s_current_state_reg_0__U1 ( .A(data_out[48]), 
        .ZN(stateFF_state_gff_13_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_13_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_13_s_next_state[0]), .CK(clk), .Q(data_out[48]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1 ( .A(data_out[44]), .B(
        stateFF_inputPar[48]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_13_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1 ( .A(data_out[45]), .B(
        stateFF_inputPar[49]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_13_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1 ( .A(data_out[46]), .B(
        stateFF_inputPar[50]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_13_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1 ( .A(data_out[47]), .B(
        stateFF_inputPar[51]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_13_s_next_state[3]) );
  INV_X1 stateFF_state_gff_14_s_current_state_reg_3__U1 ( .A(data_out[55]), 
        .ZN(stateFF_state_gff_14_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_14_s_next_state[3]), .CK(clk), .Q(data_out[55]), 
        .QN() );
  INV_X1 stateFF_state_gff_14_s_current_state_reg_2__U1 ( .A(data_out[54]), 
        .ZN(stateFF_state_gff_14_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_14_s_next_state[2]), .CK(clk), .Q(data_out[54]), 
        .QN() );
  INV_X1 stateFF_state_gff_14_s_current_state_reg_1__U1 ( .A(data_out[53]), 
        .ZN(stateFF_state_gff_14_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_14_s_next_state[1]), .CK(clk), .Q(data_out[53]), 
        .QN() );
  INV_X1 stateFF_state_gff_14_s_current_state_reg_0__U1 ( .A(data_out[52]), 
        .ZN(stateFF_state_gff_14_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_14_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_14_s_next_state[0]), .CK(clk), .Q(data_out[52]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1 ( .A(data_out[48]), .B(
        stateFF_inputPar[52]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_14_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1 ( .A(data_out[49]), .B(
        stateFF_inputPar[53]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_14_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1 ( .A(data_out[50]), .B(
        stateFF_inputPar[54]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_14_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1 ( .A(data_out[51]), .B(
        stateFF_inputPar[55]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_14_s_next_state[3]) );
  INV_X1 stateFF_state_gff_15_s_current_state_reg_3__U1 ( .A(data_out[59]), 
        .ZN(stateFF_state_gff_15_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_15_s_next_state[3]), .CK(clk), .Q(data_out[59]), 
        .QN() );
  INV_X1 stateFF_state_gff_15_s_current_state_reg_2__U1 ( .A(data_out[58]), 
        .ZN(stateFF_state_gff_15_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_15_s_next_state[2]), .CK(clk), .Q(data_out[58]), 
        .QN() );
  INV_X1 stateFF_state_gff_15_s_current_state_reg_1__U1 ( .A(data_out[57]), 
        .ZN(stateFF_state_gff_15_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_15_s_next_state[1]), .CK(clk), .Q(data_out[57]), 
        .QN() );
  INV_X1 stateFF_state_gff_15_s_current_state_reg_0__U1 ( .A(data_out[56]), 
        .ZN(stateFF_state_gff_15_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_15_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_15_s_next_state[0]), .CK(clk), .Q(data_out[56]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1 ( .A(data_out[52]), .B(
        stateFF_inputPar[56]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_15_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1 ( .A(data_out[53]), .B(
        stateFF_inputPar[57]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_15_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1 ( .A(data_out[54]), .B(
        stateFF_inputPar[58]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_15_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1 ( .A(data_out[55]), .B(
        stateFF_inputPar[59]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_15_s_next_state[3]) );
  INV_X1 stateFF_state_gff_16_s_current_state_reg_3__U1 ( .A(data_out[63]), 
        .ZN(stateFF_state_gff_16_s_current_state_reg_3__QN) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_3__FF_FF ( .D(
        stateFF_state_gff_16_s_next_state[3]), .CK(clk), .Q(data_out[63]), 
        .QN() );
  INV_X1 stateFF_state_gff_16_s_current_state_reg_2__U1 ( .A(data_out[62]), 
        .ZN(stateFF_state_gff_16_s_current_state_reg_2__QN) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_2__FF_FF ( .D(
        stateFF_state_gff_16_s_next_state[2]), .CK(clk), .Q(data_out[62]), 
        .QN() );
  INV_X1 stateFF_state_gff_16_s_current_state_reg_1__U1 ( .A(data_out[61]), 
        .ZN(stateFF_state_gff_16_s_current_state_reg_1__QN) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_1__FF_FF ( .D(
        stateFF_state_gff_16_s_next_state[1]), .CK(clk), .Q(data_out[61]), 
        .QN() );
  INV_X1 stateFF_state_gff_16_s_current_state_reg_0__U1 ( .A(data_out[60]), 
        .ZN(stateFF_state_gff_16_s_current_state_reg_0__QN) );
  DFF_X1 stateFF_state_gff_16_s_current_state_reg_0__FF_FF ( .D(
        stateFF_state_gff_16_s_next_state[0]), .CK(clk), .Q(data_out[60]), 
        .QN() );
  MUX2_X1 stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1 ( .A(data_out[56]), .B(
        stateFF_inputPar[60]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_16_s_next_state[0]) );
  MUX2_X1 stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1 ( .A(data_out[57]), .B(
        stateFF_inputPar[61]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_16_s_next_state[1]) );
  MUX2_X1 stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1 ( .A(data_out[58]), .B(
        stateFF_inputPar[62]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_16_s_next_state[2]) );
  MUX2_X1 stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1 ( .A(data_out[59]), .B(
        stateFF_inputPar[63]), .S(stateFF_state_n5), .Z(
        stateFF_state_gff_16_s_next_state[3]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_0_U1 ( .A(data_out[0]), .B(data_in[0]), 
        .S(reset), .Z(stateFF_inputPar[0]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_1_U1 ( .A(data_out[4]), .B(data_in[1]), 
        .S(reset), .Z(stateFF_inputPar[1]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_2_U1 ( .A(data_out[8]), .B(data_in[2]), 
        .S(reset), .Z(stateFF_inputPar[2]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_3_U1 ( .A(data_out[12]), .B(data_in[3]), .S(reset), .Z(stateFF_inputPar[3]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_4_U1 ( .A(data_out[16]), .B(data_in[4]), .S(reset), .Z(stateFF_inputPar[4]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_5_U1 ( .A(data_out[20]), .B(data_in[5]), .S(reset), .Z(stateFF_inputPar[5]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_6_U1 ( .A(data_out[24]), .B(data_in[6]), .S(reset), .Z(stateFF_inputPar[6]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_7_U1 ( .A(data_out[28]), .B(data_in[7]), .S(reset), .Z(stateFF_inputPar[7]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_8_U1 ( .A(data_out[32]), .B(data_in[8]), .S(reset), .Z(stateFF_inputPar[8]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_9_U1 ( .A(data_out[36]), .B(data_in[9]), .S(reset), .Z(stateFF_inputPar[9]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_10_U1 ( .A(data_out[40]), .B(
        data_in[10]), .S(reset), .Z(stateFF_inputPar[10]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_11_U1 ( .A(data_out[44]), .B(
        data_in[11]), .S(reset), .Z(stateFF_inputPar[11]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_12_U1 ( .A(data_out[48]), .B(
        data_in[12]), .S(reset), .Z(stateFF_inputPar[12]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_13_U1 ( .A(data_out[52]), .B(
        data_in[13]), .S(reset), .Z(stateFF_inputPar[13]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_14_U1 ( .A(data_out[56]), .B(
        data_in[14]), .S(reset), .Z(stateFF_inputPar[14]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_15_U1 ( .A(data_out[60]), .B(
        data_in[15]), .S(reset), .Z(stateFF_inputPar[15]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_16_U1 ( .A(data_out[1]), .B(
        data_in[16]), .S(reset), .Z(stateFF_inputPar[16]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_17_U1 ( .A(data_out[5]), .B(
        data_in[17]), .S(reset), .Z(stateFF_inputPar[17]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_18_U1 ( .A(data_out[9]), .B(
        data_in[18]), .S(reset), .Z(stateFF_inputPar[18]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_19_U1 ( .A(data_out[13]), .B(
        data_in[19]), .S(reset), .Z(stateFF_inputPar[19]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_20_U1 ( .A(data_out[17]), .B(
        data_in[20]), .S(reset), .Z(stateFF_inputPar[20]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_21_U1 ( .A(data_out[21]), .B(
        data_in[21]), .S(reset), .Z(stateFF_inputPar[21]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_22_U1 ( .A(data_out[25]), .B(
        data_in[22]), .S(reset), .Z(stateFF_inputPar[22]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_23_U1 ( .A(data_out[29]), .B(
        data_in[23]), .S(reset), .Z(stateFF_inputPar[23]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_24_U1 ( .A(data_out[33]), .B(
        data_in[24]), .S(reset), .Z(stateFF_inputPar[24]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_25_U1 ( .A(data_out[37]), .B(
        data_in[25]), .S(reset), .Z(stateFF_inputPar[25]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_26_U1 ( .A(data_out[41]), .B(
        data_in[26]), .S(reset), .Z(stateFF_inputPar[26]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_27_U1 ( .A(data_out[45]), .B(
        data_in[27]), .S(reset), .Z(stateFF_inputPar[27]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_28_U1 ( .A(data_out[49]), .B(
        data_in[28]), .S(reset), .Z(stateFF_inputPar[28]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_29_U1 ( .A(data_out[53]), .B(
        data_in[29]), .S(reset), .Z(stateFF_inputPar[29]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_30_U1 ( .A(data_out[57]), .B(
        data_in[30]), .S(reset), .Z(stateFF_inputPar[30]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_31_U1 ( .A(data_out[61]), .B(
        data_in[31]), .S(reset), .Z(stateFF_inputPar[31]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_32_U1 ( .A(data_out[2]), .B(
        data_in[32]), .S(reset), .Z(stateFF_inputPar[32]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_33_U1 ( .A(data_out[6]), .B(
        data_in[33]), .S(reset), .Z(stateFF_inputPar[33]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_34_U1 ( .A(data_out[10]), .B(
        data_in[34]), .S(reset), .Z(stateFF_inputPar[34]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_35_U1 ( .A(data_out[14]), .B(
        data_in[35]), .S(reset), .Z(stateFF_inputPar[35]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_36_U1 ( .A(data_out[18]), .B(
        data_in[36]), .S(reset), .Z(stateFF_inputPar[36]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_37_U1 ( .A(data_out[22]), .B(
        data_in[37]), .S(reset), .Z(stateFF_inputPar[37]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_38_U1 ( .A(data_out[26]), .B(
        data_in[38]), .S(reset), .Z(stateFF_inputPar[38]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_39_U1 ( .A(data_out[30]), .B(
        data_in[39]), .S(reset), .Z(stateFF_inputPar[39]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_40_U1 ( .A(data_out[34]), .B(
        data_in[40]), .S(reset), .Z(stateFF_inputPar[40]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_41_U1 ( .A(data_out[38]), .B(
        data_in[41]), .S(reset), .Z(stateFF_inputPar[41]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_42_U1 ( .A(data_out[42]), .B(
        data_in[42]), .S(reset), .Z(stateFF_inputPar[42]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_43_U1 ( .A(data_out[46]), .B(
        data_in[43]), .S(reset), .Z(stateFF_inputPar[43]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_44_U1 ( .A(data_out[50]), .B(
        data_in[44]), .S(reset), .Z(stateFF_inputPar[44]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_45_U1 ( .A(data_out[54]), .B(
        data_in[45]), .S(reset), .Z(stateFF_inputPar[45]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_46_U1 ( .A(data_out[58]), .B(
        data_in[46]), .S(reset), .Z(stateFF_inputPar[46]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_47_U1 ( .A(data_out[62]), .B(
        data_in[47]), .S(reset), .Z(stateFF_inputPar[47]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_48_U1 ( .A(data_out[3]), .B(
        data_in[48]), .S(reset), .Z(stateFF_inputPar[48]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_49_U1 ( .A(data_out[7]), .B(
        data_in[49]), .S(reset), .Z(stateFF_inputPar[49]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_50_U1 ( .A(data_out[11]), .B(
        data_in[50]), .S(reset), .Z(stateFF_inputPar[50]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_51_U1 ( .A(data_out[15]), .B(
        data_in[51]), .S(reset), .Z(stateFF_inputPar[51]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_52_U1 ( .A(data_out[19]), .B(
        data_in[52]), .S(reset), .Z(stateFF_inputPar[52]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_53_U1 ( .A(data_out[23]), .B(
        data_in[53]), .S(reset), .Z(stateFF_inputPar[53]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_54_U1 ( .A(data_out[27]), .B(
        data_in[54]), .S(reset), .Z(stateFF_inputPar[54]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_55_U1 ( .A(data_out[31]), .B(
        data_in[55]), .S(reset), .Z(stateFF_inputPar[55]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_56_U1 ( .A(data_out[35]), .B(
        data_in[56]), .S(reset), .Z(stateFF_inputPar[56]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_57_U1 ( .A(data_out[39]), .B(
        data_in[57]), .S(reset), .Z(stateFF_inputPar[57]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_58_U1 ( .A(data_out[43]), .B(
        data_in[58]), .S(reset), .Z(stateFF_inputPar[58]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_59_U1 ( .A(data_out[47]), .B(
        data_in[59]), .S(reset), .Z(stateFF_inputPar[59]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_60_U1 ( .A(data_out[51]), .B(
        data_in[60]), .S(reset), .Z(stateFF_inputPar[60]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_61_U1 ( .A(data_out[55]), .B(
        data_in[61]), .S(reset), .Z(stateFF_inputPar[61]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_62_U1 ( .A(data_out[59]), .B(
        data_in[62]), .S(reset), .Z(stateFF_inputPar[62]) );
  MUX2_X1 stateFF_MUX_inputPar_mux_inst_63_U1 ( .A(data_out[63]), .B(
        data_in[63]), .S(reset), .Z(stateFF_inputPar[63]) );
  XOR2_X1 keyFF_U5 ( .A(counter[4]), .B(keyFF_outputPar[22]), .Z(
        keyFF_counterAdd[4]) );
  XOR2_X1 keyFF_U4 ( .A(counter[3]), .B(keyFF_outputPar[21]), .Z(
        keyFF_counterAdd[3]) );
  XOR2_X1 keyFF_U3 ( .A(counter[2]), .B(keyFF_outputPar[20]), .Z(
        keyFF_counterAdd[2]) );
  XOR2_X1 keyFF_U2 ( .A(counter[1]), .B(keyFF_outputPar[19]), .Z(
        keyFF_counterAdd[1]) );
  XOR2_X1 keyFF_U1 ( .A(counter[0]), .B(keyFF_outputPar[18]), .Z(
        keyFF_counterAdd[0]) );
  INV_X2 keyFF_keystate_U3 ( .A(keyFF_keystate_n8), .ZN(keyFF_keystate_n6) );
  INV_X2 keyFF_keystate_U2 ( .A(keyFF_keystate_n8), .ZN(keyFF_keystate_n7) );
  INV_X1 keyFF_keystate_U1 ( .A(ctrlData_0_), .ZN(keyFF_keystate_n8) );
  INV_X1 keyFF_keystate_gff_1_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[3]), .ZN(
        keyFF_keystate_gff_1_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_1_s_next_state[3]), .CK(clk), .Q(keyFF_outputPar[3]), .QN() );
  INV_X1 keyFF_keystate_gff_1_s_current_state_reg_2__U1 ( .A(keyRegKS[3]), 
        .ZN(keyFF_keystate_gff_1_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_1_s_next_state[2]), .CK(clk), .Q(keyRegKS[3]), 
        .QN() );
  INV_X1 keyFF_keystate_gff_1_s_current_state_reg_1__U1 ( .A(keyRegKS[2]), 
        .ZN(keyFF_keystate_gff_1_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_1_s_next_state[1]), .CK(clk), .Q(keyRegKS[2]), 
        .QN() );
  INV_X1 keyFF_keystate_gff_1_s_current_state_reg_0__U1 ( .A(keyRegKS[1]), 
        .ZN(keyFF_keystate_gff_1_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_1_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_1_s_next_state[0]), .CK(clk), .Q(keyRegKS[1]), 
        .QN() );
  MUX2_X1 keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1 ( .A(roundkey[0]), .B(
        keyFF_inputPar[0]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_1_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1 ( .A(roundkey[1]), .B(
        keyFF_inputPar[1]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_1_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1 ( .A(roundkey[2]), .B(
        keyFF_inputPar[2]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_1_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1 ( .A(roundkey[3]), .B(
        keyFF_inputPar[3]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_1_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_2_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[7]), .ZN(
        keyFF_keystate_gff_2_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_2_s_next_state[3]), .CK(clk), .Q(keyFF_outputPar[7]), .QN() );
  INV_X1 keyFF_keystate_gff_2_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[6]), .ZN(
        keyFF_keystate_gff_2_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_2_s_next_state[2]), .CK(clk), .Q(keyFF_outputPar[6]), .QN() );
  INV_X1 keyFF_keystate_gff_2_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[5]), .ZN(
        keyFF_keystate_gff_2_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_2_s_next_state[1]), .CK(clk), .Q(keyFF_outputPar[5]), .QN() );
  INV_X1 keyFF_keystate_gff_2_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[4]), .ZN(
        keyFF_keystate_gff_2_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_2_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_2_s_next_state[0]), .CK(clk), .Q(keyFF_outputPar[4]), .QN() );
  MUX2_X1 keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1 ( .A(keyRegKS[1]), .B(
        keyFF_inputPar[4]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_2_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1 ( .A(keyRegKS[2]), .B(
        keyFF_inputPar[5]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_2_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1 ( .A(keyRegKS[3]), .B(
        keyFF_inputPar[6]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_2_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1 ( .A(keyFF_outputPar[3]), .B(keyFF_inputPar[7]), .S(keyFF_keystate_n7), .Z(
        keyFF_keystate_gff_2_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_3_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[11]), .ZN(
        keyFF_keystate_gff_3_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_3_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[11]), .QN() );
  INV_X1 keyFF_keystate_gff_3_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[10]), .ZN(
        keyFF_keystate_gff_3_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_3_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[10]), .QN() );
  INV_X1 keyFF_keystate_gff_3_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[9]), .ZN(
        keyFF_keystate_gff_3_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_3_s_next_state[1]), .CK(clk), .Q(keyFF_outputPar[9]), .QN() );
  INV_X1 keyFF_keystate_gff_3_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[8]), .ZN(
        keyFF_keystate_gff_3_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_3_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_3_s_next_state[0]), .CK(clk), .Q(keyFF_outputPar[8]), .QN() );
  MUX2_X1 keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1 ( .A(keyFF_outputPar[4]), .B(keyFF_inputPar[8]), .S(keyFF_keystate_n6), .Z(
        keyFF_keystate_gff_3_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1 ( .A(keyFF_outputPar[5]), .B(keyFF_inputPar[9]), .S(keyFF_keystate_n6), .Z(
        keyFF_keystate_gff_3_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1 ( .A(keyFF_outputPar[6]), .B(keyFF_inputPar[10]), .S(keyFF_keystate_n6), .Z(
        keyFF_keystate_gff_3_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1 ( .A(keyFF_outputPar[7]), .B(keyFF_inputPar[11]), .S(keyFF_keystate_n6), .Z(
        keyFF_keystate_gff_3_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_4_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[15]), .ZN(
        keyFF_keystate_gff_4_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_4_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[15]), .QN() );
  INV_X1 keyFF_keystate_gff_4_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[14]), .ZN(
        keyFF_keystate_gff_4_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_4_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[14]), .QN() );
  INV_X1 keyFF_keystate_gff_4_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[13]), .ZN(
        keyFF_keystate_gff_4_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_4_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[13]), .QN() );
  INV_X1 keyFF_keystate_gff_4_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[12]), .ZN(
        keyFF_keystate_gff_4_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_4_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_4_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[12]), .QN() );
  MUX2_X1 keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1 ( .A(keyFF_outputPar[8]), .B(keyFF_inputPar[12]), .S(keyFF_keystate_n6), .Z(
        keyFF_keystate_gff_4_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1 ( .A(keyFF_outputPar[9]), .B(keyFF_inputPar[13]), .S(keyFF_keystate_n6), .Z(
        keyFF_keystate_gff_4_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[10]), .B(keyFF_inputPar[14]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_4_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[11]), .B(keyFF_inputPar[15]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_4_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_5_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[19]), .ZN(
        keyFF_keystate_gff_5_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_5_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[19]), .QN() );
  INV_X1 keyFF_keystate_gff_5_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[18]), .ZN(
        keyFF_keystate_gff_5_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_5_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[18]), .QN() );
  INV_X1 keyFF_keystate_gff_5_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[17]), .ZN(
        keyFF_keystate_gff_5_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_5_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[17]), .QN() );
  INV_X1 keyFF_keystate_gff_5_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[16]), .ZN(
        keyFF_keystate_gff_5_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_5_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_5_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[16]), .QN() );
  MUX2_X1 keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[12]), .B(keyFF_inputPar[16]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_5_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[13]), .B(keyFF_inputPar[17]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_5_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[14]), .B(keyFF_inputPar[18]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_5_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[15]), .B(keyFF_inputPar[19]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_5_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_6_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[23]), .ZN(
        keyFF_keystate_gff_6_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_6_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[23]), .QN() );
  INV_X1 keyFF_keystate_gff_6_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[22]), .ZN(
        keyFF_keystate_gff_6_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_6_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[22]), .QN() );
  INV_X1 keyFF_keystate_gff_6_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[21]), .ZN(
        keyFF_keystate_gff_6_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_6_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[21]), .QN() );
  INV_X1 keyFF_keystate_gff_6_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[20]), .ZN(
        keyFF_keystate_gff_6_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_6_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_6_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[20]), .QN() );
  MUX2_X1 keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[16]), .B(keyFF_inputPar[20]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_6_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[17]), .B(keyFF_inputPar[21]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_6_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[18]), .B(keyFF_inputPar[22]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_6_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[19]), .B(keyFF_inputPar[23]), .S(ctrlData_0_), .Z(
        keyFF_keystate_gff_6_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_7_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[27]), .ZN(
        keyFF_keystate_gff_7_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_7_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[27]), .QN() );
  INV_X1 keyFF_keystate_gff_7_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[26]), .ZN(
        keyFF_keystate_gff_7_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_7_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[26]), .QN() );
  INV_X1 keyFF_keystate_gff_7_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[25]), .ZN(
        keyFF_keystate_gff_7_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_7_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[25]), .QN() );
  INV_X1 keyFF_keystate_gff_7_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[24]), .ZN(
        keyFF_keystate_gff_7_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_7_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_7_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[24]), .QN() );
  MUX2_X1 keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[20]), .B(keyFF_inputPar[24]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_7_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[21]), .B(keyFF_inputPar[25]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_7_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[22]), .B(keyFF_inputPar[26]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_7_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[23]), .B(keyFF_inputPar[27]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_7_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_8_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[31]), .ZN(
        keyFF_keystate_gff_8_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_8_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[31]), .QN() );
  INV_X1 keyFF_keystate_gff_8_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[30]), .ZN(
        keyFF_keystate_gff_8_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_8_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[30]), .QN() );
  INV_X1 keyFF_keystate_gff_8_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[29]), .ZN(
        keyFF_keystate_gff_8_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_8_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[29]), .QN() );
  INV_X1 keyFF_keystate_gff_8_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[28]), .ZN(
        keyFF_keystate_gff_8_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_8_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_8_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[28]), .QN() );
  MUX2_X1 keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[24]), .B(keyFF_inputPar[28]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_8_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[25]), .B(keyFF_inputPar[29]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_8_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[26]), .B(keyFF_inputPar[30]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_8_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[27]), .B(keyFF_inputPar[31]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_8_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_9_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[35]), .ZN(
        keyFF_keystate_gff_9_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_9_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[35]), .QN() );
  INV_X1 keyFF_keystate_gff_9_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[34]), .ZN(
        keyFF_keystate_gff_9_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_9_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[34]), .QN() );
  INV_X1 keyFF_keystate_gff_9_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[33]), .ZN(
        keyFF_keystate_gff_9_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_9_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[33]), .QN() );
  INV_X1 keyFF_keystate_gff_9_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[32]), .ZN(
        keyFF_keystate_gff_9_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_9_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_9_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[32]), .QN() );
  MUX2_X1 keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[28]), .B(keyFF_inputPar[32]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_9_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[29]), .B(keyFF_inputPar[33]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_9_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[30]), .B(keyFF_inputPar[34]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_9_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[31]), .B(keyFF_inputPar[35]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_9_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_10_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[39]), .ZN(
        keyFF_keystate_gff_10_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_10_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[39]), .QN() );
  INV_X1 keyFF_keystate_gff_10_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[38]), .ZN(
        keyFF_keystate_gff_10_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_10_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[38]), .QN() );
  INV_X1 keyFF_keystate_gff_10_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[37]), .ZN(
        keyFF_keystate_gff_10_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_10_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[37]), .QN() );
  INV_X1 keyFF_keystate_gff_10_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[36]), .ZN(
        keyFF_keystate_gff_10_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_10_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_10_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[36]), .QN() );
  MUX2_X1 keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[32]), .B(keyFF_inputPar[36]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_10_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[33]), .B(keyFF_inputPar[37]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_10_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[34]), .B(keyFF_inputPar[38]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_10_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[35]), .B(keyFF_inputPar[39]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_10_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_11_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[43]), .ZN(
        keyFF_keystate_gff_11_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_11_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[43]), .QN() );
  INV_X1 keyFF_keystate_gff_11_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[42]), .ZN(
        keyFF_keystate_gff_11_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_11_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[42]), .QN() );
  INV_X1 keyFF_keystate_gff_11_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[41]), .ZN(
        keyFF_keystate_gff_11_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_11_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[41]), .QN() );
  INV_X1 keyFF_keystate_gff_11_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[40]), .ZN(
        keyFF_keystate_gff_11_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_11_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_11_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[40]), .QN() );
  MUX2_X1 keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[36]), .B(keyFF_inputPar[40]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_11_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[37]), .B(keyFF_inputPar[41]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_11_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[38]), .B(keyFF_inputPar[42]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_11_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[39]), .B(keyFF_inputPar[43]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_11_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_12_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[47]), .ZN(
        keyFF_keystate_gff_12_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_12_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[47]), .QN() );
  INV_X1 keyFF_keystate_gff_12_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[46]), .ZN(
        keyFF_keystate_gff_12_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_12_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[46]), .QN() );
  INV_X1 keyFF_keystate_gff_12_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[45]), .ZN(
        keyFF_keystate_gff_12_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_12_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[45]), .QN() );
  INV_X1 keyFF_keystate_gff_12_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[44]), .ZN(
        keyFF_keystate_gff_12_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_12_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_12_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[44]), .QN() );
  MUX2_X1 keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[40]), .B(keyFF_inputPar[44]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_12_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[41]), .B(keyFF_inputPar[45]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_12_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[42]), .B(keyFF_inputPar[46]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_12_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[43]), .B(keyFF_inputPar[47]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_12_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_13_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[51]), .ZN(
        keyFF_keystate_gff_13_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_13_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[51]), .QN() );
  INV_X1 keyFF_keystate_gff_13_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[50]), .ZN(
        keyFF_keystate_gff_13_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_13_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[50]), .QN() );
  INV_X1 keyFF_keystate_gff_13_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[49]), .ZN(
        keyFF_keystate_gff_13_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_13_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[49]), .QN() );
  INV_X1 keyFF_keystate_gff_13_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[48]), .ZN(
        keyFF_keystate_gff_13_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_13_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_13_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[48]), .QN() );
  MUX2_X1 keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[44]), .B(keyFF_inputPar[48]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_13_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[45]), .B(keyFF_inputPar[49]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_13_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[46]), .B(keyFF_inputPar[50]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_13_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[47]), .B(keyFF_inputPar[51]), .S(keyFF_keystate_n7), 
        .Z(keyFF_keystate_gff_13_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_14_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[55]), .ZN(
        keyFF_keystate_gff_14_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_14_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[55]), .QN() );
  INV_X1 keyFF_keystate_gff_14_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[54]), .ZN(
        keyFF_keystate_gff_14_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_14_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[54]), .QN() );
  INV_X1 keyFF_keystate_gff_14_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[53]), .ZN(
        keyFF_keystate_gff_14_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_14_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[53]), .QN() );
  INV_X1 keyFF_keystate_gff_14_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[52]), .ZN(
        keyFF_keystate_gff_14_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_14_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_14_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[52]), .QN() );
  MUX2_X1 keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[48]), .B(keyFF_inputPar[52]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_14_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[49]), .B(keyFF_inputPar[53]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_14_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[50]), .B(keyFF_inputPar[54]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_14_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[51]), .B(keyFF_inputPar[55]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_14_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_15_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[59]), .ZN(
        keyFF_keystate_gff_15_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_15_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[59]), .QN() );
  INV_X1 keyFF_keystate_gff_15_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[58]), .ZN(
        keyFF_keystate_gff_15_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_15_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[58]), .QN() );
  INV_X1 keyFF_keystate_gff_15_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[57]), .ZN(
        keyFF_keystate_gff_15_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_15_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[57]), .QN() );
  INV_X1 keyFF_keystate_gff_15_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[56]), .ZN(
        keyFF_keystate_gff_15_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_15_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_15_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[56]), .QN() );
  MUX2_X1 keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[52]), .B(keyFF_inputPar[56]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_15_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[53]), .B(keyFF_inputPar[57]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_15_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[54]), .B(keyFF_inputPar[58]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_15_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[55]), .B(keyFF_inputPar[59]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_15_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_16_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[63]), .ZN(
        keyFF_keystate_gff_16_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_16_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[63]), .QN() );
  INV_X1 keyFF_keystate_gff_16_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[62]), .ZN(
        keyFF_keystate_gff_16_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_16_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[62]), .QN() );
  INV_X1 keyFF_keystate_gff_16_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[61]), .ZN(
        keyFF_keystate_gff_16_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_16_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[61]), .QN() );
  INV_X1 keyFF_keystate_gff_16_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[60]), .ZN(
        keyFF_keystate_gff_16_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_16_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_16_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[60]), .QN() );
  MUX2_X1 keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[56]), .B(keyFF_inputPar[60]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_16_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[57]), .B(keyFF_inputPar[61]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_16_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[58]), .B(keyFF_inputPar[62]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_16_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[59]), .B(keyFF_inputPar[63]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_16_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_17_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[67]), .ZN(
        keyFF_keystate_gff_17_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_17_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[67]), .QN() );
  INV_X1 keyFF_keystate_gff_17_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[66]), .ZN(
        keyFF_keystate_gff_17_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_17_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[66]), .QN() );
  INV_X1 keyFF_keystate_gff_17_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[65]), .ZN(
        keyFF_keystate_gff_17_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_17_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[65]), .QN() );
  INV_X1 keyFF_keystate_gff_17_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[64]), .ZN(
        keyFF_keystate_gff_17_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_17_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_17_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[64]), .QN() );
  MUX2_X1 keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[60]), .B(keyFF_inputPar[64]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_17_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[61]), .B(keyFF_inputPar[65]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_17_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[62]), .B(keyFF_inputPar[66]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_17_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[63]), .B(keyFF_inputPar[67]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_17_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_18_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[71]), .ZN(
        keyFF_keystate_gff_18_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_18_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[71]), .QN() );
  INV_X1 keyFF_keystate_gff_18_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[70]), .ZN(
        keyFF_keystate_gff_18_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_18_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[70]), .QN() );
  INV_X1 keyFF_keystate_gff_18_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[69]), .ZN(
        keyFF_keystate_gff_18_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_18_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[69]), .QN() );
  INV_X1 keyFF_keystate_gff_18_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[68]), .ZN(
        keyFF_keystate_gff_18_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_18_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_18_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[68]), .QN() );
  MUX2_X1 keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[64]), .B(keyFF_inputPar[68]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_18_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[65]), .B(keyFF_inputPar[69]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_18_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[66]), .B(keyFF_inputPar[70]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_18_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[67]), .B(keyFF_inputPar[71]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_18_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_19_s_current_state_reg_3__U1 ( .A(
        keyFF_outputPar[75]), .ZN(
        keyFF_keystate_gff_19_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_19_s_next_state[3]), .CK(clk), .Q(
        keyFF_outputPar[75]), .QN() );
  INV_X1 keyFF_keystate_gff_19_s_current_state_reg_2__U1 ( .A(
        keyFF_outputPar[74]), .ZN(
        keyFF_keystate_gff_19_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_19_s_next_state[2]), .CK(clk), .Q(
        keyFF_outputPar[74]), .QN() );
  INV_X1 keyFF_keystate_gff_19_s_current_state_reg_1__U1 ( .A(
        keyFF_outputPar[73]), .ZN(
        keyFF_keystate_gff_19_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_19_s_next_state[1]), .CK(clk), .Q(
        keyFF_outputPar[73]), .QN() );
  INV_X1 keyFF_keystate_gff_19_s_current_state_reg_0__U1 ( .A(
        keyFF_outputPar[72]), .ZN(
        keyFF_keystate_gff_19_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_19_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_19_s_next_state[0]), .CK(clk), .Q(
        keyFF_outputPar[72]), .QN() );
  MUX2_X1 keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[68]), .B(keyFF_inputPar[72]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_19_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[69]), .B(keyFF_inputPar[73]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_19_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[70]), .B(keyFF_inputPar[74]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_19_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[71]), .B(keyFF_inputPar[75]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_19_s_next_state[3]) );
  INV_X1 keyFF_keystate_gff_20_s_current_state_reg_3__U1 ( .A(roundkey[3]), 
        .ZN(keyFF_keystate_gff_20_s_current_state_reg_3__QN) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_3__FF_FF ( .D(
        keyFF_keystate_gff_20_s_next_state[3]), .CK(clk), .Q(roundkey[3]), 
        .QN() );
  INV_X1 keyFF_keystate_gff_20_s_current_state_reg_2__U1 ( .A(roundkey[2]), 
        .ZN(keyFF_keystate_gff_20_s_current_state_reg_2__QN) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_2__FF_FF ( .D(
        keyFF_keystate_gff_20_s_next_state[2]), .CK(clk), .Q(roundkey[2]), 
        .QN() );
  INV_X1 keyFF_keystate_gff_20_s_current_state_reg_1__U1 ( .A(roundkey[1]), 
        .ZN(keyFF_keystate_gff_20_s_current_state_reg_1__QN) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_1__FF_FF ( .D(
        keyFF_keystate_gff_20_s_next_state[1]), .CK(clk), .Q(roundkey[1]), 
        .QN() );
  INV_X1 keyFF_keystate_gff_20_s_current_state_reg_0__U1 ( .A(roundkey[0]), 
        .ZN(keyFF_keystate_gff_20_s_current_state_reg_0__QN) );
  DFF_X1 keyFF_keystate_gff_20_s_current_state_reg_0__FF_FF ( .D(
        keyFF_keystate_gff_20_s_next_state[0]), .CK(clk), .Q(roundkey[0]), 
        .QN() );
  MUX2_X1 keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1 ( .A(
        keyFF_outputPar[72]), .B(keyFF_inputPar[76]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_20_s_next_state[0]) );
  MUX2_X1 keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1 ( .A(
        keyFF_outputPar[73]), .B(keyFF_inputPar[77]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_20_s_next_state[1]) );
  MUX2_X1 keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1 ( .A(
        keyFF_outputPar[74]), .B(keyFF_inputPar[78]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_20_s_next_state[2]) );
  MUX2_X1 keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1 ( .A(
        keyFF_outputPar[75]), .B(keyFF_inputPar[79]), .S(keyFF_keystate_n6), 
        .Z(keyFF_keystate_gff_20_s_next_state[3]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_0_U1 ( .A(keyFF_outputPar[3]), .B(key[0]), .S(reset), .Z(keyFF_inputPar[0]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_1_U1 ( .A(keyFF_outputPar[4]), .B(key[1]), .S(reset), .Z(keyFF_inputPar[1]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_2_U1 ( .A(keyFF_outputPar[5]), .B(key[2]), .S(reset), .Z(keyFF_inputPar[2]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_3_U1 ( .A(keyFF_outputPar[6]), .B(key[3]), .S(reset), .Z(keyFF_inputPar[3]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_4_U1 ( .A(keyFF_outputPar[7]), .B(key[4]), .S(reset), .Z(keyFF_inputPar[4]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_5_U1 ( .A(keyFF_outputPar[8]), .B(key[5]), .S(reset), .Z(keyFF_inputPar[5]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_6_U1 ( .A(keyFF_outputPar[9]), .B(key[6]), .S(reset), .Z(keyFF_inputPar[6]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_7_U1 ( .A(keyFF_outputPar[10]), .B(
        key[7]), .S(reset), .Z(keyFF_inputPar[7]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_8_U1 ( .A(keyFF_outputPar[11]), .B(
        key[8]), .S(reset), .Z(keyFF_inputPar[8]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_9_U1 ( .A(keyFF_outputPar[12]), .B(
        key[9]), .S(reset), .Z(keyFF_inputPar[9]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_10_U1 ( .A(keyFF_outputPar[13]), .B(
        key[10]), .S(reset), .Z(keyFF_inputPar[10]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_11_U1 ( .A(keyFF_outputPar[14]), .B(
        key[11]), .S(reset), .Z(keyFF_inputPar[11]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_12_U1 ( .A(keyFF_outputPar[15]), .B(
        key[12]), .S(reset), .Z(keyFF_inputPar[12]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_13_U1 ( .A(keyFF_outputPar[16]), .B(
        key[13]), .S(reset), .Z(keyFF_inputPar[13]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_14_U1 ( .A(keyFF_outputPar[17]), .B(
        key[14]), .S(reset), .Z(keyFF_inputPar[14]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_15_U1 ( .A(keyFF_counterAdd[0]), .B(
        key[15]), .S(reset), .Z(keyFF_inputPar[15]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_16_U1 ( .A(keyFF_counterAdd[1]), .B(
        key[16]), .S(reset), .Z(keyFF_inputPar[16]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_17_U1 ( .A(keyFF_counterAdd[2]), .B(
        key[17]), .S(reset), .Z(keyFF_inputPar[17]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_18_U1 ( .A(keyFF_counterAdd[3]), .B(
        key[18]), .S(reset), .Z(keyFF_inputPar[18]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_19_U1 ( .A(keyFF_counterAdd[4]), .B(
        key[19]), .S(reset), .Z(keyFF_inputPar[19]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_20_U1 ( .A(keyFF_outputPar[23]), .B(
        key[20]), .S(reset), .Z(keyFF_inputPar[20]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_21_U1 ( .A(keyFF_outputPar[24]), .B(
        key[21]), .S(reset), .Z(keyFF_inputPar[21]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_22_U1 ( .A(keyFF_outputPar[25]), .B(
        key[22]), .S(reset), .Z(keyFF_inputPar[22]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_23_U1 ( .A(keyFF_outputPar[26]), .B(
        key[23]), .S(reset), .Z(keyFF_inputPar[23]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_24_U1 ( .A(keyFF_outputPar[27]), .B(
        key[24]), .S(reset), .Z(keyFF_inputPar[24]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_25_U1 ( .A(keyFF_outputPar[28]), .B(
        key[25]), .S(reset), .Z(keyFF_inputPar[25]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_26_U1 ( .A(keyFF_outputPar[29]), .B(
        key[26]), .S(reset), .Z(keyFF_inputPar[26]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_27_U1 ( .A(keyFF_outputPar[30]), .B(
        key[27]), .S(reset), .Z(keyFF_inputPar[27]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_28_U1 ( .A(keyFF_outputPar[31]), .B(
        key[28]), .S(reset), .Z(keyFF_inputPar[28]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_29_U1 ( .A(keyFF_outputPar[32]), .B(
        key[29]), .S(reset), .Z(keyFF_inputPar[29]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_30_U1 ( .A(keyFF_outputPar[33]), .B(
        key[30]), .S(reset), .Z(keyFF_inputPar[30]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_31_U1 ( .A(keyFF_outputPar[34]), .B(
        key[31]), .S(reset), .Z(keyFF_inputPar[31]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_32_U1 ( .A(keyFF_outputPar[35]), .B(
        key[32]), .S(reset), .Z(keyFF_inputPar[32]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_33_U1 ( .A(keyFF_outputPar[36]), .B(
        key[33]), .S(reset), .Z(keyFF_inputPar[33]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_34_U1 ( .A(keyFF_outputPar[37]), .B(
        key[34]), .S(reset), .Z(keyFF_inputPar[34]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_35_U1 ( .A(keyFF_outputPar[38]), .B(
        key[35]), .S(reset), .Z(keyFF_inputPar[35]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_36_U1 ( .A(keyFF_outputPar[39]), .B(
        key[36]), .S(reset), .Z(keyFF_inputPar[36]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_37_U1 ( .A(keyFF_outputPar[40]), .B(
        key[37]), .S(reset), .Z(keyFF_inputPar[37]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_38_U1 ( .A(keyFF_outputPar[41]), .B(
        key[38]), .S(reset), .Z(keyFF_inputPar[38]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_39_U1 ( .A(keyFF_outputPar[42]), .B(
        key[39]), .S(reset), .Z(keyFF_inputPar[39]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_40_U1 ( .A(keyFF_outputPar[43]), .B(
        key[40]), .S(reset), .Z(keyFF_inputPar[40]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_41_U1 ( .A(keyFF_outputPar[44]), .B(
        key[41]), .S(reset), .Z(keyFF_inputPar[41]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_42_U1 ( .A(keyFF_outputPar[45]), .B(
        key[42]), .S(reset), .Z(keyFF_inputPar[42]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_43_U1 ( .A(keyFF_outputPar[46]), .B(
        key[43]), .S(reset), .Z(keyFF_inputPar[43]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_44_U1 ( .A(keyFF_outputPar[47]), .B(
        key[44]), .S(reset), .Z(keyFF_inputPar[44]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_45_U1 ( .A(keyFF_outputPar[48]), .B(
        key[45]), .S(reset), .Z(keyFF_inputPar[45]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_46_U1 ( .A(keyFF_outputPar[49]), .B(
        key[46]), .S(reset), .Z(keyFF_inputPar[46]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_47_U1 ( .A(keyFF_outputPar[50]), .B(
        key[47]), .S(reset), .Z(keyFF_inputPar[47]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_48_U1 ( .A(keyFF_outputPar[51]), .B(
        key[48]), .S(reset), .Z(keyFF_inputPar[48]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_49_U1 ( .A(keyFF_outputPar[52]), .B(
        key[49]), .S(reset), .Z(keyFF_inputPar[49]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_50_U1 ( .A(keyFF_outputPar[53]), .B(
        key[50]), .S(reset), .Z(keyFF_inputPar[50]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_51_U1 ( .A(keyFF_outputPar[54]), .B(
        key[51]), .S(reset), .Z(keyFF_inputPar[51]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_52_U1 ( .A(keyFF_outputPar[55]), .B(
        key[52]), .S(reset), .Z(keyFF_inputPar[52]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_53_U1 ( .A(keyFF_outputPar[56]), .B(
        key[53]), .S(reset), .Z(keyFF_inputPar[53]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_54_U1 ( .A(keyFF_outputPar[57]), .B(
        key[54]), .S(reset), .Z(keyFF_inputPar[54]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_55_U1 ( .A(keyFF_outputPar[58]), .B(
        key[55]), .S(reset), .Z(keyFF_inputPar[55]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_56_U1 ( .A(keyFF_outputPar[59]), .B(
        key[56]), .S(reset), .Z(keyFF_inputPar[56]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_57_U1 ( .A(keyFF_outputPar[60]), .B(
        key[57]), .S(reset), .Z(keyFF_inputPar[57]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_58_U1 ( .A(keyFF_outputPar[61]), .B(
        key[58]), .S(reset), .Z(keyFF_inputPar[58]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_59_U1 ( .A(keyFF_outputPar[62]), .B(
        key[59]), .S(reset), .Z(keyFF_inputPar[59]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_60_U1 ( .A(keyFF_outputPar[63]), .B(
        key[60]), .S(reset), .Z(keyFF_inputPar[60]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_61_U1 ( .A(keyFF_outputPar[64]), .B(
        key[61]), .S(reset), .Z(keyFF_inputPar[61]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_62_U1 ( .A(keyFF_outputPar[65]), .B(
        key[62]), .S(reset), .Z(keyFF_inputPar[62]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_63_U1 ( .A(keyFF_outputPar[66]), .B(
        key[63]), .S(reset), .Z(keyFF_inputPar[63]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_64_U1 ( .A(keyFF_outputPar[67]), .B(
        key[64]), .S(reset), .Z(keyFF_inputPar[64]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_65_U1 ( .A(keyFF_outputPar[68]), .B(
        key[65]), .S(reset), .Z(keyFF_inputPar[65]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_66_U1 ( .A(keyFF_outputPar[69]), .B(
        key[66]), .S(reset), .Z(keyFF_inputPar[66]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_67_U1 ( .A(keyFF_outputPar[70]), .B(
        key[67]), .S(reset), .Z(keyFF_inputPar[67]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_68_U1 ( .A(keyFF_outputPar[71]), .B(
        key[68]), .S(reset), .Z(keyFF_inputPar[68]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_69_U1 ( .A(keyFF_outputPar[72]), .B(
        key[69]), .S(reset), .Z(keyFF_inputPar[69]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_70_U1 ( .A(keyFF_outputPar[73]), .B(
        key[70]), .S(reset), .Z(keyFF_inputPar[70]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_71_U1 ( .A(keyFF_outputPar[74]), .B(
        key[71]), .S(reset), .Z(keyFF_inputPar[71]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_72_U1 ( .A(keyFF_outputPar[75]), .B(
        key[72]), .S(reset), .Z(keyFF_inputPar[72]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_73_U1 ( .A(roundkey[0]), .B(key[73]), 
        .S(reset), .Z(keyFF_inputPar[73]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_74_U1 ( .A(roundkey[1]), .B(key[74]), 
        .S(reset), .Z(keyFF_inputPar[74]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_75_U1 ( .A(roundkey[2]), .B(key[75]), 
        .S(reset), .Z(keyFF_inputPar[75]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_76_U1 ( .A(sboxOut[0]), .B(key[76]), .S(
        reset), .Z(keyFF_inputPar[76]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_77_U1 ( .A(sboxOut[1]), .B(key[77]), .S(
        reset), .Z(keyFF_inputPar[77]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_78_U1 ( .A(sboxOut[2]), .B(key[78]), .S(
        reset), .Z(keyFF_inputPar[78]) );
  MUX2_X1 keyFF_MUX_inputPar_mux_inst_79_U1 ( .A(sboxOut[3]), .B(key[79]), .S(
        reset), .Z(keyFF_inputPar[79]) );
  INV_X1 sboxInst_U3 ( .A(sboxInst_L0), .ZN(sboxInst_n1) );
  INV_X1 sboxInst_U2 ( .A(sboxIn[3]), .ZN(sboxInst_n2) );
  INV_X1 sboxInst_U1 ( .A(sboxIn[1]), .ZN(sboxInst_n3) );
  XOR2_X1 sboxInst_XOR1_U1 ( .A(sboxIn[2]), .B(sboxIn[1]), .Z(sboxInst_L0) );
  XOR2_X1 sboxInst_XOR2_U1 ( .A(sboxIn[1]), .B(sboxIn[0]), .Z(sboxInst_L1) );
  XOR2_X1 sboxInst_XOR3_U1 ( .A(sboxInst_L1), .B(sboxIn[3]), .Z(sboxInst_L2)
         );
  XNOR2_X1 sboxInst_XOR16_U1 ( .A(sboxInst_T0), .B(sboxInst_L2), .ZN(
        sboxInst_Q2) );
  XOR2_X1 sboxInst_XOR4_U1 ( .A(sboxIn[3]), .B(sboxIn[0]), .Z(sboxInst_L3) );
  XOR2_X1 sboxInst_XOR5_U1 ( .A(sboxInst_L3), .B(sboxInst_L0), .Z(sboxInst_Q3)
         );
  XOR2_X1 sboxInst_XOR6_U1 ( .A(sboxIn[3]), .B(sboxIn[1]), .Z(sboxInst_L4) );
  XOR2_X1 sboxInst_XOR7_U1 ( .A(sboxInst_T0), .B(sboxInst_T2), .Z(sboxInst_L5)
         );
  XNOR2_X1 sboxInst_XOR8_U1 ( .A(sboxInst_L4), .B(sboxInst_L5), .ZN(
        sboxInst_Q6) );
  XOR2_X1 sboxInst_XOR9_U1 ( .A(sboxInst_L1), .B(sboxIn[2]), .Z(sboxInst_Q7)
         );
  AND2_X1 sboxInst_AND1_U1 ( .A1(sboxInst_n1), .A2(sboxInst_n2), .ZN(
        sboxInst_T0) );
  AND2_X1 sboxInst_AND2_U1 ( .A1(sboxInst_Q2), .A2(sboxInst_Q3), .ZN(
        sboxInst_T1) );
  AND2_X1 sboxInst_AND3_U1 ( .A1(sboxInst_n3), .A2(sboxIn[2]), .ZN(sboxInst_T2) );
  AND2_X1 sboxInst_AND4_U1 ( .A1(sboxInst_Q6), .A2(sboxInst_Q7), .ZN(
        sboxInst_T3) );
  XOR2_X1 sboxInst_XOR10_U1 ( .A(sboxInst_L5), .B(sboxInst_T3), .Z(sboxInst_L7) );
  XOR2_X1 sboxInst_XOR11_U1 ( .A(sboxIn[0]), .B(sboxInst_L7), .Z(sboxOut[3])
         );
  XOR2_X1 sboxInst_XOR12_U1 ( .A(sboxInst_L5), .B(sboxInst_T1), .Z(sboxInst_L8) );
  XOR2_X1 sboxInst_XOR13_U1 ( .A(sboxInst_L1), .B(sboxInst_L8), .Z(sboxOut[2])
         );
  XOR2_X1 sboxInst_XOR14_U1 ( .A(sboxInst_L4), .B(sboxInst_T3), .Z(sboxOut[1])
         );
  XOR2_X1 sboxInst_XOR15_U1 ( .A(sboxInst_L3), .B(sboxInst_T2), .Z(sboxOut[0])
         );
  MUX2_X1 MUX_sboxin_mux_inst_0_U1 ( .A(stateXORroundkey[0]), .B(roundkey[3]), 
        .S(selSbox), .Z(sboxIn[0]) );
  MUX2_X1 MUX_sboxin_mux_inst_1_U1 ( .A(stateXORroundkey[1]), .B(keyRegKS[1]), 
        .S(selSbox), .Z(sboxIn[1]) );
  MUX2_X1 MUX_sboxin_mux_inst_2_U1 ( .A(stateXORroundkey[2]), .B(keyRegKS[2]), 
        .S(selSbox), .Z(sboxIn[2]) );
  MUX2_X1 MUX_sboxin_mux_inst_3_U1 ( .A(stateXORroundkey[3]), .B(keyRegKS[3]), 
        .S(selSbox), .Z(sboxIn[3]) );
  MUX2_X1 MUX_serialIn_mux_inst_0_U1 ( .A(sboxOut[0]), .B(stateXORroundkey[0]), 
        .S(intDone), .Z(serialIn[0]) );
  MUX2_X1 MUX_serialIn_mux_inst_1_U1 ( .A(sboxOut[1]), .B(stateXORroundkey[1]), 
        .S(intDone), .Z(serialIn[1]) );
  MUX2_X1 MUX_serialIn_mux_inst_2_U1 ( .A(sboxOut[2]), .B(stateXORroundkey[2]), 
        .S(intDone), .Z(serialIn[2]) );
  MUX2_X1 MUX_serialIn_mux_inst_3_U1 ( .A(sboxOut[3]), .B(stateXORroundkey[3]), 
        .S(intDone), .Z(serialIn[3]) );
endmodule

