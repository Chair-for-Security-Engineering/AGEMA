
module Sbox(X, Y);
  input  [7:0] X;
  output [7:0] Y;

  wire [3:0] b0, b1, b2, b3, b4, b5, b6, b7;

  
  LUT6 #(.INIT(64'hB14EDE67096C6EED)) b0_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b0[0]));
  LUT6 #(.INIT(64'h68AB4BFA8ACB7A13)) b0_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b0[1]));
  LUT6 #(.INIT(64'h10BDB210C006EAB5)) b0_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b0[2]));
  LUT6 #(.INIT(64'h4F1EAD396F247A04)) b0_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b0[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b0_4 (.I0(b0[0]), .I1(b0[1]), .I2(b0[2]), .I3(b0[3]), .I4(X[6]), .I5(X[7]), .O(Y[0]));

  LUT6 #(.INIT(64'h7BAE007D4C53FC7D)) b1_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b1[0]));
  LUT6 #(.INIT(64'hE61A4C5E97816F7A)) b1_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b1[1]));
  LUT6 #(.INIT(64'h6A450B2EF33486B4)) b1_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b1[2]));
  LUT6 #(.INIT(64'hC870974094EAD8A9)) b1_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b1[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b1_4 (.I0(b1[0]), .I1(b1[1]), .I2(b1[2]), .I3(b1[3]), .I4(X[6]), .I5(X[7]), .O(Y[1]));

  LUT6 #(.INIT(64'hA16387FB3B48B4C6)) b2_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b2[0]));
  LUT6 #(.INIT(64'h23A869A2A428C424)) b2_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b2[1]));
  LUT6 #(.INIT(64'h577D64E03B0C3FFB)) b2_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b2[2]));
  LUT6 #(.INIT(64'hAC39B6C0D6CE2EFC)) b2_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b2[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b2_4 (.I0(b2[0]), .I1(b2[1]), .I2(b2[2]), .I3(b2[3]), .I4(X[6]), .I5(X[7]), .O(Y[2]));

  LUT6 #(.INIT(64'h109020A2193D586A)) b3_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b3[0]));
  LUT6 #(.INIT(64'h2568EA2EFFA8527D)) b3_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b3[1]));
  LUT6 #(.INIT(64'hE9DA849CF6AC6C1B)) b3_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b3[2]));
  LUT6 #(.INIT(64'h4E9DDB76C892FB1B)) b3_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b3[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b3_4 (.I0(b3[0]), .I1(b3[1]), .I2(b3[2]), .I3(b3[3]), .I4(X[6]), .I5(X[7]), .O(Y[3]));

  LUT6 #(.INIT(64'hC2B0F97752B8B11E)) b4_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b4[0]));
  LUT6 #(.INIT(64'hF7F17A494CE30F58)) b4_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b4[1]));
  LUT6 #(.INIT(64'h2624B286BC48ECB4)) b4_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b4[2]));
  LUT6 #(.INIT(64'hF210A3AECE472E53)) b4_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b4[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b4_4 (.I0(b4[0]), .I1(b4[1]), .I2(b4[2]), .I3(b4[3]), .I4(X[6]), .I5(X[7]), .O(Y[4]));

  LUT6 #(.INIT(64'hF8045F7B6D98DD7F)) b5_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b5[0]));
  LUT6 #(.INIT(64'h6BC2AA4E0D787AA4)) b5_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b5[1]));
  LUT6 #(.INIT(64'h7D8DCC4706319E08)) b5_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b5[2]));
  LUT6 #(.INIT(64'h54B248130B4F256F)) b5_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b5[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b5_4 (.I0(b5[0]), .I1(b5[1]), .I2(b5[2]), .I3(b5[3]), .I4(X[6]), .I5(X[7]), .O(Y[5]));

  LUT6 #(.INIT(64'h980A3CC2C2FDB4FF)) b6_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b6[0]));
  LUT6 #(.INIT(64'hE4851B3BF3AB2560)) b6_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b6[1]));
  LUT6 #(.INIT(64'h3F6BCB91B30DB559)) b6_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b6[2]));
  LUT6 #(.INIT(64'h21E0B83325591782)) b6_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b6[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b6_4 (.I0(b6[0]), .I1(b6[1]), .I2(b6[2]), .I3(b6[3]), .I4(X[6]), .I5(X[7]), .O(Y[6]));

  LUT6 #(.INIT(64'h5CAA2EC7BF977090)) b7_0 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b7[0]));
  LUT6 #(.INIT(64'hE7BAC28F866AAC82)) b7_1 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b7[1]));
  LUT6 #(.INIT(64'h4CB3770196CA0329)) b7_2 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b7[2]));
  LUT6 #(.INIT(64'h52379DE7B844E3E1)) b7_3 (.I0(X[0]),  .I1(X[1]),  .I2(X[2]),  .I3(X[3]),  .I4(X[4]), .I5(X[5]), .O(b7[3]));
  LUT6 #(.INIT(64'hFF00F0F0CCCCAAAA)) b7_4 (.I0(b7[0]), .I1(b7[1]), .I2(b7[2]), .I3(b7[3]), .I4(X[6]), .I5(X[7]), .O(Y[7]));

endmodule
