/* modified netlist. Source: module LED in file /LED_round-based/AGEMA/LED.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module LED_GHPC_ANF_Pipeline_d1 (IN_plaintext_s0, IN_key_s0, IN_reset, CLK, IN_key_s1, IN_plaintext_s1, Fresh, OUT_ciphertext_s0, OUT_done, OUT_ciphertext_s1);
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input IN_reset ;
    input CLK ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [63:0] Fresh ;
    output [63:0] OUT_ciphertext_s0 ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_356 ;
    wire signal_375 ;
    wire signal_394 ;
    wire signal_413 ;
    wire signal_432 ;
    wire signal_451 ;
    wire signal_470 ;
    wire signal_489 ;
    wire signal_508 ;
    wire signal_527 ;
    wire signal_546 ;
    wire signal_565 ;
    wire signal_584 ;
    wire signal_603 ;
    wire signal_622 ;
    wire signal_641 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1330 ;
    wire signal_1333 ;
    wire signal_1336 ;
    wire signal_1339 ;
    wire signal_1342 ;
    wire signal_1345 ;
    wire signal_1348 ;
    wire signal_1351 ;
    wire signal_1354 ;
    wire signal_1357 ;
    wire signal_1360 ;
    wire signal_1363 ;
    wire signal_1366 ;
    wire signal_1368 ;
    wire signal_1370 ;
    wire signal_1372 ;
    wire signal_1374 ;
    wire signal_1376 ;
    wire signal_1378 ;
    wire signal_1380 ;
    wire signal_1382 ;
    wire signal_1384 ;
    wire signal_1386 ;
    wire signal_1388 ;
    wire signal_1390 ;
    wire signal_1392 ;
    wire signal_1395 ;
    wire signal_1398 ;
    wire signal_1401 ;
    wire signal_1404 ;
    wire signal_1407 ;
    wire signal_1410 ;
    wire signal_1413 ;
    wire signal_1416 ;
    wire signal_1419 ;
    wire signal_1422 ;
    wire signal_1425 ;
    wire signal_1428 ;
    wire signal_1431 ;
    wire signal_1434 ;
    wire signal_1437 ;
    wire signal_1440 ;
    wire signal_1443 ;
    wire signal_1446 ;
    wire signal_1449 ;
    wire signal_1452 ;
    wire signal_1455 ;
    wire signal_1458 ;
    wire signal_1461 ;
    wire signal_1464 ;
    wire signal_1467 ;
    wire signal_1470 ;
    wire signal_1473 ;
    wire signal_1476 ;
    wire signal_1479 ;
    wire signal_1482 ;
    wire signal_1485 ;
    wire signal_1488 ;
    wire signal_1491 ;
    wire signal_1494 ;
    wire signal_1497 ;
    wire signal_1500 ;
    wire signal_1503 ;
    wire signal_1506 ;
    wire signal_1509 ;
    wire signal_1512 ;
    wire signal_1515 ;
    wire signal_1518 ;
    wire signal_1521 ;
    wire signal_1524 ;
    wire signal_1527 ;
    wire signal_1530 ;
    wire signal_1533 ;
    wire signal_1536 ;
    wire signal_1539 ;
    wire signal_1542 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1554 ;
    wire signal_1556 ;
    wire signal_1558 ;
    wire signal_1560 ;
    wire signal_1562 ;
    wire signal_1564 ;
    wire signal_1566 ;
    wire signal_1568 ;
    wire signal_1570 ;
    wire signal_1572 ;
    wire signal_1574 ;
    wire signal_1576 ;
    wire signal_1578 ;
    wire signal_1580 ;
    wire signal_1582 ;
    wire signal_1584 ;
    wire signal_1586 ;
    wire signal_1588 ;
    wire signal_1590 ;
    wire signal_1592 ;
    wire signal_1594 ;
    wire signal_1596 ;
    wire signal_1598 ;
    wire signal_1600 ;
    wire signal_1602 ;
    wire signal_1604 ;
    wire signal_1606 ;
    wire signal_1608 ;
    wire signal_1610 ;
    wire signal_1612 ;
    wire signal_1614 ;
    wire signal_1616 ;
    wire signal_1618 ;
    wire signal_1620 ;
    wire signal_1622 ;
    wire signal_1624 ;
    wire signal_1626 ;
    wire signal_1628 ;
    wire signal_1630 ;
    wire signal_1632 ;
    wire signal_1634 ;
    wire signal_1636 ;
    wire signal_1638 ;
    wire signal_1640 ;
    wire signal_1642 ;
    wire signal_1644 ;
    wire signal_1646 ;
    wire signal_1648 ;
    wire signal_1650 ;
    wire signal_1652 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1917 ;
    wire signal_1919 ;
    wire signal_1921 ;
    wire signal_1923 ;
    wire signal_1925 ;
    wire signal_1927 ;
    wire signal_1929 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1965 ;
    wire signal_1967 ;
    wire signal_1969 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2001 ;
    wire signal_2003 ;
    wire signal_2005 ;
    wire signal_2007 ;
    wire signal_2009 ;
    wire signal_2011 ;
    wire signal_2013 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2061 ;
    wire signal_2063 ;
    wire signal_2065 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2085 ;
    wire signal_2087 ;
    wire signal_2089 ;
    wire signal_2091 ;
    wire signal_2093 ;
    wire signal_2095 ;
    wire signal_2097 ;
    wire signal_2099 ;
    wire signal_2101 ;
    wire signal_2103 ;
    wire signal_2105 ;
    wire signal_2107 ;
    wire signal_2109 ;
    wire signal_2111 ;
    wire signal_2113 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2141 ;
    wire signal_2143 ;
    wire signal_2145 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2153 ;
    wire signal_2155 ;
    wire signal_2157 ;
    wire signal_2159 ;
    wire signal_2161 ;
    wire signal_2163 ;
    wire signal_2165 ;
    wire signal_2167 ;
    wire signal_2169 ;
    wire signal_2171 ;
    wire signal_2173 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2205 ;
    wire signal_2207 ;
    wire signal_2209 ;
    wire signal_2211 ;
    wire signal_2213 ;
    wire signal_2215 ;
    wire signal_2217 ;
    wire signal_2219 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;

    /* cells in depth 0 */
    NOR2_X1 cell_0 ( .A1 (signal_875), .A2 (signal_878), .ZN (signal_266) ) ;
    NAND2_X1 cell_1 ( .A1 (signal_879), .A2 (signal_266), .ZN (signal_267) ) ;
    NOR2_X1 cell_2 ( .A1 (signal_874), .A2 (signal_267), .ZN (signal_268) ) ;
    NAND2_X1 cell_3 ( .A1 (signal_876), .A2 (signal_268), .ZN (signal_269) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_877), .A2 (signal_269), .ZN (signal_270) ) ;
    NOR2_X1 cell_5 ( .A1 (OUT_done), .A2 (signal_270), .ZN (signal_271) ) ;
    NOR2_X1 cell_6 ( .A1 (IN_reset), .A2 (signal_271), .ZN (signal_265) ) ;
    NAND2_X1 cell_7 ( .A1 (signal_273), .A2 (signal_274), .ZN (signal_272) ) ;
    XNOR2_X1 cell_8 ( .A (signal_304), .B (signal_275), .ZN (signal_274) ) ;
    XOR2_X1 cell_9 ( .A (signal_309), .B (signal_307), .Z (signal_275) ) ;
    NAND2_X1 cell_10 ( .A1 (signal_276), .A2 (signal_277), .ZN (signal_273) ) ;
    NAND2_X1 cell_11 ( .A1 (signal_278), .A2 (signal_279), .ZN (signal_277) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_302), .A2 (signal_289), .ZN (signal_279) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_278) ) ;
    NAND2_X1 cell_14 ( .A1 (signal_289), .A2 (signal_280), .ZN (signal_276) ) ;
    AND2_X1 cell_15 ( .A1 (signal_306), .A2 (signal_309), .ZN (signal_280) ) ;
    NAND2_X1 cell_16 ( .A1 (signal_298), .A2 (signal_283), .ZN (signal_282) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_300), .A2 (signal_284), .ZN (signal_283) ) ;
    NAND2_X1 cell_18 ( .A1 (signal_296), .A2 (signal_876), .ZN (signal_284) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_292), .A2 (signal_290), .ZN (signal_281) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_292), .A2 (IN_reset), .ZN (signal_291) ) ;
    NOR2_X1 cell_21 ( .A1 (IN_reset), .A2 (signal_294), .ZN (signal_293) ) ;
    NOR2_X1 cell_22 ( .A1 (IN_reset), .A2 (signal_296), .ZN (signal_295) ) ;
    NOR2_X1 cell_23 ( .A1 (IN_reset), .A2 (signal_298), .ZN (signal_297) ) ;
    NOR2_X1 cell_24 ( .A1 (IN_reset), .A2 (signal_300), .ZN (signal_299) ) ;
    NOR2_X1 cell_25 ( .A1 (signal_289), .A2 (IN_reset), .ZN (signal_303) ) ;
    NOR2_X1 cell_26 ( .A1 (signal_306), .A2 (IN_reset), .ZN (signal_305) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_309), .A2 (IN_reset), .ZN (signal_308) ) ;
    NOR2_X1 cell_28 ( .A1 (signal_288), .A2 (IN_reset), .ZN (signal_310) ) ;
    OR2_X1 cell_29 ( .A1 (signal_288), .A2 (signal_276), .ZN (signal_286) ) ;
    NAND2_X1 cell_30 ( .A1 (signal_272), .A2 (signal_286), .ZN (signal_311) ) ;
    NOR2_X1 cell_31 ( .A1 (signal_281), .A2 (signal_282), .ZN (signal_340) ) ;
    INV_X1 cell_32 ( .A (signal_286), .ZN (signal_285) ) ;
    OR2_X1 cell_33 ( .A1 (IN_reset), .A2 (signal_287), .ZN (signal_301) ) ;
    XNOR2_X1 cell_34 ( .A (signal_292), .B (signal_290), .ZN (signal_287) ) ;
    INV_X1 cell_35 ( .A (signal_340), .ZN (signal_341) ) ;
    INV_X1 cell_36 ( .A (signal_341), .ZN (signal_344) ) ;
    INV_X1 cell_37 ( .A (signal_341), .ZN (signal_342) ) ;
    INV_X1 cell_38 ( .A (signal_341), .ZN (signal_343) ) ;
    INV_X1 cell_167 ( .A (signal_345), .ZN (signal_346) ) ;
    INV_X1 cell_168 ( .A (signal_285), .ZN (signal_345) ) ;
    INV_X1 cell_169 ( .A (signal_345), .ZN (signal_348) ) ;
    INV_X1 cell_170 ( .A (signal_345), .ZN (signal_347) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_171 ( .s (signal_285), .b ({IN_key_s1[64], IN_key_s0[64]}), .a ({IN_key_s1[0], IN_key_s0[0]}), .c ({signal_1330, signal_1135}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_172 ( .s (signal_346), .b ({IN_key_s1[65], IN_key_s0[65]}), .a ({IN_key_s1[1], IN_key_s0[1]}), .c ({signal_1395, signal_1134}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_173 ( .s (signal_346), .b ({IN_key_s1[66], IN_key_s0[66]}), .a ({IN_key_s1[2], IN_key_s0[2]}), .c ({signal_1398, signal_1133}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_174 ( .s (signal_285), .b ({IN_key_s1[67], IN_key_s0[67]}), .a ({IN_key_s1[3], IN_key_s0[3]}), .c ({signal_1333, signal_1132}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_175 ( .s (signal_346), .b ({IN_key_s1[68], IN_key_s0[68]}), .a ({IN_key_s1[4], IN_key_s0[4]}), .c ({signal_1401, signal_1131}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_176 ( .s (signal_346), .b ({IN_key_s1[69], IN_key_s0[69]}), .a ({IN_key_s1[5], IN_key_s0[5]}), .c ({signal_1404, signal_1130}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_177 ( .s (signal_346), .b ({IN_key_s1[70], IN_key_s0[70]}), .a ({IN_key_s1[6], IN_key_s0[6]}), .c ({signal_1407, signal_1129}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_178 ( .s (signal_346), .b ({IN_key_s1[71], IN_key_s0[71]}), .a ({IN_key_s1[7], IN_key_s0[7]}), .c ({signal_1410, signal_1128}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_179 ( .s (signal_346), .b ({IN_key_s1[72], IN_key_s0[72]}), .a ({IN_key_s1[8], IN_key_s0[8]}), .c ({signal_1413, signal_1127}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_180 ( .s (signal_346), .b ({IN_key_s1[73], IN_key_s0[73]}), .a ({IN_key_s1[9], IN_key_s0[9]}), .c ({signal_1416, signal_1126}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_181 ( .s (signal_346), .b ({IN_key_s1[74], IN_key_s0[74]}), .a ({IN_key_s1[10], IN_key_s0[10]}), .c ({signal_1419, signal_1125}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_182 ( .s (signal_346), .b ({IN_key_s1[75], IN_key_s0[75]}), .a ({IN_key_s1[11], IN_key_s0[11]}), .c ({signal_1422, signal_1124}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_183 ( .s (signal_346), .b ({IN_key_s1[76], IN_key_s0[76]}), .a ({IN_key_s1[12], IN_key_s0[12]}), .c ({signal_1425, signal_1123}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_184 ( .s (signal_346), .b ({IN_key_s1[77], IN_key_s0[77]}), .a ({IN_key_s1[13], IN_key_s0[13]}), .c ({signal_1428, signal_1122}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_185 ( .s (signal_346), .b ({IN_key_s1[78], IN_key_s0[78]}), .a ({IN_key_s1[14], IN_key_s0[14]}), .c ({signal_1431, signal_1121}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_186 ( .s (signal_346), .b ({IN_key_s1[79], IN_key_s0[79]}), .a ({IN_key_s1[15], IN_key_s0[15]}), .c ({signal_1434, signal_1120}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_187 ( .s (signal_285), .b ({IN_key_s1[80], IN_key_s0[80]}), .a ({IN_key_s1[16], IN_key_s0[16]}), .c ({signal_1336, signal_1119}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_188 ( .s (signal_347), .b ({IN_key_s1[81], IN_key_s0[81]}), .a ({IN_key_s1[17], IN_key_s0[17]}), .c ({signal_1437, signal_1118}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_189 ( .s (signal_348), .b ({IN_key_s1[82], IN_key_s0[82]}), .a ({IN_key_s1[18], IN_key_s0[18]}), .c ({signal_1440, signal_1117}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_190 ( .s (signal_285), .b ({IN_key_s1[83], IN_key_s0[83]}), .a ({IN_key_s1[19], IN_key_s0[19]}), .c ({signal_1339, signal_1116}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_191 ( .s (signal_346), .b ({IN_key_s1[84], IN_key_s0[84]}), .a ({IN_key_s1[20], IN_key_s0[20]}), .c ({signal_1443, signal_1115}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_192 ( .s (signal_348), .b ({IN_key_s1[85], IN_key_s0[85]}), .a ({IN_key_s1[21], IN_key_s0[21]}), .c ({signal_1446, signal_1114}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_193 ( .s (signal_285), .b ({IN_key_s1[86], IN_key_s0[86]}), .a ({IN_key_s1[22], IN_key_s0[22]}), .c ({signal_1342, signal_1113}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_194 ( .s (signal_348), .b ({IN_key_s1[87], IN_key_s0[87]}), .a ({IN_key_s1[23], IN_key_s0[23]}), .c ({signal_1449, signal_1112}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_195 ( .s (signal_285), .b ({IN_key_s1[88], IN_key_s0[88]}), .a ({IN_key_s1[24], IN_key_s0[24]}), .c ({signal_1345, signal_1111}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_196 ( .s (signal_348), .b ({IN_key_s1[89], IN_key_s0[89]}), .a ({IN_key_s1[25], IN_key_s0[25]}), .c ({signal_1452, signal_1110}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_197 ( .s (signal_285), .b ({IN_key_s1[90], IN_key_s0[90]}), .a ({IN_key_s1[26], IN_key_s0[26]}), .c ({signal_1348, signal_1109}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_198 ( .s (signal_348), .b ({IN_key_s1[91], IN_key_s0[91]}), .a ({IN_key_s1[27], IN_key_s0[27]}), .c ({signal_1455, signal_1108}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_199 ( .s (signal_285), .b ({IN_key_s1[92], IN_key_s0[92]}), .a ({IN_key_s1[28], IN_key_s0[28]}), .c ({signal_1351, signal_1107}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_200 ( .s (signal_347), .b ({IN_key_s1[93], IN_key_s0[93]}), .a ({IN_key_s1[29], IN_key_s0[29]}), .c ({signal_1458, signal_1106}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_201 ( .s (signal_347), .b ({IN_key_s1[94], IN_key_s0[94]}), .a ({IN_key_s1[30], IN_key_s0[30]}), .c ({signal_1461, signal_1105}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_202 ( .s (signal_347), .b ({IN_key_s1[95], IN_key_s0[95]}), .a ({IN_key_s1[31], IN_key_s0[31]}), .c ({signal_1464, signal_1104}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_203 ( .s (signal_285), .b ({IN_key_s1[96], IN_key_s0[96]}), .a ({IN_key_s1[32], IN_key_s0[32]}), .c ({signal_1354, signal_1103}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_204 ( .s (signal_348), .b ({IN_key_s1[97], IN_key_s0[97]}), .a ({IN_key_s1[33], IN_key_s0[33]}), .c ({signal_1467, signal_1102}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_205 ( .s (signal_285), .b ({IN_key_s1[98], IN_key_s0[98]}), .a ({IN_key_s1[34], IN_key_s0[34]}), .c ({signal_1357, signal_1101}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_206 ( .s (signal_285), .b ({IN_key_s1[99], IN_key_s0[99]}), .a ({IN_key_s1[35], IN_key_s0[35]}), .c ({signal_1360, signal_1100}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_207 ( .s (signal_285), .b ({IN_key_s1[100], IN_key_s0[100]}), .a ({IN_key_s1[36], IN_key_s0[36]}), .c ({signal_1363, signal_1099}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_208 ( .s (signal_347), .b ({IN_key_s1[101], IN_key_s0[101]}), .a ({IN_key_s1[37], IN_key_s0[37]}), .c ({signal_1470, signal_1098}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_209 ( .s (signal_347), .b ({IN_key_s1[102], IN_key_s0[102]}), .a ({IN_key_s1[38], IN_key_s0[38]}), .c ({signal_1473, signal_1097}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_210 ( .s (signal_285), .b ({IN_key_s1[103], IN_key_s0[103]}), .a ({IN_key_s1[39], IN_key_s0[39]}), .c ({signal_1366, signal_1096}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_211 ( .s (signal_347), .b ({IN_key_s1[104], IN_key_s0[104]}), .a ({IN_key_s1[40], IN_key_s0[40]}), .c ({signal_1476, signal_1095}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_212 ( .s (signal_347), .b ({IN_key_s1[105], IN_key_s0[105]}), .a ({IN_key_s1[41], IN_key_s0[41]}), .c ({signal_1479, signal_1094}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_213 ( .s (signal_347), .b ({IN_key_s1[106], IN_key_s0[106]}), .a ({IN_key_s1[42], IN_key_s0[42]}), .c ({signal_1482, signal_1093}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_214 ( .s (signal_347), .b ({IN_key_s1[107], IN_key_s0[107]}), .a ({IN_key_s1[43], IN_key_s0[43]}), .c ({signal_1485, signal_1092}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_215 ( .s (signal_347), .b ({IN_key_s1[108], IN_key_s0[108]}), .a ({IN_key_s1[44], IN_key_s0[44]}), .c ({signal_1488, signal_1091}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_216 ( .s (signal_347), .b ({IN_key_s1[109], IN_key_s0[109]}), .a ({IN_key_s1[45], IN_key_s0[45]}), .c ({signal_1491, signal_1090}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_217 ( .s (signal_347), .b ({IN_key_s1[110], IN_key_s0[110]}), .a ({IN_key_s1[46], IN_key_s0[46]}), .c ({signal_1494, signal_1089}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_218 ( .s (signal_347), .b ({IN_key_s1[111], IN_key_s0[111]}), .a ({IN_key_s1[47], IN_key_s0[47]}), .c ({signal_1497, signal_1088}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_219 ( .s (signal_347), .b ({IN_key_s1[112], IN_key_s0[112]}), .a ({IN_key_s1[48], IN_key_s0[48]}), .c ({signal_1500, signal_1087}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_220 ( .s (signal_347), .b ({IN_key_s1[113], IN_key_s0[113]}), .a ({IN_key_s1[49], IN_key_s0[49]}), .c ({signal_1503, signal_1086}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_221 ( .s (signal_347), .b ({IN_key_s1[114], IN_key_s0[114]}), .a ({IN_key_s1[50], IN_key_s0[50]}), .c ({signal_1506, signal_1085}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_222 ( .s (signal_347), .b ({IN_key_s1[115], IN_key_s0[115]}), .a ({IN_key_s1[51], IN_key_s0[51]}), .c ({signal_1509, signal_1084}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_223 ( .s (signal_348), .b ({IN_key_s1[116], IN_key_s0[116]}), .a ({IN_key_s1[52], IN_key_s0[52]}), .c ({signal_1512, signal_1083}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_224 ( .s (signal_348), .b ({IN_key_s1[117], IN_key_s0[117]}), .a ({IN_key_s1[53], IN_key_s0[53]}), .c ({signal_1515, signal_1082}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_225 ( .s (signal_348), .b ({IN_key_s1[118], IN_key_s0[118]}), .a ({IN_key_s1[54], IN_key_s0[54]}), .c ({signal_1518, signal_1081}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_226 ( .s (signal_348), .b ({IN_key_s1[119], IN_key_s0[119]}), .a ({IN_key_s1[55], IN_key_s0[55]}), .c ({signal_1521, signal_1080}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_227 ( .s (signal_348), .b ({IN_key_s1[120], IN_key_s0[120]}), .a ({IN_key_s1[56], IN_key_s0[56]}), .c ({signal_1524, signal_1079}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_228 ( .s (signal_348), .b ({IN_key_s1[121], IN_key_s0[121]}), .a ({IN_key_s1[57], IN_key_s0[57]}), .c ({signal_1527, signal_1078}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_229 ( .s (signal_348), .b ({IN_key_s1[122], IN_key_s0[122]}), .a ({IN_key_s1[58], IN_key_s0[58]}), .c ({signal_1530, signal_1077}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_230 ( .s (signal_348), .b ({IN_key_s1[123], IN_key_s0[123]}), .a ({IN_key_s1[59], IN_key_s0[59]}), .c ({signal_1533, signal_1076}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_231 ( .s (signal_348), .b ({IN_key_s1[124], IN_key_s0[124]}), .a ({IN_key_s1[60], IN_key_s0[60]}), .c ({signal_1536, signal_1075}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_232 ( .s (signal_348), .b ({IN_key_s1[125], IN_key_s0[125]}), .a ({IN_key_s1[61], IN_key_s0[61]}), .c ({signal_1539, signal_1074}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_233 ( .s (signal_348), .b ({IN_key_s1[126], IN_key_s0[126]}), .a ({IN_key_s1[62], IN_key_s0[62]}), .c ({signal_1542, signal_1073}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_234 ( .s (signal_348), .b ({IN_key_s1[127], IN_key_s0[127]}), .a ({IN_key_s1[63], IN_key_s0[63]}), .c ({signal_1545, signal_1072}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_235 ( .a ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .b ({signal_1416, signal_1126}), .c ({signal_1554, signal_1062}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_236 ( .a ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .b ({signal_1413, signal_1127}), .c ({signal_1556, signal_1063}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_237 ( .a ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .b ({signal_1410, signal_1128}), .c ({signal_1558, signal_1064}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_238 ( .a ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .b ({signal_1407, signal_1129}), .c ({signal_1560, signal_1065}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_239 ( .a ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .b ({signal_1545, signal_1072}), .c ({signal_1562, signal_1008}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_240 ( .a ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .b ({signal_1542, signal_1073}), .c ({signal_1564, signal_1009}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_241 ( .a ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .b ({signal_1539, signal_1074}), .c ({signal_1566, signal_1010}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_242 ( .a ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .b ({signal_1536, signal_1075}), .c ({signal_1568, signal_1011}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_243 ( .a ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .b ({signal_1404, signal_1130}), .c ({signal_1570, signal_1066}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_244 ( .a ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .b ({signal_1533, signal_1076}), .c ({signal_1572, signal_1012}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_245 ( .a ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .b ({signal_1530, signal_1077}), .c ({signal_1574, signal_1013}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_246 ( .a ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .b ({signal_1527, signal_1078}), .c ({signal_1576, signal_1014}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_247 ( .a ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .b ({signal_1524, signal_1079}), .c ({signal_1578, signal_1015}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_248 ( .a ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .b ({signal_1521, signal_1080}), .c ({signal_1580, signal_1016}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_249 ( .a ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .b ({signal_1518, signal_1081}), .c ({signal_1582, signal_1017}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_250 ( .a ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .b ({signal_1515, signal_1082}), .c ({signal_1584, signal_1018}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_251 ( .a ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .b ({signal_1512, signal_1083}), .c ({signal_1586, signal_1019}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_252 ( .a ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .b ({signal_1509, signal_1084}), .c ({signal_1588, signal_1020}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_253 ( .a ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .b ({signal_1506, signal_1085}), .c ({signal_1590, signal_1021}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_254 ( .a ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .b ({signal_1401, signal_1131}), .c ({signal_1592, signal_1067}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_255 ( .a ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .b ({signal_1503, signal_1086}), .c ({signal_1594, signal_1022}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_256 ( .a ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .b ({signal_1500, signal_1087}), .c ({signal_1596, signal_1023}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_257 ( .a ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .b ({signal_1497, signal_1088}), .c ({signal_1598, signal_1024}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_258 ( .a ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .b ({signal_1494, signal_1089}), .c ({signal_1600, signal_1025}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_259 ( .a ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .b ({signal_1491, signal_1090}), .c ({signal_1602, signal_1026}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_260 ( .a ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .b ({signal_1488, signal_1091}), .c ({signal_1604, signal_1027}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_261 ( .a ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .b ({signal_1485, signal_1092}), .c ({signal_1606, signal_1028}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_262 ( .a ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .b ({signal_1482, signal_1093}), .c ({signal_1608, signal_1029}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_263 ( .a ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .b ({signal_1479, signal_1094}), .c ({signal_1610, signal_1030}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_264 ( .a ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .b ({signal_1476, signal_1095}), .c ({signal_1612, signal_1031}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_265 ( .a ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .b ({signal_1333, signal_1132}), .c ({signal_1368, signal_1068}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_266 ( .a ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .b ({signal_1366, signal_1096}), .c ({signal_1370, signal_1032}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_267 ( .a ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .b ({signal_1473, signal_1097}), .c ({signal_1614, signal_1033}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_268 ( .a ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .b ({signal_1470, signal_1098}), .c ({signal_1616, signal_1034}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_269 ( .a ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .b ({signal_1363, signal_1099}), .c ({signal_1372, signal_1035}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_270 ( .a ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .b ({signal_1360, signal_1100}), .c ({signal_1374, signal_1036}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_271 ( .a ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .b ({signal_1357, signal_1101}), .c ({signal_1376, signal_1037}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_272 ( .a ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .b ({signal_1467, signal_1102}), .c ({signal_1618, signal_1038}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_273 ( .a ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .b ({signal_1354, signal_1103}), .c ({signal_1378, signal_1039}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_274 ( .a ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .b ({signal_1464, signal_1104}), .c ({signal_1620, signal_1040}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_275 ( .a ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .b ({signal_1461, signal_1105}), .c ({signal_1622, signal_1041}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_276 ( .a ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .b ({signal_1398, signal_1133}), .c ({signal_1624, signal_1069}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_277 ( .a ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .b ({signal_1458, signal_1106}), .c ({signal_1626, signal_1042}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_278 ( .a ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .b ({signal_1351, signal_1107}), .c ({signal_1380, signal_1043}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_279 ( .a ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .b ({signal_1455, signal_1108}), .c ({signal_1628, signal_1044}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_280 ( .a ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .b ({signal_1348, signal_1109}), .c ({signal_1382, signal_1045}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_281 ( .a ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .b ({signal_1452, signal_1110}), .c ({signal_1630, signal_1046}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_282 ( .a ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .b ({signal_1345, signal_1111}), .c ({signal_1384, signal_1047}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_283 ( .a ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .b ({signal_1449, signal_1112}), .c ({signal_1632, signal_1048}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_284 ( .a ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .b ({signal_1342, signal_1113}), .c ({signal_1386, signal_1049}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_285 ( .a ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .b ({signal_1446, signal_1114}), .c ({signal_1634, signal_1050}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_286 ( .a ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .b ({signal_1443, signal_1115}), .c ({signal_1636, signal_1051}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_287 ( .a ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .b ({signal_1395, signal_1134}), .c ({signal_1638, signal_1070}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_288 ( .a ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .b ({signal_1339, signal_1116}), .c ({signal_1388, signal_1052}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_289 ( .a ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .b ({signal_1440, signal_1117}), .c ({signal_1640, signal_1053}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_290 ( .a ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .b ({signal_1437, signal_1118}), .c ({signal_1642, signal_1054}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_291 ( .a ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .b ({signal_1336, signal_1119}), .c ({signal_1390, signal_1055}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_292 ( .a ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .b ({signal_1434, signal_1120}), .c ({signal_1644, signal_1056}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_293 ( .a ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .b ({signal_1431, signal_1121}), .c ({signal_1646, signal_1057}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_294 ( .a ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .b ({signal_1428, signal_1122}), .c ({signal_1648, signal_1058}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_295 ( .a ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .b ({signal_1425, signal_1123}), .c ({signal_1650, signal_1059}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_296 ( .a ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .b ({signal_1422, signal_1124}), .c ({signal_1652, signal_1060}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_297 ( .a ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .b ({signal_1419, signal_1125}), .c ({signal_1654, signal_1061}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_298 ( .a ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .b ({signal_1330, signal_1135}), .c ({signal_1392, signal_1071}) ) ;
    INV_X1 cell_299 ( .A (signal_349), .ZN (signal_351) ) ;
    INV_X1 cell_300 ( .A (signal_311), .ZN (signal_349) ) ;
    INV_X1 cell_301 ( .A (signal_349), .ZN (signal_350) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_302 ( .s (signal_311), .b ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .a ({signal_1392, signal_1071}), .c ({signal_1546, signal_312}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_303 ( .s (signal_311), .b ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .a ({signal_1638, signal_1070}), .c ({signal_1666, signal_313}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_304 ( .s (signal_311), .b ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .a ({signal_1624, signal_1069}), .c ({signal_1667, signal_314}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_305 ( .s (signal_311), .b ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .a ({signal_1368, signal_1068}), .c ({signal_1547, signal_315}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_306 ( .s (signal_350), .b ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .a ({signal_1592, signal_1067}), .c ({signal_1668, signal_316}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_307 ( .s (signal_350), .b ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .a ({signal_1570, signal_1066}), .c ({signal_1669, signal_317}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_308 ( .s (signal_350), .b ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .a ({signal_1560, signal_1065}), .c ({signal_1670, signal_318}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_309 ( .s (signal_350), .b ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .a ({signal_1558, signal_1064}), .c ({signal_1671, signal_1000}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_310 ( .s (signal_350), .b ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .a ({signal_1556, signal_1063}), .c ({signal_1672, signal_999}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_311 ( .s (signal_350), .b ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .a ({signal_1554, signal_1062}), .c ({signal_1673, signal_998}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_312 ( .s (signal_350), .b ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .a ({signal_1654, signal_1061}), .c ({signal_1674, signal_997}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_313 ( .s (signal_350), .b ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .a ({signal_1652, signal_1060}), .c ({signal_1675, signal_996}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_314 ( .s (signal_350), .b ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .a ({signal_1650, signal_1059}), .c ({signal_1676, signal_995}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_315 ( .s (signal_350), .b ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .a ({signal_1648, signal_1058}), .c ({signal_1677, signal_994}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_316 ( .s (signal_350), .b ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .a ({signal_1646, signal_1057}), .c ({signal_1678, signal_993}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_317 ( .s (signal_350), .b ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .a ({signal_1644, signal_1056}), .c ({signal_1679, signal_992}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_318 ( .s (signal_311), .b ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .a ({signal_1390, signal_1055}), .c ({signal_1548, signal_319}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_319 ( .s (signal_311), .b ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .a ({signal_1642, signal_1054}), .c ({signal_1680, signal_320}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_320 ( .s (signal_311), .b ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .a ({signal_1640, signal_1053}), .c ({signal_1681, signal_321}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_321 ( .s (signal_311), .b ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .a ({signal_1388, signal_1052}), .c ({signal_1549, signal_322}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_322 ( .s (signal_350), .b ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .a ({signal_1636, signal_1051}), .c ({signal_1682, signal_323}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_323 ( .s (signal_311), .b ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .a ({signal_1634, signal_1050}), .c ({signal_1683, signal_324}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_324 ( .s (signal_311), .b ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .a ({signal_1386, signal_1049}), .c ({signal_1550, signal_325}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_325 ( .s (signal_311), .b ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .a ({signal_1632, signal_1048}), .c ({signal_1684, signal_984}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_326 ( .s (signal_311), .b ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .a ({signal_1384, signal_1047}), .c ({signal_1551, signal_983}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_327 ( .s (signal_311), .b ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .a ({signal_1630, signal_1046}), .c ({signal_1685, signal_982}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_328 ( .s (signal_311), .b ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .a ({signal_1382, signal_1045}), .c ({signal_1552, signal_981}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_329 ( .s (signal_311), .b ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .a ({signal_1628, signal_1044}), .c ({signal_1686, signal_980}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_330 ( .s (signal_351), .b ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .a ({signal_1380, signal_1043}), .c ({signal_1655, signal_979}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_331 ( .s (signal_351), .b ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .a ({signal_1626, signal_1042}), .c ({signal_1687, signal_978}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_332 ( .s (signal_351), .b ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .a ({signal_1622, signal_1041}), .c ({signal_1688, signal_977}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_333 ( .s (signal_351), .b ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .a ({signal_1620, signal_1040}), .c ({signal_1689, signal_976}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_334 ( .s (signal_351), .b ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .a ({signal_1378, signal_1039}), .c ({signal_1656, signal_326}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_335 ( .s (signal_351), .b ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .a ({signal_1618, signal_1038}), .c ({signal_1690, signal_327}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_336 ( .s (signal_351), .b ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .a ({signal_1376, signal_1037}), .c ({signal_1657, signal_328}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_337 ( .s (signal_351), .b ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .a ({signal_1374, signal_1036}), .c ({signal_1658, signal_329}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_338 ( .s (signal_351), .b ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .a ({signal_1372, signal_1035}), .c ({signal_1659, signal_330}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_339 ( .s (signal_311), .b ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .a ({signal_1616, signal_1034}), .c ({signal_1691, signal_331}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_340 ( .s (signal_351), .b ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .a ({signal_1614, signal_1033}), .c ({signal_1692, signal_332}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_341 ( .s (signal_351), .b ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .a ({signal_1370, signal_1032}), .c ({signal_1660, signal_968}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_342 ( .s (signal_351), .b ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .a ({signal_1612, signal_1031}), .c ({signal_1693, signal_967}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_343 ( .s (signal_351), .b ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .a ({signal_1610, signal_1030}), .c ({signal_1694, signal_966}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_344 ( .s (signal_351), .b ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .a ({signal_1608, signal_1029}), .c ({signal_1695, signal_965}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_345 ( .s (signal_351), .b ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .a ({signal_1606, signal_1028}), .c ({signal_1696, signal_964}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_346 ( .s (signal_351), .b ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .a ({signal_1604, signal_1027}), .c ({signal_1697, signal_963}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_347 ( .s (signal_351), .b ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .a ({signal_1602, signal_1026}), .c ({signal_1698, signal_962}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_348 ( .s (signal_351), .b ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .a ({signal_1600, signal_1025}), .c ({signal_1699, signal_961}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_349 ( .s (signal_351), .b ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .a ({signal_1598, signal_1024}), .c ({signal_1700, signal_960}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_350 ( .s (signal_351), .b ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .a ({signal_1596, signal_1023}), .c ({signal_1701, signal_333}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_351 ( .s (signal_351), .b ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .a ({signal_1594, signal_1022}), .c ({signal_1702, signal_334}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_352 ( .s (signal_311), .b ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .a ({signal_1590, signal_1021}), .c ({signal_1703, signal_335}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_353 ( .s (signal_351), .b ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .a ({signal_1588, signal_1020}), .c ({signal_1704, signal_336}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_354 ( .s (signal_351), .b ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .a ({signal_1586, signal_1019}), .c ({signal_1705, signal_337}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_355 ( .s (signal_351), .b ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .a ({signal_1584, signal_1018}), .c ({signal_1706, signal_338}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_356 ( .s (signal_351), .b ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .a ({signal_1582, signal_1017}), .c ({signal_1707, signal_339}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_357 ( .s (signal_351), .b ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .a ({signal_1580, signal_1016}), .c ({signal_1708, signal_952}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_358 ( .s (signal_351), .b ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .a ({signal_1578, signal_1015}), .c ({signal_1709, signal_951}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_359 ( .s (signal_351), .b ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .a ({signal_1576, signal_1014}), .c ({signal_1710, signal_950}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_360 ( .s (signal_351), .b ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .a ({signal_1574, signal_1013}), .c ({signal_1711, signal_949}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_361 ( .s (signal_351), .b ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .a ({signal_1572, signal_1012}), .c ({signal_1712, signal_948}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_362 ( .s (signal_351), .b ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .a ({signal_1568, signal_1011}), .c ({signal_1713, signal_947}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_363 ( .s (signal_351), .b ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .a ({signal_1566, signal_1010}), .c ({signal_1714, signal_946}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_364 ( .s (signal_351), .b ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .a ({signal_1564, signal_1009}), .c ({signal_1715, signal_945}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_365 ( .s (signal_351), .b ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .a ({signal_1562, signal_1008}), .c ({signal_1716, signal_944}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_366 ( .a ({1'b0, signal_874}), .b ({signal_1670, signal_318}), .c ({signal_1721, signal_1001}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_367 ( .a ({1'b0, signal_875}), .b ({signal_1669, signal_317}), .c ({signal_1722, signal_1002}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_368 ( .a ({1'b0, signal_877}), .b ({signal_1707, signal_339}), .c ({signal_1723, signal_953}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_369 ( .a ({1'b0, signal_878}), .b ({signal_1706, signal_338}), .c ({signal_1724, signal_954}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_370 ( .a ({1'b0, signal_879}), .b ({signal_1705, signal_337}), .c ({signal_1725, signal_955}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_371 ( .a ({1'b0, 1'b0}), .b ({signal_1704, signal_336}), .c ({signal_1726, signal_956}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_372 ( .a ({1'b0, 1'b0}), .b ({signal_1703, signal_335}), .c ({signal_1727, signal_957}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_373 ( .a ({1'b0, signal_876}), .b ({signal_1668, signal_316}), .c ({signal_1728, signal_1003}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_374 ( .a ({1'b0, 1'b0}), .b ({signal_1702, signal_334}), .c ({signal_1729, signal_958}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_375 ( .a ({1'b0, 1'b0}), .b ({signal_1701, signal_333}), .c ({signal_1730, signal_959}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_376 ( .a ({1'b0, 1'b1}), .b ({signal_1547, signal_315}), .c ({signal_1661, signal_1004}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_377 ( .a ({1'b0, signal_874}), .b ({signal_1692, signal_332}), .c ({signal_1731, signal_969}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_378 ( .a ({1'b0, signal_875}), .b ({signal_1691, signal_331}), .c ({signal_1732, signal_970}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_379 ( .a ({1'b0, signal_876}), .b ({signal_1659, signal_330}), .c ({signal_1717, signal_971}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_380 ( .a ({1'b0, 1'b0}), .b ({signal_1658, signal_329}), .c ({signal_1718, signal_972}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_381 ( .a ({1'b0, 1'b0}), .b ({signal_1657, signal_328}), .c ({signal_1719, signal_973}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_382 ( .a ({1'b0, 1'b0}), .b ({signal_1690, signal_327}), .c ({signal_1733, signal_974}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_383 ( .a ({1'b0, 1'b0}), .b ({signal_1656, signal_326}), .c ({signal_1720, signal_975}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_384 ( .a ({1'b0, 1'b0}), .b ({signal_1667, signal_314}), .c ({signal_1734, signal_1005}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_385 ( .a ({1'b0, signal_877}), .b ({signal_1550, signal_325}), .c ({signal_1662, signal_985}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_386 ( .a ({1'b0, signal_878}), .b ({signal_1683, signal_324}), .c ({signal_1735, signal_986}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_387 ( .a ({1'b0, signal_879}), .b ({signal_1682, signal_323}), .c ({signal_1736, signal_987}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_388 ( .a ({1'b0, 1'b0}), .b ({signal_1666, signal_313}), .c ({signal_1737, signal_1006}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_389 ( .a ({1'b0, 1'b1}), .b ({signal_1549, signal_322}), .c ({signal_1663, signal_988}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_390 ( .a ({1'b0, 1'b0}), .b ({signal_1681, signal_321}), .c ({signal_1738, signal_989}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_391 ( .a ({1'b0, 1'b0}), .b ({signal_1680, signal_320}), .c ({signal_1739, signal_990}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_392 ( .a ({1'b0, 1'b0}), .b ({signal_1548, signal_319}), .c ({signal_1664, signal_991}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_393 ( .a ({1'b0, 1'b0}), .b ({signal_1546, signal_312}), .c ({signal_1665, signal_1007}) ) ;
    INV_X1 cell_978 ( .A (signal_808), .ZN (signal_309) ) ;
    INV_X1 cell_980 ( .A (signal_307), .ZN (signal_306) ) ;
    INV_X1 cell_982 ( .A (signal_304), .ZN (signal_289) ) ;
    INV_X1 cell_984 ( .A (signal_288), .ZN (signal_302) ) ;
    INV_X1 cell_986 ( .A (signal_879), .ZN (signal_300) ) ;
    INV_X1 cell_988 ( .A (signal_878), .ZN (signal_298) ) ;
    INV_X1 cell_990 ( .A (signal_877), .ZN (signal_296) ) ;
    INV_X1 cell_992 ( .A (signal_876), .ZN (signal_294) ) ;
    INV_X1 cell_994 ( .A (signal_875), .ZN (signal_292) ) ;
    INV_X1 cell_996 ( .A (signal_874), .ZN (signal_290) ) ;

    /* cells in depth 1 */
    buf_clk cell_1129 ( .C (CLK), .D (signal_343), .Q (signal_2284) ) ;
    buf_clk cell_1131 ( .C (CLK), .D (signal_312), .Q (signal_2286) ) ;
    buf_clk cell_1133 ( .C (CLK), .D (signal_1546), .Q (signal_2288) ) ;
    buf_clk cell_1135 ( .C (CLK), .D (signal_313), .Q (signal_2290) ) ;
    buf_clk cell_1137 ( .C (CLK), .D (signal_1666), .Q (signal_2292) ) ;
    buf_clk cell_1139 ( .C (CLK), .D (signal_344), .Q (signal_2294) ) ;
    buf_clk cell_1141 ( .C (CLK), .D (signal_314), .Q (signal_2296) ) ;
    buf_clk cell_1143 ( .C (CLK), .D (signal_1667), .Q (signal_2298) ) ;
    buf_clk cell_1145 ( .C (CLK), .D (signal_342), .Q (signal_2300) ) ;
    buf_clk cell_1147 ( .C (CLK), .D (signal_315), .Q (signal_2302) ) ;
    buf_clk cell_1149 ( .C (CLK), .D (signal_1547), .Q (signal_2304) ) ;
    buf_clk cell_1151 ( .C (CLK), .D (signal_316), .Q (signal_2306) ) ;
    buf_clk cell_1153 ( .C (CLK), .D (signal_1668), .Q (signal_2308) ) ;
    buf_clk cell_1155 ( .C (CLK), .D (signal_317), .Q (signal_2310) ) ;
    buf_clk cell_1157 ( .C (CLK), .D (signal_1669), .Q (signal_2312) ) ;
    buf_clk cell_1159 ( .C (CLK), .D (signal_318), .Q (signal_2314) ) ;
    buf_clk cell_1161 ( .C (CLK), .D (signal_1670), .Q (signal_2316) ) ;
    buf_clk cell_1163 ( .C (CLK), .D (signal_1000), .Q (signal_2318) ) ;
    buf_clk cell_1165 ( .C (CLK), .D (signal_1671), .Q (signal_2320) ) ;
    buf_clk cell_1167 ( .C (CLK), .D (signal_999), .Q (signal_2322) ) ;
    buf_clk cell_1169 ( .C (CLK), .D (signal_1672), .Q (signal_2324) ) ;
    buf_clk cell_1171 ( .C (CLK), .D (signal_998), .Q (signal_2326) ) ;
    buf_clk cell_1173 ( .C (CLK), .D (signal_1673), .Q (signal_2328) ) ;
    buf_clk cell_1175 ( .C (CLK), .D (signal_997), .Q (signal_2330) ) ;
    buf_clk cell_1177 ( .C (CLK), .D (signal_1674), .Q (signal_2332) ) ;
    buf_clk cell_1179 ( .C (CLK), .D (signal_996), .Q (signal_2334) ) ;
    buf_clk cell_1181 ( .C (CLK), .D (signal_1675), .Q (signal_2336) ) ;
    buf_clk cell_1183 ( .C (CLK), .D (signal_995), .Q (signal_2338) ) ;
    buf_clk cell_1185 ( .C (CLK), .D (signal_1676), .Q (signal_2340) ) ;
    buf_clk cell_1187 ( .C (CLK), .D (signal_994), .Q (signal_2342) ) ;
    buf_clk cell_1189 ( .C (CLK), .D (signal_1677), .Q (signal_2344) ) ;
    buf_clk cell_1191 ( .C (CLK), .D (signal_993), .Q (signal_2346) ) ;
    buf_clk cell_1193 ( .C (CLK), .D (signal_1678), .Q (signal_2348) ) ;
    buf_clk cell_1195 ( .C (CLK), .D (signal_992), .Q (signal_2350) ) ;
    buf_clk cell_1197 ( .C (CLK), .D (signal_1679), .Q (signal_2352) ) ;
    buf_clk cell_1199 ( .C (CLK), .D (signal_319), .Q (signal_2354) ) ;
    buf_clk cell_1201 ( .C (CLK), .D (signal_1548), .Q (signal_2356) ) ;
    buf_clk cell_1203 ( .C (CLK), .D (signal_320), .Q (signal_2358) ) ;
    buf_clk cell_1205 ( .C (CLK), .D (signal_1680), .Q (signal_2360) ) ;
    buf_clk cell_1207 ( .C (CLK), .D (signal_321), .Q (signal_2362) ) ;
    buf_clk cell_1209 ( .C (CLK), .D (signal_1681), .Q (signal_2364) ) ;
    buf_clk cell_1211 ( .C (CLK), .D (signal_322), .Q (signal_2366) ) ;
    buf_clk cell_1213 ( .C (CLK), .D (signal_1549), .Q (signal_2368) ) ;
    buf_clk cell_1215 ( .C (CLK), .D (signal_323), .Q (signal_2370) ) ;
    buf_clk cell_1217 ( .C (CLK), .D (signal_1682), .Q (signal_2372) ) ;
    buf_clk cell_1219 ( .C (CLK), .D (signal_324), .Q (signal_2374) ) ;
    buf_clk cell_1221 ( .C (CLK), .D (signal_1683), .Q (signal_2376) ) ;
    buf_clk cell_1223 ( .C (CLK), .D (signal_325), .Q (signal_2378) ) ;
    buf_clk cell_1225 ( .C (CLK), .D (signal_1550), .Q (signal_2380) ) ;
    buf_clk cell_1227 ( .C (CLK), .D (signal_984), .Q (signal_2382) ) ;
    buf_clk cell_1229 ( .C (CLK), .D (signal_1684), .Q (signal_2384) ) ;
    buf_clk cell_1231 ( .C (CLK), .D (signal_983), .Q (signal_2386) ) ;
    buf_clk cell_1233 ( .C (CLK), .D (signal_1551), .Q (signal_2388) ) ;
    buf_clk cell_1235 ( .C (CLK), .D (signal_982), .Q (signal_2390) ) ;
    buf_clk cell_1237 ( .C (CLK), .D (signal_1685), .Q (signal_2392) ) ;
    buf_clk cell_1239 ( .C (CLK), .D (signal_981), .Q (signal_2394) ) ;
    buf_clk cell_1241 ( .C (CLK), .D (signal_1552), .Q (signal_2396) ) ;
    buf_clk cell_1243 ( .C (CLK), .D (signal_980), .Q (signal_2398) ) ;
    buf_clk cell_1245 ( .C (CLK), .D (signal_1686), .Q (signal_2400) ) ;
    buf_clk cell_1247 ( .C (CLK), .D (signal_979), .Q (signal_2402) ) ;
    buf_clk cell_1249 ( .C (CLK), .D (signal_1655), .Q (signal_2404) ) ;
    buf_clk cell_1251 ( .C (CLK), .D (signal_978), .Q (signal_2406) ) ;
    buf_clk cell_1253 ( .C (CLK), .D (signal_1687), .Q (signal_2408) ) ;
    buf_clk cell_1255 ( .C (CLK), .D (signal_977), .Q (signal_2410) ) ;
    buf_clk cell_1257 ( .C (CLK), .D (signal_1688), .Q (signal_2412) ) ;
    buf_clk cell_1259 ( .C (CLK), .D (signal_976), .Q (signal_2414) ) ;
    buf_clk cell_1261 ( .C (CLK), .D (signal_1689), .Q (signal_2416) ) ;
    buf_clk cell_1263 ( .C (CLK), .D (signal_326), .Q (signal_2418) ) ;
    buf_clk cell_1265 ( .C (CLK), .D (signal_1656), .Q (signal_2420) ) ;
    buf_clk cell_1267 ( .C (CLK), .D (signal_327), .Q (signal_2422) ) ;
    buf_clk cell_1269 ( .C (CLK), .D (signal_1690), .Q (signal_2424) ) ;
    buf_clk cell_1271 ( .C (CLK), .D (signal_328), .Q (signal_2426) ) ;
    buf_clk cell_1273 ( .C (CLK), .D (signal_1657), .Q (signal_2428) ) ;
    buf_clk cell_1275 ( .C (CLK), .D (signal_329), .Q (signal_2430) ) ;
    buf_clk cell_1277 ( .C (CLK), .D (signal_1658), .Q (signal_2432) ) ;
    buf_clk cell_1279 ( .C (CLK), .D (signal_330), .Q (signal_2434) ) ;
    buf_clk cell_1281 ( .C (CLK), .D (signal_1659), .Q (signal_2436) ) ;
    buf_clk cell_1283 ( .C (CLK), .D (signal_331), .Q (signal_2438) ) ;
    buf_clk cell_1285 ( .C (CLK), .D (signal_1691), .Q (signal_2440) ) ;
    buf_clk cell_1287 ( .C (CLK), .D (signal_332), .Q (signal_2442) ) ;
    buf_clk cell_1289 ( .C (CLK), .D (signal_1692), .Q (signal_2444) ) ;
    buf_clk cell_1291 ( .C (CLK), .D (signal_968), .Q (signal_2446) ) ;
    buf_clk cell_1293 ( .C (CLK), .D (signal_1660), .Q (signal_2448) ) ;
    buf_clk cell_1295 ( .C (CLK), .D (signal_967), .Q (signal_2450) ) ;
    buf_clk cell_1297 ( .C (CLK), .D (signal_1693), .Q (signal_2452) ) ;
    buf_clk cell_1299 ( .C (CLK), .D (signal_966), .Q (signal_2454) ) ;
    buf_clk cell_1301 ( .C (CLK), .D (signal_1694), .Q (signal_2456) ) ;
    buf_clk cell_1303 ( .C (CLK), .D (signal_965), .Q (signal_2458) ) ;
    buf_clk cell_1305 ( .C (CLK), .D (signal_1695), .Q (signal_2460) ) ;
    buf_clk cell_1307 ( .C (CLK), .D (signal_340), .Q (signal_2462) ) ;
    buf_clk cell_1309 ( .C (CLK), .D (signal_964), .Q (signal_2464) ) ;
    buf_clk cell_1311 ( .C (CLK), .D (signal_1696), .Q (signal_2466) ) ;
    buf_clk cell_1313 ( .C (CLK), .D (signal_963), .Q (signal_2468) ) ;
    buf_clk cell_1315 ( .C (CLK), .D (signal_1697), .Q (signal_2470) ) ;
    buf_clk cell_1317 ( .C (CLK), .D (signal_962), .Q (signal_2472) ) ;
    buf_clk cell_1319 ( .C (CLK), .D (signal_1698), .Q (signal_2474) ) ;
    buf_clk cell_1321 ( .C (CLK), .D (signal_961), .Q (signal_2476) ) ;
    buf_clk cell_1323 ( .C (CLK), .D (signal_1699), .Q (signal_2478) ) ;
    buf_clk cell_1325 ( .C (CLK), .D (signal_960), .Q (signal_2480) ) ;
    buf_clk cell_1327 ( .C (CLK), .D (signal_1700), .Q (signal_2482) ) ;
    buf_clk cell_1329 ( .C (CLK), .D (signal_333), .Q (signal_2484) ) ;
    buf_clk cell_1331 ( .C (CLK), .D (signal_1701), .Q (signal_2486) ) ;
    buf_clk cell_1333 ( .C (CLK), .D (signal_334), .Q (signal_2488) ) ;
    buf_clk cell_1335 ( .C (CLK), .D (signal_1702), .Q (signal_2490) ) ;
    buf_clk cell_1337 ( .C (CLK), .D (signal_335), .Q (signal_2492) ) ;
    buf_clk cell_1339 ( .C (CLK), .D (signal_1703), .Q (signal_2494) ) ;
    buf_clk cell_1341 ( .C (CLK), .D (signal_336), .Q (signal_2496) ) ;
    buf_clk cell_1343 ( .C (CLK), .D (signal_1704), .Q (signal_2498) ) ;
    buf_clk cell_1345 ( .C (CLK), .D (signal_337), .Q (signal_2500) ) ;
    buf_clk cell_1347 ( .C (CLK), .D (signal_1705), .Q (signal_2502) ) ;
    buf_clk cell_1349 ( .C (CLK), .D (signal_338), .Q (signal_2504) ) ;
    buf_clk cell_1351 ( .C (CLK), .D (signal_1706), .Q (signal_2506) ) ;
    buf_clk cell_1353 ( .C (CLK), .D (signal_339), .Q (signal_2508) ) ;
    buf_clk cell_1355 ( .C (CLK), .D (signal_1707), .Q (signal_2510) ) ;
    buf_clk cell_1357 ( .C (CLK), .D (signal_952), .Q (signal_2512) ) ;
    buf_clk cell_1359 ( .C (CLK), .D (signal_1708), .Q (signal_2514) ) ;
    buf_clk cell_1361 ( .C (CLK), .D (signal_951), .Q (signal_2516) ) ;
    buf_clk cell_1363 ( .C (CLK), .D (signal_1709), .Q (signal_2518) ) ;
    buf_clk cell_1365 ( .C (CLK), .D (signal_950), .Q (signal_2520) ) ;
    buf_clk cell_1367 ( .C (CLK), .D (signal_1710), .Q (signal_2522) ) ;
    buf_clk cell_1369 ( .C (CLK), .D (signal_949), .Q (signal_2524) ) ;
    buf_clk cell_1371 ( .C (CLK), .D (signal_1711), .Q (signal_2526) ) ;
    buf_clk cell_1373 ( .C (CLK), .D (signal_948), .Q (signal_2528) ) ;
    buf_clk cell_1375 ( .C (CLK), .D (signal_1712), .Q (signal_2530) ) ;
    buf_clk cell_1377 ( .C (CLK), .D (signal_947), .Q (signal_2532) ) ;
    buf_clk cell_1379 ( .C (CLK), .D (signal_1713), .Q (signal_2534) ) ;
    buf_clk cell_1381 ( .C (CLK), .D (signal_946), .Q (signal_2536) ) ;
    buf_clk cell_1383 ( .C (CLK), .D (signal_1714), .Q (signal_2538) ) ;
    buf_clk cell_1385 ( .C (CLK), .D (signal_945), .Q (signal_2540) ) ;
    buf_clk cell_1387 ( .C (CLK), .D (signal_1715), .Q (signal_2542) ) ;
    buf_clk cell_1389 ( .C (CLK), .D (signal_944), .Q (signal_2544) ) ;
    buf_clk cell_1391 ( .C (CLK), .D (signal_1716), .Q (signal_2546) ) ;
    buf_clk cell_1393 ( .C (CLK), .D (IN_reset), .Q (signal_2548) ) ;
    buf_clk cell_1395 ( .C (CLK), .D (IN_plaintext_s0[0]), .Q (signal_2550) ) ;
    buf_clk cell_1397 ( .C (CLK), .D (IN_plaintext_s1[0]), .Q (signal_2552) ) ;
    buf_clk cell_1399 ( .C (CLK), .D (IN_plaintext_s0[1]), .Q (signal_2554) ) ;
    buf_clk cell_1401 ( .C (CLK), .D (IN_plaintext_s1[1]), .Q (signal_2556) ) ;
    buf_clk cell_1403 ( .C (CLK), .D (IN_plaintext_s0[2]), .Q (signal_2558) ) ;
    buf_clk cell_1405 ( .C (CLK), .D (IN_plaintext_s1[2]), .Q (signal_2560) ) ;
    buf_clk cell_1407 ( .C (CLK), .D (IN_plaintext_s0[3]), .Q (signal_2562) ) ;
    buf_clk cell_1409 ( .C (CLK), .D (IN_plaintext_s1[3]), .Q (signal_2564) ) ;
    buf_clk cell_1411 ( .C (CLK), .D (IN_plaintext_s0[4]), .Q (signal_2566) ) ;
    buf_clk cell_1413 ( .C (CLK), .D (IN_plaintext_s1[4]), .Q (signal_2568) ) ;
    buf_clk cell_1415 ( .C (CLK), .D (IN_plaintext_s0[5]), .Q (signal_2570) ) ;
    buf_clk cell_1417 ( .C (CLK), .D (IN_plaintext_s1[5]), .Q (signal_2572) ) ;
    buf_clk cell_1419 ( .C (CLK), .D (IN_plaintext_s0[6]), .Q (signal_2574) ) ;
    buf_clk cell_1421 ( .C (CLK), .D (IN_plaintext_s1[6]), .Q (signal_2576) ) ;
    buf_clk cell_1423 ( .C (CLK), .D (IN_plaintext_s0[7]), .Q (signal_2578) ) ;
    buf_clk cell_1425 ( .C (CLK), .D (IN_plaintext_s1[7]), .Q (signal_2580) ) ;
    buf_clk cell_1427 ( .C (CLK), .D (IN_plaintext_s0[8]), .Q (signal_2582) ) ;
    buf_clk cell_1429 ( .C (CLK), .D (IN_plaintext_s1[8]), .Q (signal_2584) ) ;
    buf_clk cell_1431 ( .C (CLK), .D (IN_plaintext_s0[9]), .Q (signal_2586) ) ;
    buf_clk cell_1433 ( .C (CLK), .D (IN_plaintext_s1[9]), .Q (signal_2588) ) ;
    buf_clk cell_1435 ( .C (CLK), .D (IN_plaintext_s0[10]), .Q (signal_2590) ) ;
    buf_clk cell_1437 ( .C (CLK), .D (IN_plaintext_s1[10]), .Q (signal_2592) ) ;
    buf_clk cell_1439 ( .C (CLK), .D (IN_plaintext_s0[11]), .Q (signal_2594) ) ;
    buf_clk cell_1441 ( .C (CLK), .D (IN_plaintext_s1[11]), .Q (signal_2596) ) ;
    buf_clk cell_1443 ( .C (CLK), .D (IN_plaintext_s0[12]), .Q (signal_2598) ) ;
    buf_clk cell_1445 ( .C (CLK), .D (IN_plaintext_s1[12]), .Q (signal_2600) ) ;
    buf_clk cell_1447 ( .C (CLK), .D (IN_plaintext_s0[13]), .Q (signal_2602) ) ;
    buf_clk cell_1449 ( .C (CLK), .D (IN_plaintext_s1[13]), .Q (signal_2604) ) ;
    buf_clk cell_1451 ( .C (CLK), .D (IN_plaintext_s0[14]), .Q (signal_2606) ) ;
    buf_clk cell_1453 ( .C (CLK), .D (IN_plaintext_s1[14]), .Q (signal_2608) ) ;
    buf_clk cell_1455 ( .C (CLK), .D (IN_plaintext_s0[15]), .Q (signal_2610) ) ;
    buf_clk cell_1457 ( .C (CLK), .D (IN_plaintext_s1[15]), .Q (signal_2612) ) ;
    buf_clk cell_1459 ( .C (CLK), .D (IN_plaintext_s0[16]), .Q (signal_2614) ) ;
    buf_clk cell_1461 ( .C (CLK), .D (IN_plaintext_s1[16]), .Q (signal_2616) ) ;
    buf_clk cell_1463 ( .C (CLK), .D (IN_plaintext_s0[17]), .Q (signal_2618) ) ;
    buf_clk cell_1465 ( .C (CLK), .D (IN_plaintext_s1[17]), .Q (signal_2620) ) ;
    buf_clk cell_1467 ( .C (CLK), .D (IN_plaintext_s0[18]), .Q (signal_2622) ) ;
    buf_clk cell_1469 ( .C (CLK), .D (IN_plaintext_s1[18]), .Q (signal_2624) ) ;
    buf_clk cell_1471 ( .C (CLK), .D (IN_plaintext_s0[19]), .Q (signal_2626) ) ;
    buf_clk cell_1473 ( .C (CLK), .D (IN_plaintext_s1[19]), .Q (signal_2628) ) ;
    buf_clk cell_1475 ( .C (CLK), .D (IN_plaintext_s0[20]), .Q (signal_2630) ) ;
    buf_clk cell_1477 ( .C (CLK), .D (IN_plaintext_s1[20]), .Q (signal_2632) ) ;
    buf_clk cell_1479 ( .C (CLK), .D (IN_plaintext_s0[21]), .Q (signal_2634) ) ;
    buf_clk cell_1481 ( .C (CLK), .D (IN_plaintext_s1[21]), .Q (signal_2636) ) ;
    buf_clk cell_1483 ( .C (CLK), .D (IN_plaintext_s0[22]), .Q (signal_2638) ) ;
    buf_clk cell_1485 ( .C (CLK), .D (IN_plaintext_s1[22]), .Q (signal_2640) ) ;
    buf_clk cell_1487 ( .C (CLK), .D (IN_plaintext_s0[23]), .Q (signal_2642) ) ;
    buf_clk cell_1489 ( .C (CLK), .D (IN_plaintext_s1[23]), .Q (signal_2644) ) ;
    buf_clk cell_1491 ( .C (CLK), .D (IN_plaintext_s0[24]), .Q (signal_2646) ) ;
    buf_clk cell_1493 ( .C (CLK), .D (IN_plaintext_s1[24]), .Q (signal_2648) ) ;
    buf_clk cell_1495 ( .C (CLK), .D (IN_plaintext_s0[25]), .Q (signal_2650) ) ;
    buf_clk cell_1497 ( .C (CLK), .D (IN_plaintext_s1[25]), .Q (signal_2652) ) ;
    buf_clk cell_1499 ( .C (CLK), .D (IN_plaintext_s0[26]), .Q (signal_2654) ) ;
    buf_clk cell_1501 ( .C (CLK), .D (IN_plaintext_s1[26]), .Q (signal_2656) ) ;
    buf_clk cell_1503 ( .C (CLK), .D (IN_plaintext_s0[27]), .Q (signal_2658) ) ;
    buf_clk cell_1505 ( .C (CLK), .D (IN_plaintext_s1[27]), .Q (signal_2660) ) ;
    buf_clk cell_1507 ( .C (CLK), .D (IN_plaintext_s0[28]), .Q (signal_2662) ) ;
    buf_clk cell_1509 ( .C (CLK), .D (IN_plaintext_s1[28]), .Q (signal_2664) ) ;
    buf_clk cell_1511 ( .C (CLK), .D (IN_plaintext_s0[29]), .Q (signal_2666) ) ;
    buf_clk cell_1513 ( .C (CLK), .D (IN_plaintext_s1[29]), .Q (signal_2668) ) ;
    buf_clk cell_1515 ( .C (CLK), .D (IN_plaintext_s0[30]), .Q (signal_2670) ) ;
    buf_clk cell_1517 ( .C (CLK), .D (IN_plaintext_s1[30]), .Q (signal_2672) ) ;
    buf_clk cell_1519 ( .C (CLK), .D (IN_plaintext_s0[31]), .Q (signal_2674) ) ;
    buf_clk cell_1521 ( .C (CLK), .D (IN_plaintext_s1[31]), .Q (signal_2676) ) ;
    buf_clk cell_1523 ( .C (CLK), .D (IN_plaintext_s0[32]), .Q (signal_2678) ) ;
    buf_clk cell_1525 ( .C (CLK), .D (IN_plaintext_s1[32]), .Q (signal_2680) ) ;
    buf_clk cell_1527 ( .C (CLK), .D (IN_plaintext_s0[33]), .Q (signal_2682) ) ;
    buf_clk cell_1529 ( .C (CLK), .D (IN_plaintext_s1[33]), .Q (signal_2684) ) ;
    buf_clk cell_1531 ( .C (CLK), .D (IN_plaintext_s0[34]), .Q (signal_2686) ) ;
    buf_clk cell_1533 ( .C (CLK), .D (IN_plaintext_s1[34]), .Q (signal_2688) ) ;
    buf_clk cell_1535 ( .C (CLK), .D (IN_plaintext_s0[35]), .Q (signal_2690) ) ;
    buf_clk cell_1537 ( .C (CLK), .D (IN_plaintext_s1[35]), .Q (signal_2692) ) ;
    buf_clk cell_1539 ( .C (CLK), .D (IN_plaintext_s0[36]), .Q (signal_2694) ) ;
    buf_clk cell_1541 ( .C (CLK), .D (IN_plaintext_s1[36]), .Q (signal_2696) ) ;
    buf_clk cell_1543 ( .C (CLK), .D (IN_plaintext_s0[37]), .Q (signal_2698) ) ;
    buf_clk cell_1545 ( .C (CLK), .D (IN_plaintext_s1[37]), .Q (signal_2700) ) ;
    buf_clk cell_1547 ( .C (CLK), .D (IN_plaintext_s0[38]), .Q (signal_2702) ) ;
    buf_clk cell_1549 ( .C (CLK), .D (IN_plaintext_s1[38]), .Q (signal_2704) ) ;
    buf_clk cell_1551 ( .C (CLK), .D (IN_plaintext_s0[39]), .Q (signal_2706) ) ;
    buf_clk cell_1553 ( .C (CLK), .D (IN_plaintext_s1[39]), .Q (signal_2708) ) ;
    buf_clk cell_1555 ( .C (CLK), .D (IN_plaintext_s0[40]), .Q (signal_2710) ) ;
    buf_clk cell_1557 ( .C (CLK), .D (IN_plaintext_s1[40]), .Q (signal_2712) ) ;
    buf_clk cell_1559 ( .C (CLK), .D (IN_plaintext_s0[41]), .Q (signal_2714) ) ;
    buf_clk cell_1561 ( .C (CLK), .D (IN_plaintext_s1[41]), .Q (signal_2716) ) ;
    buf_clk cell_1563 ( .C (CLK), .D (IN_plaintext_s0[42]), .Q (signal_2718) ) ;
    buf_clk cell_1565 ( .C (CLK), .D (IN_plaintext_s1[42]), .Q (signal_2720) ) ;
    buf_clk cell_1567 ( .C (CLK), .D (IN_plaintext_s0[43]), .Q (signal_2722) ) ;
    buf_clk cell_1569 ( .C (CLK), .D (IN_plaintext_s1[43]), .Q (signal_2724) ) ;
    buf_clk cell_1571 ( .C (CLK), .D (IN_plaintext_s0[44]), .Q (signal_2726) ) ;
    buf_clk cell_1573 ( .C (CLK), .D (IN_plaintext_s1[44]), .Q (signal_2728) ) ;
    buf_clk cell_1575 ( .C (CLK), .D (IN_plaintext_s0[45]), .Q (signal_2730) ) ;
    buf_clk cell_1577 ( .C (CLK), .D (IN_plaintext_s1[45]), .Q (signal_2732) ) ;
    buf_clk cell_1579 ( .C (CLK), .D (IN_plaintext_s0[46]), .Q (signal_2734) ) ;
    buf_clk cell_1581 ( .C (CLK), .D (IN_plaintext_s1[46]), .Q (signal_2736) ) ;
    buf_clk cell_1583 ( .C (CLK), .D (IN_plaintext_s0[47]), .Q (signal_2738) ) ;
    buf_clk cell_1585 ( .C (CLK), .D (IN_plaintext_s1[47]), .Q (signal_2740) ) ;
    buf_clk cell_1587 ( .C (CLK), .D (IN_plaintext_s0[48]), .Q (signal_2742) ) ;
    buf_clk cell_1589 ( .C (CLK), .D (IN_plaintext_s1[48]), .Q (signal_2744) ) ;
    buf_clk cell_1591 ( .C (CLK), .D (IN_plaintext_s0[49]), .Q (signal_2746) ) ;
    buf_clk cell_1593 ( .C (CLK), .D (IN_plaintext_s1[49]), .Q (signal_2748) ) ;
    buf_clk cell_1595 ( .C (CLK), .D (IN_plaintext_s0[50]), .Q (signal_2750) ) ;
    buf_clk cell_1597 ( .C (CLK), .D (IN_plaintext_s1[50]), .Q (signal_2752) ) ;
    buf_clk cell_1599 ( .C (CLK), .D (IN_plaintext_s0[51]), .Q (signal_2754) ) ;
    buf_clk cell_1601 ( .C (CLK), .D (IN_plaintext_s1[51]), .Q (signal_2756) ) ;
    buf_clk cell_1603 ( .C (CLK), .D (IN_plaintext_s0[52]), .Q (signal_2758) ) ;
    buf_clk cell_1605 ( .C (CLK), .D (IN_plaintext_s1[52]), .Q (signal_2760) ) ;
    buf_clk cell_1607 ( .C (CLK), .D (IN_plaintext_s0[53]), .Q (signal_2762) ) ;
    buf_clk cell_1609 ( .C (CLK), .D (IN_plaintext_s1[53]), .Q (signal_2764) ) ;
    buf_clk cell_1611 ( .C (CLK), .D (IN_plaintext_s0[54]), .Q (signal_2766) ) ;
    buf_clk cell_1613 ( .C (CLK), .D (IN_plaintext_s1[54]), .Q (signal_2768) ) ;
    buf_clk cell_1615 ( .C (CLK), .D (IN_plaintext_s0[55]), .Q (signal_2770) ) ;
    buf_clk cell_1617 ( .C (CLK), .D (IN_plaintext_s1[55]), .Q (signal_2772) ) ;
    buf_clk cell_1619 ( .C (CLK), .D (IN_plaintext_s0[56]), .Q (signal_2774) ) ;
    buf_clk cell_1621 ( .C (CLK), .D (IN_plaintext_s1[56]), .Q (signal_2776) ) ;
    buf_clk cell_1623 ( .C (CLK), .D (IN_plaintext_s0[57]), .Q (signal_2778) ) ;
    buf_clk cell_1625 ( .C (CLK), .D (IN_plaintext_s1[57]), .Q (signal_2780) ) ;
    buf_clk cell_1627 ( .C (CLK), .D (IN_plaintext_s0[58]), .Q (signal_2782) ) ;
    buf_clk cell_1629 ( .C (CLK), .D (IN_plaintext_s1[58]), .Q (signal_2784) ) ;
    buf_clk cell_1631 ( .C (CLK), .D (IN_plaintext_s0[59]), .Q (signal_2786) ) ;
    buf_clk cell_1633 ( .C (CLK), .D (IN_plaintext_s1[59]), .Q (signal_2788) ) ;
    buf_clk cell_1635 ( .C (CLK), .D (IN_plaintext_s0[60]), .Q (signal_2790) ) ;
    buf_clk cell_1637 ( .C (CLK), .D (IN_plaintext_s1[60]), .Q (signal_2792) ) ;
    buf_clk cell_1639 ( .C (CLK), .D (IN_plaintext_s0[61]), .Q (signal_2794) ) ;
    buf_clk cell_1641 ( .C (CLK), .D (IN_plaintext_s1[61]), .Q (signal_2796) ) ;
    buf_clk cell_1643 ( .C (CLK), .D (IN_plaintext_s0[62]), .Q (signal_2798) ) ;
    buf_clk cell_1645 ( .C (CLK), .D (IN_plaintext_s1[62]), .Q (signal_2800) ) ;
    buf_clk cell_1647 ( .C (CLK), .D (IN_plaintext_s0[63]), .Q (signal_2802) ) ;
    buf_clk cell_1649 ( .C (CLK), .D (IN_plaintext_s1[63]), .Q (signal_2804) ) ;
    buf_clk cell_1651 ( .C (CLK), .D (signal_1007), .Q (signal_2806) ) ;
    buf_clk cell_1653 ( .C (CLK), .D (signal_1665), .Q (signal_2808) ) ;
    buf_clk cell_1655 ( .C (CLK), .D (signal_1003), .Q (signal_2810) ) ;
    buf_clk cell_1657 ( .C (CLK), .D (signal_1728), .Q (signal_2812) ) ;
    buf_clk cell_1659 ( .C (CLK), .D (signal_991), .Q (signal_2814) ) ;
    buf_clk cell_1661 ( .C (CLK), .D (signal_1664), .Q (signal_2816) ) ;
    buf_clk cell_1663 ( .C (CLK), .D (signal_987), .Q (signal_2818) ) ;
    buf_clk cell_1665 ( .C (CLK), .D (signal_1736), .Q (signal_2820) ) ;
    buf_clk cell_1667 ( .C (CLK), .D (signal_975), .Q (signal_2822) ) ;
    buf_clk cell_1669 ( .C (CLK), .D (signal_1720), .Q (signal_2824) ) ;
    buf_clk cell_1671 ( .C (CLK), .D (signal_971), .Q (signal_2826) ) ;
    buf_clk cell_1673 ( .C (CLK), .D (signal_1717), .Q (signal_2828) ) ;
    buf_clk cell_1675 ( .C (CLK), .D (signal_959), .Q (signal_2830) ) ;
    buf_clk cell_1677 ( .C (CLK), .D (signal_1730), .Q (signal_2832) ) ;
    buf_clk cell_1679 ( .C (CLK), .D (signal_955), .Q (signal_2834) ) ;
    buf_clk cell_1681 ( .C (CLK), .D (signal_1725), .Q (signal_2836) ) ;
    buf_clk cell_1683 ( .C (CLK), .D (signal_310), .Q (signal_2838) ) ;
    buf_clk cell_1685 ( .C (CLK), .D (signal_308), .Q (signal_2840) ) ;
    buf_clk cell_1687 ( .C (CLK), .D (signal_305), .Q (signal_2842) ) ;
    buf_clk cell_1689 ( .C (CLK), .D (signal_303), .Q (signal_2844) ) ;
    buf_clk cell_1691 ( .C (CLK), .D (signal_301), .Q (signal_2846) ) ;
    buf_clk cell_1693 ( .C (CLK), .D (signal_299), .Q (signal_2848) ) ;
    buf_clk cell_1695 ( .C (CLK), .D (signal_297), .Q (signal_2850) ) ;
    buf_clk cell_1697 ( .C (CLK), .D (signal_295), .Q (signal_2852) ) ;
    buf_clk cell_1699 ( .C (CLK), .D (signal_293), .Q (signal_2854) ) ;
    buf_clk cell_1701 ( .C (CLK), .D (signal_291), .Q (signal_2856) ) ;
    buf_clk cell_1703 ( .C (CLK), .D (signal_265), .Q (signal_2858) ) ;

    /* cells in depth 2 */
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_39 ( .s (signal_2285), .b ({signal_1871, signal_1327}), .a ({signal_2289, signal_2287}), .c ({signal_1888, signal_1263}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_40 ( .s (signal_2285), .b ({signal_1934, signal_1326}), .a ({signal_2293, signal_2291}), .c ({signal_1956, signal_1262}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_41 ( .s (signal_2295), .b ({signal_1870, signal_1325}), .a ({signal_2299, signal_2297}), .c ({signal_1889, signal_1261}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_42 ( .s (signal_2301), .b ({signal_1899, signal_1324}), .a ({signal_2305, signal_2303}), .c ({signal_1912, signal_1260}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_43 ( .s (signal_2301), .b ({signal_1876, signal_1323}), .a ({signal_2309, signal_2307}), .c ({signal_1890, signal_1259}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_44 ( .s (signal_2301), .b ({signal_1940, signal_1322}), .a ({signal_2313, signal_2311}), .c ({signal_1957, signal_1258}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_45 ( .s (signal_2301), .b ({signal_1875, signal_1321}), .a ({signal_2317, signal_2315}), .c ({signal_1891, signal_1257}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_46 ( .s (signal_2301), .b ({signal_1903, signal_1320}), .a ({signal_2321, signal_2319}), .c ({signal_1913, signal_1256}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_47 ( .s (signal_2301), .b ({signal_1881, signal_1319}), .a ({signal_2325, signal_2323}), .c ({signal_1892, signal_1255}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_48 ( .s (signal_2301), .b ({signal_1946, signal_1318}), .a ({signal_2329, signal_2327}), .c ({signal_1958, signal_1254}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_49 ( .s (signal_2301), .b ({signal_1880, signal_1317}), .a ({signal_2333, signal_2331}), .c ({signal_1893, signal_1253}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_50 ( .s (signal_2301), .b ({signal_1907, signal_1316}), .a ({signal_2337, signal_2335}), .c ({signal_1914, signal_1252}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_51 ( .s (signal_2301), .b ({signal_1886, signal_1315}), .a ({signal_2341, signal_2339}), .c ({signal_1894, signal_1251}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_52 ( .s (signal_2301), .b ({signal_1952, signal_1314}), .a ({signal_2345, signal_2343}), .c ({signal_1959, signal_1250}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_53 ( .s (signal_2301), .b ({signal_1885, signal_1313}), .a ({signal_2349, signal_2347}), .c ({signal_1895, signal_1249}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_54 ( .s (signal_2301), .b ({signal_1911, signal_1312}), .a ({signal_2353, signal_2351}), .c ({signal_1915, signal_1248}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_55 ( .s (signal_2285), .b ({signal_1976, signal_1311}), .a ({signal_2357, signal_2355}), .c ({signal_1996, signal_1247}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_56 ( .s (signal_2285), .b ({signal_2022, signal_1310}), .a ({signal_2361, signal_2359}), .c ({signal_2044, signal_1246}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_57 ( .s (signal_2285), .b ({signal_2019, signal_1309}), .a ({signal_2365, signal_2363}), .c ({signal_2045, signal_1245}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_58 ( .s (signal_2285), .b ({signal_1936, signal_1308}), .a ({signal_2369, signal_2367}), .c ({signal_1960, signal_1244}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_59 ( .s (signal_2285), .b ({signal_1982, signal_1307}), .a ({signal_2373, signal_2371}), .c ({signal_1997, signal_1243}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_60 ( .s (signal_2285), .b ({signal_2029, signal_1306}), .a ({signal_2377, signal_2375}), .c ({signal_2046, signal_1242}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_61 ( .s (signal_2285), .b ({signal_2026, signal_1305}), .a ({signal_2381, signal_2379}), .c ({signal_2047, signal_1241}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_62 ( .s (signal_2285), .b ({signal_1942, signal_1304}), .a ({signal_2385, signal_2383}), .c ({signal_1961, signal_1240}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_63 ( .s (signal_2285), .b ({signal_1988, signal_1303}), .a ({signal_2389, signal_2387}), .c ({signal_1998, signal_1239}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_64 ( .s (signal_2285), .b ({signal_2036, signal_1302}), .a ({signal_2393, signal_2391}), .c ({signal_2048, signal_1238}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_65 ( .s (signal_2285), .b ({signal_2033, signal_1301}), .a ({signal_2397, signal_2395}), .c ({signal_2049, signal_1237}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_66 ( .s (signal_2285), .b ({signal_1948, signal_1300}), .a ({signal_2401, signal_2399}), .c ({signal_1962, signal_1236}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_67 ( .s (signal_2295), .b ({signal_1994, signal_1299}), .a ({signal_2405, signal_2403}), .c ({signal_1999, signal_1235}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_68 ( .s (signal_2295), .b ({signal_2043, signal_1298}), .a ({signal_2409, signal_2407}), .c ({signal_2050, signal_1234}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_69 ( .s (signal_2295), .b ({signal_2040, signal_1297}), .a ({signal_2413, signal_2411}), .c ({signal_2051, signal_1233}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_70 ( .s (signal_2295), .b ({signal_1954, signal_1296}), .a ({signal_2417, signal_2415}), .c ({signal_1963, signal_1232}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_71 ( .s (signal_2295), .b ({signal_2018, signal_1295}), .a ({signal_2421, signal_2419}), .c ({signal_2052, signal_1231}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_72 ( .s (signal_2295), .b ({signal_2070, signal_1294}), .a ({signal_2425, signal_2423}), .c ({signal_2080, signal_1230}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_73 ( .s (signal_2295), .b ({signal_2016, signal_1293}), .a ({signal_2429, signal_2427}), .c ({signal_2053, signal_1229}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_74 ( .s (signal_2295), .b ({signal_2118, signal_1292}), .a ({signal_2433, signal_2431}), .c ({signal_2128, signal_1228}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_75 ( .s (signal_2295), .b ({signal_2025, signal_1291}), .a ({signal_2437, signal_2435}), .c ({signal_2054, signal_1227}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_76 ( .s (signal_2295), .b ({signal_2073, signal_1290}), .a ({signal_2441, signal_2439}), .c ({signal_2081, signal_1226}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_77 ( .s (signal_2295), .b ({signal_2023, signal_1289}), .a ({signal_2445, signal_2443}), .c ({signal_2055, signal_1225}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_78 ( .s (signal_2295), .b ({signal_2121, signal_1288}), .a ({signal_2449, signal_2447}), .c ({signal_2129, signal_1224}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_79 ( .s (signal_2295), .b ({signal_2032, signal_1287}), .a ({signal_2453, signal_2451}), .c ({signal_2056, signal_1223}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_80 ( .s (signal_2285), .b ({signal_2076, signal_1286}), .a ({signal_2457, signal_2455}), .c ({signal_2082, signal_1222}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_81 ( .s (signal_2301), .b ({signal_2030, signal_1285}), .a ({signal_2461, signal_2459}), .c ({signal_2057, signal_1221}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_82 ( .s (signal_2463), .b ({signal_2124, signal_1284}), .a ({signal_2467, signal_2465}), .c ({signal_2130, signal_1220}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_83 ( .s (signal_2285), .b ({signal_2039, signal_1283}), .a ({signal_2471, signal_2469}), .c ({signal_2058, signal_1219}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_84 ( .s (signal_2301), .b ({signal_2079, signal_1282}), .a ({signal_2475, signal_2473}), .c ({signal_2083, signal_1218}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_85 ( .s (signal_2295), .b ({signal_2037, signal_1281}), .a ({signal_2479, signal_2477}), .c ({signal_2059, signal_1217}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_86 ( .s (signal_2463), .b ({signal_2127, signal_1280}), .a ({signal_2483, signal_2481}), .c ({signal_2131, signal_1216}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_87 ( .s (signal_2463), .b ({signal_2185, signal_1279}), .a ({signal_2487, signal_2485}), .c ({signal_2192, signal_1215}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_88 ( .s (signal_2463), .b ({signal_2196, signal_1278}), .a ({signal_2491, signal_2489}), .c ({signal_2200, signal_1214}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_89 ( .s (signal_2463), .b ({signal_2117, signal_1277}), .a ({signal_2495, signal_2493}), .c ({signal_2132, signal_1213}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_90 ( .s (signal_2463), .b ({signal_2116, signal_1276}), .a ({signal_2499, signal_2497}), .c ({signal_2133, signal_1212}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_91 ( .s (signal_2463), .b ({signal_2187, signal_1275}), .a ({signal_2503, signal_2501}), .c ({signal_2193, signal_1211}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_92 ( .s (signal_2463), .b ({signal_2197, signal_1274}), .a ({signal_2507, signal_2505}), .c ({signal_2201, signal_1210}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_93 ( .s (signal_2295), .b ({signal_2120, signal_1273}), .a ({signal_2511, signal_2509}), .c ({signal_2134, signal_1209}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_94 ( .s (signal_2285), .b ({signal_2119, signal_1272}), .a ({signal_2515, signal_2513}), .c ({signal_2135, signal_1208}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_95 ( .s (signal_2301), .b ({signal_2189, signal_1271}), .a ({signal_2519, signal_2517}), .c ({signal_2194, signal_1207}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_96 ( .s (signal_2295), .b ({signal_2198, signal_1270}), .a ({signal_2523, signal_2521}), .c ({signal_2202, signal_1206}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_97 ( .s (signal_2285), .b ({signal_2123, signal_1269}), .a ({signal_2527, signal_2525}), .c ({signal_2136, signal_1205}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_98 ( .s (signal_2301), .b ({signal_2122, signal_1268}), .a ({signal_2531, signal_2529}), .c ({signal_2137, signal_1204}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_99 ( .s (signal_2285), .b ({signal_2191, signal_1267}), .a ({signal_2535, signal_2533}), .c ({signal_2195, signal_1203}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_100 ( .s (signal_2301), .b ({signal_2199, signal_1266}), .a ({signal_2539, signal_2537}), .c ({signal_2203, signal_1202}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_101 ( .s (signal_2295), .b ({signal_2126, signal_1265}), .a ({signal_2543, signal_2541}), .c ({signal_2138, signal_1201}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_102 ( .s (signal_2295), .b ({signal_2125, signal_1264}), .a ({signal_2547, signal_2545}), .c ({signal_2139, signal_1200}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_103 ( .s (signal_2549), .b ({signal_1888, signal_1263}), .a ({signal_2553, signal_2551}), .c ({signal_1917, signal_1199}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_104 ( .s (signal_2549), .b ({signal_1956, signal_1262}), .a ({signal_2557, signal_2555}), .c ({signal_2001, signal_1198}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_105 ( .s (signal_2549), .b ({signal_1889, signal_1261}), .a ({signal_2561, signal_2559}), .c ({signal_1919, signal_1197}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_106 ( .s (signal_2549), .b ({signal_1912, signal_1260}), .a ({signal_2565, signal_2563}), .c ({signal_1965, signal_1196}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_107 ( .s (signal_2549), .b ({signal_1890, signal_1259}), .a ({signal_2569, signal_2567}), .c ({signal_1921, signal_1195}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_108 ( .s (signal_2549), .b ({signal_1957, signal_1258}), .a ({signal_2573, signal_2571}), .c ({signal_2003, signal_1194}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_109 ( .s (signal_2549), .b ({signal_1891, signal_1257}), .a ({signal_2577, signal_2575}), .c ({signal_1923, signal_1193}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_110 ( .s (signal_2549), .b ({signal_1913, signal_1256}), .a ({signal_2581, signal_2579}), .c ({signal_1967, signal_1192}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_111 ( .s (signal_2549), .b ({signal_1892, signal_1255}), .a ({signal_2585, signal_2583}), .c ({signal_1925, signal_1191}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_112 ( .s (signal_2549), .b ({signal_1958, signal_1254}), .a ({signal_2589, signal_2587}), .c ({signal_2005, signal_1190}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_113 ( .s (signal_2549), .b ({signal_1893, signal_1253}), .a ({signal_2593, signal_2591}), .c ({signal_1927, signal_1189}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_114 ( .s (signal_2549), .b ({signal_1914, signal_1252}), .a ({signal_2597, signal_2595}), .c ({signal_1969, signal_1188}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_115 ( .s (signal_2549), .b ({signal_1894, signal_1251}), .a ({signal_2601, signal_2599}), .c ({signal_1929, signal_1187}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_116 ( .s (signal_2549), .b ({signal_1959, signal_1250}), .a ({signal_2605, signal_2603}), .c ({signal_2007, signal_1186}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_117 ( .s (signal_2549), .b ({signal_1895, signal_1249}), .a ({signal_2609, signal_2607}), .c ({signal_1931, signal_1185}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_118 ( .s (signal_2549), .b ({signal_1915, signal_1248}), .a ({signal_2613, signal_2611}), .c ({signal_1971, signal_1184}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_119 ( .s (signal_2549), .b ({signal_1996, signal_1247}), .a ({signal_2617, signal_2615}), .c ({signal_2061, signal_1183}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_120 ( .s (signal_2549), .b ({signal_2044, signal_1246}), .a ({signal_2621, signal_2619}), .c ({signal_2085, signal_1182}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_121 ( .s (signal_2549), .b ({signal_2045, signal_1245}), .a ({signal_2625, signal_2623}), .c ({signal_2087, signal_1181}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_122 ( .s (signal_2549), .b ({signal_1960, signal_1244}), .a ({signal_2629, signal_2627}), .c ({signal_2009, signal_1180}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_123 ( .s (signal_2549), .b ({signal_1997, signal_1243}), .a ({signal_2633, signal_2631}), .c ({signal_2063, signal_1179}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_124 ( .s (signal_2549), .b ({signal_2046, signal_1242}), .a ({signal_2637, signal_2635}), .c ({signal_2089, signal_1178}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_125 ( .s (signal_2549), .b ({signal_2047, signal_1241}), .a ({signal_2641, signal_2639}), .c ({signal_2091, signal_1177}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_126 ( .s (signal_2549), .b ({signal_1961, signal_1240}), .a ({signal_2645, signal_2643}), .c ({signal_2011, signal_1176}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_127 ( .s (signal_2549), .b ({signal_1998, signal_1239}), .a ({signal_2649, signal_2647}), .c ({signal_2065, signal_1175}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_128 ( .s (signal_2549), .b ({signal_2048, signal_1238}), .a ({signal_2653, signal_2651}), .c ({signal_2093, signal_1174}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_129 ( .s (signal_2549), .b ({signal_2049, signal_1237}), .a ({signal_2657, signal_2655}), .c ({signal_2095, signal_1173}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_130 ( .s (signal_2549), .b ({signal_1962, signal_1236}), .a ({signal_2661, signal_2659}), .c ({signal_2013, signal_1172}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_131 ( .s (signal_2549), .b ({signal_1999, signal_1235}), .a ({signal_2665, signal_2663}), .c ({signal_2067, signal_1171}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_132 ( .s (signal_2549), .b ({signal_2050, signal_1234}), .a ({signal_2669, signal_2667}), .c ({signal_2097, signal_1170}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_133 ( .s (signal_2549), .b ({signal_2051, signal_1233}), .a ({signal_2673, signal_2671}), .c ({signal_2099, signal_1169}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_134 ( .s (signal_2549), .b ({signal_1963, signal_1232}), .a ({signal_2677, signal_2675}), .c ({signal_2015, signal_1168}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_135 ( .s (signal_2549), .b ({signal_2052, signal_1231}), .a ({signal_2681, signal_2679}), .c ({signal_2101, signal_1167}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_136 ( .s (signal_2549), .b ({signal_2080, signal_1230}), .a ({signal_2685, signal_2683}), .c ({signal_2141, signal_1166}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_137 ( .s (signal_2549), .b ({signal_2053, signal_1229}), .a ({signal_2689, signal_2687}), .c ({signal_2103, signal_1165}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_138 ( .s (signal_2549), .b ({signal_2128, signal_1228}), .a ({signal_2693, signal_2691}), .c ({signal_2153, signal_1164}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_139 ( .s (signal_2549), .b ({signal_2054, signal_1227}), .a ({signal_2697, signal_2695}), .c ({signal_2105, signal_1163}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_140 ( .s (signal_2549), .b ({signal_2081, signal_1226}), .a ({signal_2701, signal_2699}), .c ({signal_2143, signal_1162}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_141 ( .s (signal_2549), .b ({signal_2055, signal_1225}), .a ({signal_2705, signal_2703}), .c ({signal_2107, signal_1161}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_142 ( .s (signal_2549), .b ({signal_2129, signal_1224}), .a ({signal_2709, signal_2707}), .c ({signal_2155, signal_1160}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_143 ( .s (signal_2549), .b ({signal_2056, signal_1223}), .a ({signal_2713, signal_2711}), .c ({signal_2109, signal_1159}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_144 ( .s (signal_2549), .b ({signal_2082, signal_1222}), .a ({signal_2717, signal_2715}), .c ({signal_2145, signal_1158}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_145 ( .s (signal_2549), .b ({signal_2057, signal_1221}), .a ({signal_2721, signal_2719}), .c ({signal_2111, signal_1157}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_146 ( .s (signal_2549), .b ({signal_2130, signal_1220}), .a ({signal_2725, signal_2723}), .c ({signal_2157, signal_1156}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_147 ( .s (signal_2549), .b ({signal_2058, signal_1219}), .a ({signal_2729, signal_2727}), .c ({signal_2113, signal_1155}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_148 ( .s (signal_2549), .b ({signal_2083, signal_1218}), .a ({signal_2733, signal_2731}), .c ({signal_2147, signal_1154}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_149 ( .s (signal_2549), .b ({signal_2059, signal_1217}), .a ({signal_2737, signal_2735}), .c ({signal_2115, signal_1153}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_150 ( .s (signal_2549), .b ({signal_2131, signal_1216}), .a ({signal_2741, signal_2739}), .c ({signal_2159, signal_1152}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_151 ( .s (signal_2549), .b ({signal_2192, signal_1215}), .a ({signal_2745, signal_2743}), .c ({signal_2205, signal_1151}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_152 ( .s (signal_2549), .b ({signal_2200, signal_1214}), .a ({signal_2749, signal_2747}), .c ({signal_2213, signal_1150}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_153 ( .s (signal_2549), .b ({signal_2132, signal_1213}), .a ({signal_2753, signal_2751}), .c ({signal_2161, signal_1149}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_154 ( .s (signal_2549), .b ({signal_2133, signal_1212}), .a ({signal_2757, signal_2755}), .c ({signal_2163, signal_1148}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_155 ( .s (signal_2549), .b ({signal_2193, signal_1211}), .a ({signal_2761, signal_2759}), .c ({signal_2207, signal_1147}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_156 ( .s (signal_2549), .b ({signal_2201, signal_1210}), .a ({signal_2765, signal_2763}), .c ({signal_2215, signal_1146}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_157 ( .s (signal_2549), .b ({signal_2134, signal_1209}), .a ({signal_2769, signal_2767}), .c ({signal_2165, signal_1145}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_158 ( .s (signal_2549), .b ({signal_2135, signal_1208}), .a ({signal_2773, signal_2771}), .c ({signal_2167, signal_1144}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_159 ( .s (signal_2549), .b ({signal_2194, signal_1207}), .a ({signal_2777, signal_2775}), .c ({signal_2209, signal_1143}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_160 ( .s (signal_2549), .b ({signal_2202, signal_1206}), .a ({signal_2781, signal_2779}), .c ({signal_2217, signal_1142}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_161 ( .s (signal_2549), .b ({signal_2136, signal_1205}), .a ({signal_2785, signal_2783}), .c ({signal_2169, signal_1141}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_162 ( .s (signal_2549), .b ({signal_2137, signal_1204}), .a ({signal_2789, signal_2787}), .c ({signal_2171, signal_1140}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_163 ( .s (signal_2549), .b ({signal_2195, signal_1203}), .a ({signal_2793, signal_2791}), .c ({signal_2211, signal_1139}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_164 ( .s (signal_2549), .b ({signal_2203, signal_1202}), .a ({signal_2797, signal_2795}), .c ({signal_2219, signal_1138}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_165 ( .s (signal_2549), .b ({signal_2138, signal_1201}), .a ({signal_2801, signal_2799}), .c ({signal_2173, signal_1137}) ) ;
    mux2_masked #(.low_latency(0), .pipeline(1)) cell_166 ( .s (signal_2549), .b ({signal_2139, signal_1200}), .a ({signal_2805, signal_2803}), .c ({signal_2175, signal_1136}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_412 ( .a ({signal_2809, signal_2807}), .b ({signal_1740, signal_356}), .c ({signal_1812, signal_940}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_435 ( .a ({signal_2813, signal_2811}), .b ({signal_1741, signal_375}), .c ({signal_1813, signal_936}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_458 ( .a ({signal_2325, signal_2323}), .b ({signal_1742, signal_394}), .c ({signal_1814, signal_932}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_481 ( .a ({signal_2341, signal_2339}), .b ({signal_1743, signal_413}), .c ({signal_1815, signal_928}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_504 ( .a ({signal_2817, signal_2815}), .b ({signal_1744, signal_432}), .c ({signal_1816, signal_924}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_527 ( .a ({signal_2821, signal_2819}), .b ({signal_1745, signal_451}), .c ({signal_1817, signal_920}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_550 ( .a ({signal_2389, signal_2387}), .b ({signal_1746, signal_470}), .c ({signal_1818, signal_916}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_573 ( .a ({signal_2405, signal_2403}), .b ({signal_1747, signal_489}), .c ({signal_1819, signal_912}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_596 ( .a ({signal_2825, signal_2823}), .b ({signal_1748, signal_508}), .c ({signal_1820, signal_908}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_619 ( .a ({signal_2829, signal_2827}), .b ({signal_1749, signal_527}), .c ({signal_1821, signal_904}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_642 ( .a ({signal_2453, signal_2451}), .b ({signal_1750, signal_546}), .c ({signal_1822, signal_900}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_665 ( .a ({signal_2471, signal_2469}), .b ({signal_1751, signal_565}), .c ({signal_1823, signal_896}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_688 ( .a ({signal_2833, signal_2831}), .b ({signal_1752, signal_584}), .c ({signal_1824, signal_892}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_711 ( .a ({signal_2837, signal_2835}), .b ({signal_1753, signal_603}), .c ({signal_1825, signal_888}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_734 ( .a ({signal_2519, signal_2517}), .b ({signal_1754, signal_622}), .c ({signal_1826, signal_884}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_757 ( .a ({signal_2535, signal_2533}), .b ({signal_1755, signal_641}), .c ({signal_1827, signal_880}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_762 ( .a ({signal_2068, signal_656}), .b ({signal_1932, signal_657}), .c ({signal_2116, signal_1276}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_763 ( .a ({signal_1899, signal_1324}), .b ({signal_1773, signal_882}), .c ({signal_1932, signal_657}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_764 ( .a ({signal_2016, signal_1293}), .b ({signal_2019, signal_1309}), .c ({signal_2068, signal_656}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_765 ( .a ({signal_1896, signal_658}), .b ({signal_1977, signal_659}), .c ({signal_2016, signal_1293}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_766 ( .a ({signal_1772, signal_881}), .b ({signal_1869, signal_660}), .c ({signal_1896, signal_658}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_767 ( .a ({signal_2017, signal_661}), .b ({signal_2070, signal_1294}), .c ({signal_2117, signal_1277}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_768 ( .a ({signal_1870, signal_1325}), .b ({signal_1977, signal_659}), .c ({signal_2017, signal_661}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_769 ( .a ({signal_2184, signal_662}), .b ({signal_2020, signal_663}), .c ({signal_2196, signal_1278}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_770 ( .a ({signal_2176, signal_664}), .b ({signal_1972, signal_665}), .c ({signal_2184, signal_662}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_771 ( .a ({signal_1827, signal_880}), .b ({signal_1934, signal_1326}), .c ({signal_1972, signal_665}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_772 ( .a ({signal_2018, signal_1295}), .b ({signal_2148, signal_666}), .c ({signal_2176, signal_664}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_773 ( .a ({signal_1973, signal_667}), .b ({signal_1933, signal_668}), .c ({signal_2018, signal_1295}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_774 ( .a ({signal_1787, signal_901}), .b ({signal_1899, signal_1324}), .c ({signal_1933, signal_668}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_775 ( .a ({signal_1774, signal_883}), .b ({signal_1936, signal_1308}), .c ({signal_1973, signal_667}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_776 ( .a ({signal_2177, signal_669}), .b ({signal_1871, signal_1327}), .c ({signal_2185, signal_1279}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_777 ( .a ({signal_1936, signal_1308}), .b ({signal_2148, signal_666}), .c ({signal_2177, signal_669}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_778 ( .a ({signal_1772, signal_881}), .b ({signal_2118, signal_1292}), .c ({signal_2148, signal_666}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_779 ( .a ({signal_2069, signal_670}), .b ({signal_1828, signal_671}), .c ({signal_2118, signal_1292}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_780 ( .a ({signal_1827, signal_880}), .b ({signal_1788, signal_902}), .c ({signal_1828, signal_671}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_781 ( .a ({signal_2019, signal_1309}), .b ({signal_1870, signal_1325}), .c ({signal_2069, signal_670}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_782 ( .a ({signal_1974, signal_672}), .b ({signal_1868, signal_673}), .c ({signal_2019, signal_1309}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_783 ( .a ({signal_1837, signal_674}), .b ({signal_1773, signal_882}), .c ({signal_1868, signal_673}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_784 ( .a ({signal_1934, signal_1326}), .b ({signal_1801, signal_923}), .c ({signal_1974, signal_672}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_785 ( .a ({signal_1897, signal_675}), .b ({signal_1829, signal_676}), .c ({signal_1934, signal_1326}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_786 ( .a ({signal_1789, signal_903}), .b ({signal_1822, signal_900}), .c ({signal_1829, signal_676}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_787 ( .a ({signal_1835, signal_677}), .b ({signal_1869, signal_660}), .c ({signal_1897, signal_675}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_788 ( .a ({signal_1830, signal_678}), .b ({signal_1810, signal_941}), .c ({signal_1869, signal_660}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_789 ( .a ({signal_1800, signal_922}), .b ({signal_1812, signal_940}), .c ({signal_1830, signal_678}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_790 ( .a ({signal_2021, signal_679}), .b ({signal_2020, signal_663}), .c ({signal_2070, signal_1294}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_791 ( .a ({signal_1976, signal_1311}), .b ({signal_1936, signal_1308}), .c ({signal_2020, signal_663}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_792 ( .a ({signal_1975, signal_680}), .b ({signal_1831, signal_681}), .c ({signal_2021, signal_679}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_793 ( .a ({signal_1787, signal_901}), .b ({signal_1822, signal_900}), .c ({signal_1831, signal_681}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_794 ( .a ({signal_1937, signal_682}), .b ({signal_1773, signal_882}), .c ({signal_1975, signal_680}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_795 ( .a ({signal_1756, signal_683}), .b ({signal_1935, signal_684}), .c ({signal_1976, signal_1311}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_796 ( .a ({signal_1899, signal_1324}), .b ({signal_1827, signal_880}), .c ({signal_1935, signal_684}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_798 ( .a ({signal_1898, signal_685}), .b ({signal_1832, signal_686}), .c ({signal_1936, signal_1308}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_799 ( .a ({signal_1772, signal_881}), .b ({signal_1822, signal_900}), .c ({signal_1832, signal_686}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_800 ( .a ({signal_1870, signal_1325}), .b ({signal_1800, signal_922}), .c ({signal_1898, signal_685}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_801 ( .a ({signal_1757, signal_687}), .b ({signal_1833, signal_688}), .c ({signal_1870, signal_1325}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_802 ( .a ({signal_1758, signal_689}), .b ({signal_1812, signal_940}), .c ({signal_1833, signal_688}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_804 ( .a ({signal_1835, signal_677}), .b ({signal_1977, signal_659}), .c ({signal_2022, signal_1310}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_805 ( .a ({signal_1834, signal_690}), .b ({signal_1937, signal_682}), .c ({signal_1977, signal_659}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_806 ( .a ({signal_1899, signal_1324}), .b ({signal_1871, signal_1327}), .c ({signal_1937, signal_682}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_807 ( .a ({signal_1817, signal_920}), .b ({signal_1758, signal_689}), .c ({signal_1834, signal_690}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_809 ( .a ({signal_1827, signal_880}), .b ({signal_1774, signal_883}), .c ({signal_1835, signal_677}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_810 ( .a ({signal_1759, signal_691}), .b ({signal_1836, signal_692}), .c ({signal_1871, signal_1327}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_811 ( .a ({signal_1827, signal_880}), .b ({signal_1822, signal_900}), .c ({signal_1836, signal_692}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_813 ( .a ({signal_1872, signal_693}), .b ({signal_1772, signal_881}), .c ({signal_1899, signal_1324}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_814 ( .a ({signal_1837, signal_674}), .b ({signal_1811, signal_942}), .c ({signal_1872, signal_693}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_815 ( .a ({signal_1787, signal_901}), .b ({signal_1817, signal_920}), .c ({signal_1837, signal_674}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_816 ( .a ({signal_2071, signal_694}), .b ({signal_1938, signal_695}), .c ({signal_2119, signal_1272}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_817 ( .a ({signal_1903, signal_1320}), .b ({signal_1782, signal_894}), .c ({signal_1938, signal_695}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_818 ( .a ({signal_2023, signal_1289}), .b ({signal_2026, signal_1305}), .c ({signal_2071, signal_694}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_819 ( .a ({signal_1900, signal_696}), .b ({signal_1983, signal_697}), .c ({signal_2023, signal_1289}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_820 ( .a ({signal_1781, signal_893}), .b ({signal_1874, signal_698}), .c ({signal_1900, signal_696}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_821 ( .a ({signal_2024, signal_699}), .b ({signal_2073, signal_1290}), .c ({signal_2120, signal_1273}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_822 ( .a ({signal_1875, signal_1321}), .b ({signal_1983, signal_697}), .c ({signal_2024, signal_699}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_823 ( .a ({signal_2186, signal_700}), .b ({signal_2027, signal_701}), .c ({signal_2197, signal_1274}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_824 ( .a ({signal_2178, signal_702}), .b ({signal_1978, signal_703}), .c ({signal_2186, signal_700}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_825 ( .a ({signal_1824, signal_892}), .b ({signal_1940, signal_1322}), .c ({signal_1978, signal_703}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_826 ( .a ({signal_2025, signal_1291}), .b ({signal_2149, signal_704}), .c ({signal_2178, signal_702}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_827 ( .a ({signal_1979, signal_705}), .b ({signal_1939, signal_706}), .c ({signal_2025, signal_1291}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_828 ( .a ({signal_1784, signal_897}), .b ({signal_1903, signal_1320}), .c ({signal_1939, signal_706}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_829 ( .a ({signal_1783, signal_895}), .b ({signal_1942, signal_1304}), .c ({signal_1979, signal_705}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_830 ( .a ({signal_2179, signal_707}), .b ({signal_1876, signal_1323}), .c ({signal_2187, signal_1275}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_831 ( .a ({signal_1942, signal_1304}), .b ({signal_2149, signal_704}), .c ({signal_2179, signal_707}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_832 ( .a ({signal_1781, signal_893}), .b ({signal_2121, signal_1288}), .c ({signal_2149, signal_704}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_833 ( .a ({signal_2072, signal_708}), .b ({signal_1838, signal_709}), .c ({signal_2121, signal_1288}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_834 ( .a ({signal_1824, signal_892}), .b ({signal_1785, signal_898}), .c ({signal_1838, signal_709}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_835 ( .a ({signal_2026, signal_1305}), .b ({signal_1875, signal_1321}), .c ({signal_2072, signal_708}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_836 ( .a ({signal_1980, signal_710}), .b ({signal_1873, signal_711}), .c ({signal_2026, signal_1305}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_837 ( .a ({signal_1847, signal_712}), .b ({signal_1782, signal_894}), .c ({signal_1873, signal_711}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_838 ( .a ({signal_1940, signal_1322}), .b ({signal_1799, signal_919}), .c ({signal_1980, signal_710}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_839 ( .a ({signal_1901, signal_713}), .b ({signal_1839, signal_714}), .c ({signal_1940, signal_1322}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_840 ( .a ({signal_1786, signal_899}), .b ({signal_1823, signal_896}), .c ({signal_1839, signal_714}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_841 ( .a ({signal_1845, signal_715}), .b ({signal_1874, signal_698}), .c ({signal_1901, signal_713}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_842 ( .a ({signal_1840, signal_716}), .b ({signal_1808, signal_937}), .c ({signal_1874, signal_698}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_843 ( .a ({signal_1798, signal_918}), .b ({signal_1813, signal_936}), .c ({signal_1840, signal_716}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_844 ( .a ({signal_2028, signal_717}), .b ({signal_2027, signal_701}), .c ({signal_2073, signal_1290}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_845 ( .a ({signal_1982, signal_1307}), .b ({signal_1942, signal_1304}), .c ({signal_2027, signal_701}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_846 ( .a ({signal_1981, signal_718}), .b ({signal_1841, signal_719}), .c ({signal_2028, signal_717}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_847 ( .a ({signal_1784, signal_897}), .b ({signal_1823, signal_896}), .c ({signal_1841, signal_719}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_848 ( .a ({signal_1943, signal_720}), .b ({signal_1782, signal_894}), .c ({signal_1981, signal_718}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_849 ( .a ({signal_1760, signal_721}), .b ({signal_1941, signal_722}), .c ({signal_1982, signal_1307}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_850 ( .a ({signal_1903, signal_1320}), .b ({signal_1824, signal_892}), .c ({signal_1941, signal_722}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_852 ( .a ({signal_1902, signal_723}), .b ({signal_1842, signal_724}), .c ({signal_1942, signal_1304}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_853 ( .a ({signal_1781, signal_893}), .b ({signal_1823, signal_896}), .c ({signal_1842, signal_724}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_854 ( .a ({signal_1875, signal_1321}), .b ({signal_1798, signal_918}), .c ({signal_1902, signal_723}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_855 ( .a ({signal_1761, signal_725}), .b ({signal_1843, signal_726}), .c ({signal_1875, signal_1321}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_856 ( .a ({signal_1762, signal_727}), .b ({signal_1813, signal_936}), .c ({signal_1843, signal_726}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_858 ( .a ({signal_1845, signal_715}), .b ({signal_1983, signal_697}), .c ({signal_2029, signal_1306}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_859 ( .a ({signal_1844, signal_728}), .b ({signal_1943, signal_720}), .c ({signal_1983, signal_697}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_860 ( .a ({signal_1903, signal_1320}), .b ({signal_1876, signal_1323}), .c ({signal_1943, signal_720}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_861 ( .a ({signal_1818, signal_916}), .b ({signal_1762, signal_727}), .c ({signal_1844, signal_728}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_863 ( .a ({signal_1824, signal_892}), .b ({signal_1783, signal_895}), .c ({signal_1845, signal_715}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_864 ( .a ({signal_1763, signal_729}), .b ({signal_1846, signal_730}), .c ({signal_1876, signal_1323}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_865 ( .a ({signal_1824, signal_892}), .b ({signal_1823, signal_896}), .c ({signal_1846, signal_730}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_867 ( .a ({signal_1877, signal_731}), .b ({signal_1781, signal_893}), .c ({signal_1903, signal_1320}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_868 ( .a ({signal_1847, signal_712}), .b ({signal_1809, signal_938}), .c ({signal_1877, signal_731}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_869 ( .a ({signal_1784, signal_897}), .b ({signal_1818, signal_916}), .c ({signal_1847, signal_712}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_870 ( .a ({signal_2074, signal_732}), .b ({signal_1944, signal_733}), .c ({signal_2122, signal_1268}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_871 ( .a ({signal_1907, signal_1316}), .b ({signal_1779, signal_890}), .c ({signal_1944, signal_733}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_872 ( .a ({signal_2030, signal_1285}), .b ({signal_2033, signal_1301}), .c ({signal_2074, signal_732}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_873 ( .a ({signal_1904, signal_734}), .b ({signal_1989, signal_735}), .c ({signal_2030, signal_1285}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_874 ( .a ({signal_1778, signal_889}), .b ({signal_1879, signal_736}), .c ({signal_1904, signal_734}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_875 ( .a ({signal_2031, signal_737}), .b ({signal_2076, signal_1286}), .c ({signal_2123, signal_1269}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_876 ( .a ({signal_1880, signal_1317}), .b ({signal_1989, signal_735}), .c ({signal_2031, signal_737}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_877 ( .a ({signal_2188, signal_738}), .b ({signal_2034, signal_739}), .c ({signal_2198, signal_1270}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_878 ( .a ({signal_2180, signal_740}), .b ({signal_1984, signal_741}), .c ({signal_2188, signal_738}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_879 ( .a ({signal_1825, signal_888}), .b ({signal_1946, signal_1318}), .c ({signal_1984, signal_741}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_880 ( .a ({signal_2032, signal_1287}), .b ({signal_2150, signal_742}), .c ({signal_2180, signal_740}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_881 ( .a ({signal_1985, signal_743}), .b ({signal_1945, signal_744}), .c ({signal_2032, signal_1287}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_882 ( .a ({signal_1793, signal_909}), .b ({signal_1907, signal_1316}), .c ({signal_1945, signal_744}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_883 ( .a ({signal_1780, signal_891}), .b ({signal_1948, signal_1300}), .c ({signal_1985, signal_743}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_884 ( .a ({signal_2181, signal_745}), .b ({signal_1881, signal_1319}), .c ({signal_2189, signal_1271}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_885 ( .a ({signal_1948, signal_1300}), .b ({signal_2150, signal_742}), .c ({signal_2181, signal_745}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_886 ( .a ({signal_1778, signal_889}), .b ({signal_2124, signal_1284}), .c ({signal_2150, signal_742}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_887 ( .a ({signal_2075, signal_746}), .b ({signal_1848, signal_747}), .c ({signal_2124, signal_1284}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_888 ( .a ({signal_1825, signal_888}), .b ({signal_1794, signal_910}), .c ({signal_1848, signal_747}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_889 ( .a ({signal_2033, signal_1301}), .b ({signal_1880, signal_1317}), .c ({signal_2075, signal_746}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_890 ( .a ({signal_1986, signal_748}), .b ({signal_1878, signal_749}), .c ({signal_2033, signal_1301}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_891 ( .a ({signal_1857, signal_750}), .b ({signal_1779, signal_890}), .c ({signal_1878, signal_749}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_892 ( .a ({signal_1946, signal_1318}), .b ({signal_1797, signal_915}), .c ({signal_1986, signal_748}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_893 ( .a ({signal_1905, signal_751}), .b ({signal_1849, signal_752}), .c ({signal_1946, signal_1318}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_894 ( .a ({signal_1795, signal_911}), .b ({signal_1820, signal_908}), .c ({signal_1849, signal_752}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_895 ( .a ({signal_1855, signal_753}), .b ({signal_1879, signal_736}), .c ({signal_1905, signal_751}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_896 ( .a ({signal_1850, signal_754}), .b ({signal_1806, signal_933}), .c ({signal_1879, signal_736}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_897 ( .a ({signal_1796, signal_914}), .b ({signal_1814, signal_932}), .c ({signal_1850, signal_754}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_898 ( .a ({signal_2035, signal_755}), .b ({signal_2034, signal_739}), .c ({signal_2076, signal_1286}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_899 ( .a ({signal_1988, signal_1303}), .b ({signal_1948, signal_1300}), .c ({signal_2034, signal_739}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_900 ( .a ({signal_1987, signal_756}), .b ({signal_1851, signal_757}), .c ({signal_2035, signal_755}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_901 ( .a ({signal_1793, signal_909}), .b ({signal_1820, signal_908}), .c ({signal_1851, signal_757}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_902 ( .a ({signal_1949, signal_758}), .b ({signal_1779, signal_890}), .c ({signal_1987, signal_756}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_903 ( .a ({signal_1764, signal_759}), .b ({signal_1947, signal_760}), .c ({signal_1988, signal_1303}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_904 ( .a ({signal_1907, signal_1316}), .b ({signal_1825, signal_888}), .c ({signal_1947, signal_760}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_906 ( .a ({signal_1906, signal_761}), .b ({signal_1852, signal_762}), .c ({signal_1948, signal_1300}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_907 ( .a ({signal_1778, signal_889}), .b ({signal_1820, signal_908}), .c ({signal_1852, signal_762}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_908 ( .a ({signal_1880, signal_1317}), .b ({signal_1796, signal_914}), .c ({signal_1906, signal_761}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_909 ( .a ({signal_1765, signal_763}), .b ({signal_1853, signal_764}), .c ({signal_1880, signal_1317}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_910 ( .a ({signal_1766, signal_765}), .b ({signal_1814, signal_932}), .c ({signal_1853, signal_764}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_912 ( .a ({signal_1855, signal_753}), .b ({signal_1989, signal_735}), .c ({signal_2036, signal_1302}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_913 ( .a ({signal_1854, signal_766}), .b ({signal_1949, signal_758}), .c ({signal_1989, signal_735}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_914 ( .a ({signal_1907, signal_1316}), .b ({signal_1881, signal_1319}), .c ({signal_1949, signal_758}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_915 ( .a ({signal_1819, signal_912}), .b ({signal_1766, signal_765}), .c ({signal_1854, signal_766}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_917 ( .a ({signal_1825, signal_888}), .b ({signal_1780, signal_891}), .c ({signal_1855, signal_753}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_918 ( .a ({signal_1767, signal_767}), .b ({signal_1856, signal_768}), .c ({signal_1881, signal_1319}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_919 ( .a ({signal_1825, signal_888}), .b ({signal_1820, signal_908}), .c ({signal_1856, signal_768}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_921 ( .a ({signal_1882, signal_769}), .b ({signal_1778, signal_889}), .c ({signal_1907, signal_1316}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_922 ( .a ({signal_1857, signal_750}), .b ({signal_1807, signal_934}), .c ({signal_1882, signal_769}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_923 ( .a ({signal_1793, signal_909}), .b ({signal_1819, signal_912}), .c ({signal_1857, signal_750}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_924 ( .a ({signal_2077, signal_770}), .b ({signal_1950, signal_771}), .c ({signal_2125, signal_1264}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_925 ( .a ({signal_1911, signal_1312}), .b ({signal_1776, signal_886}), .c ({signal_1950, signal_771}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_926 ( .a ({signal_2037, signal_1281}), .b ({signal_2040, signal_1297}), .c ({signal_2077, signal_770}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_927 ( .a ({signal_1908, signal_772}), .b ({signal_1995, signal_773}), .c ({signal_2037, signal_1281}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_928 ( .a ({signal_1775, signal_885}), .b ({signal_1884, signal_774}), .c ({signal_1908, signal_772}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_929 ( .a ({signal_2038, signal_775}), .b ({signal_2079, signal_1282}), .c ({signal_2126, signal_1265}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_930 ( .a ({signal_1885, signal_1313}), .b ({signal_1995, signal_773}), .c ({signal_2038, signal_775}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_931 ( .a ({signal_2190, signal_776}), .b ({signal_2041, signal_777}), .c ({signal_2199, signal_1266}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_932 ( .a ({signal_2182, signal_778}), .b ({signal_1990, signal_779}), .c ({signal_2190, signal_776}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_933 ( .a ({signal_1826, signal_884}), .b ({signal_1952, signal_1314}), .c ({signal_1990, signal_779}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_934 ( .a ({signal_2039, signal_1283}), .b ({signal_2151, signal_780}), .c ({signal_2182, signal_778}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_935 ( .a ({signal_1991, signal_781}), .b ({signal_1951, signal_782}), .c ({signal_2039, signal_1283}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_936 ( .a ({signal_1790, signal_905}), .b ({signal_1911, signal_1312}), .c ({signal_1951, signal_782}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_937 ( .a ({signal_1777, signal_887}), .b ({signal_1954, signal_1296}), .c ({signal_1991, signal_781}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_938 ( .a ({signal_2183, signal_783}), .b ({signal_1886, signal_1315}), .c ({signal_2191, signal_1267}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_939 ( .a ({signal_1954, signal_1296}), .b ({signal_2151, signal_780}), .c ({signal_2183, signal_783}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_940 ( .a ({signal_1775, signal_885}), .b ({signal_2127, signal_1280}), .c ({signal_2151, signal_780}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_941 ( .a ({signal_2078, signal_784}), .b ({signal_1858, signal_785}), .c ({signal_2127, signal_1280}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_942 ( .a ({signal_1826, signal_884}), .b ({signal_1791, signal_906}), .c ({signal_1858, signal_785}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_943 ( .a ({signal_2040, signal_1297}), .b ({signal_1885, signal_1313}), .c ({signal_2078, signal_784}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_944 ( .a ({signal_1992, signal_786}), .b ({signal_1883, signal_787}), .c ({signal_2040, signal_1297}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_945 ( .a ({signal_1867, signal_788}), .b ({signal_1776, signal_886}), .c ({signal_1883, signal_787}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_946 ( .a ({signal_1952, signal_1314}), .b ({signal_1803, signal_927}), .c ({signal_1992, signal_786}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_947 ( .a ({signal_1909, signal_789}), .b ({signal_1859, signal_790}), .c ({signal_1952, signal_1314}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_948 ( .a ({signal_1792, signal_907}), .b ({signal_1821, signal_904}), .c ({signal_1859, signal_790}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_949 ( .a ({signal_1865, signal_791}), .b ({signal_1884, signal_774}), .c ({signal_1909, signal_789}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_950 ( .a ({signal_1860, signal_792}), .b ({signal_1804, signal_929}), .c ({signal_1884, signal_774}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_951 ( .a ({signal_1802, signal_926}), .b ({signal_1815, signal_928}), .c ({signal_1860, signal_792}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_952 ( .a ({signal_2042, signal_793}), .b ({signal_2041, signal_777}), .c ({signal_2079, signal_1282}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_953 ( .a ({signal_1994, signal_1299}), .b ({signal_1954, signal_1296}), .c ({signal_2041, signal_777}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_954 ( .a ({signal_1993, signal_794}), .b ({signal_1861, signal_795}), .c ({signal_2042, signal_793}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_955 ( .a ({signal_1790, signal_905}), .b ({signal_1821, signal_904}), .c ({signal_1861, signal_795}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_956 ( .a ({signal_1955, signal_796}), .b ({signal_1776, signal_886}), .c ({signal_1993, signal_794}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_957 ( .a ({signal_1768, signal_797}), .b ({signal_1953, signal_798}), .c ({signal_1994, signal_1299}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_958 ( .a ({signal_1911, signal_1312}), .b ({signal_1826, signal_884}), .c ({signal_1953, signal_798}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_960 ( .a ({signal_1910, signal_799}), .b ({signal_1862, signal_800}), .c ({signal_1954, signal_1296}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_961 ( .a ({signal_1775, signal_885}), .b ({signal_1821, signal_904}), .c ({signal_1862, signal_800}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_962 ( .a ({signal_1885, signal_1313}), .b ({signal_1802, signal_926}), .c ({signal_1910, signal_799}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_963 ( .a ({signal_1769, signal_801}), .b ({signal_1863, signal_802}), .c ({signal_1885, signal_1313}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_964 ( .a ({signal_1770, signal_803}), .b ({signal_1815, signal_928}), .c ({signal_1863, signal_802}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_966 ( .a ({signal_1865, signal_791}), .b ({signal_1995, signal_773}), .c ({signal_2043, signal_1298}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_967 ( .a ({signal_1864, signal_804}), .b ({signal_1955, signal_796}), .c ({signal_1995, signal_773}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_968 ( .a ({signal_1911, signal_1312}), .b ({signal_1886, signal_1315}), .c ({signal_1955, signal_796}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_969 ( .a ({signal_1816, signal_924}), .b ({signal_1770, signal_803}), .c ({signal_1864, signal_804}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_971 ( .a ({signal_1826, signal_884}), .b ({signal_1777, signal_887}), .c ({signal_1865, signal_791}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_972 ( .a ({signal_1771, signal_805}), .b ({signal_1866, signal_806}), .c ({signal_1886, signal_1315}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_973 ( .a ({signal_1826, signal_884}), .b ({signal_1821, signal_904}), .c ({signal_1866, signal_806}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_975 ( .a ({signal_1887, signal_807}), .b ({signal_1775, signal_885}), .c ({signal_1911, signal_1312}) ) ;
    xnor_GHPC #(.low_latency(0), .pipeline(1)) cell_976 ( .a ({signal_1867, signal_788}), .b ({signal_1805, signal_930}), .c ({signal_1887, signal_807}) ) ;
    xor_GHPC #(.low_latency(0), .pipeline(1)) cell_977 ( .a ({signal_1790, signal_905}), .b ({signal_1816, signal_924}), .c ({signal_1867, signal_788}) ) ;
    LED_step2_ANF #(.low_latency(0), .pipeline(1)) cell_1128 ( .in0 ({signal_999, signal_998, signal_997, signal_996, signal_995, signal_994, signal_993, signal_992, signal_991, signal_990, signal_989, signal_988, signal_987, signal_986, signal_985, signal_984, signal_983, signal_982, signal_981, signal_980, signal_979, signal_978, signal_977, signal_976, signal_975, signal_974, signal_973, signal_972, signal_971, signal_970, signal_969, signal_968, signal_967, signal_966, signal_965, signal_964, signal_963, signal_962, signal_961, signal_960, signal_959, signal_958, signal_957, signal_956, signal_955, signal_954, signal_953, signal_952, signal_951, signal_950, signal_949, signal_948, signal_947, signal_946, signal_945, signal_944, signal_1007, signal_1006, signal_1005, signal_1004, signal_1003, signal_1002, signal_1001, signal_1000}), .in1 ({signal_1672, signal_1673, signal_1674, signal_1675, signal_1676, signal_1677, signal_1678, signal_1679, signal_1664, signal_1739, signal_1738, signal_1663, signal_1736, signal_1735, signal_1662, signal_1684, signal_1551, signal_1685, signal_1552, signal_1686, signal_1655, signal_1687, signal_1688, signal_1689, signal_1720, signal_1733, signal_1719, signal_1718, signal_1717, signal_1732, signal_1731, signal_1660, signal_1693, signal_1694, signal_1695, signal_1696, signal_1697, signal_1698, signal_1699, signal_1700, signal_1730, signal_1729, signal_1727, signal_1726, signal_1725, signal_1724, signal_1723, signal_1708, signal_1709, signal_1710, signal_1711, signal_1712, signal_1713, signal_1714, signal_1715, signal_1716, signal_1665, signal_1737, signal_1734, signal_1661, signal_1728, signal_1722, signal_1721, signal_1671}), .clk (CLK), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_942, signal_941, signal_938, signal_937, signal_934, signal_933, signal_930, signal_929, signal_927, signal_926, signal_923, signal_922, signal_919, signal_918, signal_915, signal_914, signal_911, signal_910, signal_909, signal_907, signal_906, signal_905, signal_903, signal_902, signal_901, signal_899, signal_898, signal_897, signal_895, signal_894, signal_893, signal_891, signal_890, signal_889, signal_887, signal_886, signal_885, signal_883, signal_882, signal_881, signal_805, signal_803, signal_801, signal_797, signal_767, signal_765, signal_763, signal_759, signal_729, signal_727, signal_725, signal_721, signal_691, signal_689, signal_687, signal_683, signal_641, signal_622, signal_603, signal_584, signal_565, signal_546, signal_527, signal_508, signal_489, signal_470, signal_451, signal_432, signal_413, signal_394, signal_375, signal_356}), .out1 ({signal_1811, signal_1810, signal_1809, signal_1808, signal_1807, signal_1806, signal_1805, signal_1804, signal_1803, signal_1802, signal_1801, signal_1800, signal_1799, signal_1798, signal_1797, signal_1796, signal_1795, signal_1794, signal_1793, signal_1792, signal_1791, signal_1790, signal_1789, signal_1788, signal_1787, signal_1786, signal_1785, signal_1784, signal_1783, signal_1782, signal_1781, signal_1780, signal_1779, signal_1778, signal_1777, signal_1776, signal_1775, signal_1774, signal_1773, signal_1772, signal_1771, signal_1770, signal_1769, signal_1768, signal_1767, signal_1766, signal_1765, signal_1764, signal_1763, signal_1762, signal_1761, signal_1760, signal_1759, signal_1758, signal_1757, signal_1756, signal_1755, signal_1754, signal_1753, signal_1752, signal_1751, signal_1750, signal_1749, signal_1748, signal_1747, signal_1746, signal_1745, signal_1744, signal_1743, signal_1742, signal_1741, signal_1740}) ) ;
    buf_clk cell_1130 ( .C (CLK), .D (signal_2284), .Q (signal_2285) ) ;
    buf_clk cell_1132 ( .C (CLK), .D (signal_2286), .Q (signal_2287) ) ;
    buf_clk cell_1134 ( .C (CLK), .D (signal_2288), .Q (signal_2289) ) ;
    buf_clk cell_1136 ( .C (CLK), .D (signal_2290), .Q (signal_2291) ) ;
    buf_clk cell_1138 ( .C (CLK), .D (signal_2292), .Q (signal_2293) ) ;
    buf_clk cell_1140 ( .C (CLK), .D (signal_2294), .Q (signal_2295) ) ;
    buf_clk cell_1142 ( .C (CLK), .D (signal_2296), .Q (signal_2297) ) ;
    buf_clk cell_1144 ( .C (CLK), .D (signal_2298), .Q (signal_2299) ) ;
    buf_clk cell_1146 ( .C (CLK), .D (signal_2300), .Q (signal_2301) ) ;
    buf_clk cell_1148 ( .C (CLK), .D (signal_2302), .Q (signal_2303) ) ;
    buf_clk cell_1150 ( .C (CLK), .D (signal_2304), .Q (signal_2305) ) ;
    buf_clk cell_1152 ( .C (CLK), .D (signal_2306), .Q (signal_2307) ) ;
    buf_clk cell_1154 ( .C (CLK), .D (signal_2308), .Q (signal_2309) ) ;
    buf_clk cell_1156 ( .C (CLK), .D (signal_2310), .Q (signal_2311) ) ;
    buf_clk cell_1158 ( .C (CLK), .D (signal_2312), .Q (signal_2313) ) ;
    buf_clk cell_1160 ( .C (CLK), .D (signal_2314), .Q (signal_2315) ) ;
    buf_clk cell_1162 ( .C (CLK), .D (signal_2316), .Q (signal_2317) ) ;
    buf_clk cell_1164 ( .C (CLK), .D (signal_2318), .Q (signal_2319) ) ;
    buf_clk cell_1166 ( .C (CLK), .D (signal_2320), .Q (signal_2321) ) ;
    buf_clk cell_1168 ( .C (CLK), .D (signal_2322), .Q (signal_2323) ) ;
    buf_clk cell_1170 ( .C (CLK), .D (signal_2324), .Q (signal_2325) ) ;
    buf_clk cell_1172 ( .C (CLK), .D (signal_2326), .Q (signal_2327) ) ;
    buf_clk cell_1174 ( .C (CLK), .D (signal_2328), .Q (signal_2329) ) ;
    buf_clk cell_1176 ( .C (CLK), .D (signal_2330), .Q (signal_2331) ) ;
    buf_clk cell_1178 ( .C (CLK), .D (signal_2332), .Q (signal_2333) ) ;
    buf_clk cell_1180 ( .C (CLK), .D (signal_2334), .Q (signal_2335) ) ;
    buf_clk cell_1182 ( .C (CLK), .D (signal_2336), .Q (signal_2337) ) ;
    buf_clk cell_1184 ( .C (CLK), .D (signal_2338), .Q (signal_2339) ) ;
    buf_clk cell_1186 ( .C (CLK), .D (signal_2340), .Q (signal_2341) ) ;
    buf_clk cell_1188 ( .C (CLK), .D (signal_2342), .Q (signal_2343) ) ;
    buf_clk cell_1190 ( .C (CLK), .D (signal_2344), .Q (signal_2345) ) ;
    buf_clk cell_1192 ( .C (CLK), .D (signal_2346), .Q (signal_2347) ) ;
    buf_clk cell_1194 ( .C (CLK), .D (signal_2348), .Q (signal_2349) ) ;
    buf_clk cell_1196 ( .C (CLK), .D (signal_2350), .Q (signal_2351) ) ;
    buf_clk cell_1198 ( .C (CLK), .D (signal_2352), .Q (signal_2353) ) ;
    buf_clk cell_1200 ( .C (CLK), .D (signal_2354), .Q (signal_2355) ) ;
    buf_clk cell_1202 ( .C (CLK), .D (signal_2356), .Q (signal_2357) ) ;
    buf_clk cell_1204 ( .C (CLK), .D (signal_2358), .Q (signal_2359) ) ;
    buf_clk cell_1206 ( .C (CLK), .D (signal_2360), .Q (signal_2361) ) ;
    buf_clk cell_1208 ( .C (CLK), .D (signal_2362), .Q (signal_2363) ) ;
    buf_clk cell_1210 ( .C (CLK), .D (signal_2364), .Q (signal_2365) ) ;
    buf_clk cell_1212 ( .C (CLK), .D (signal_2366), .Q (signal_2367) ) ;
    buf_clk cell_1214 ( .C (CLK), .D (signal_2368), .Q (signal_2369) ) ;
    buf_clk cell_1216 ( .C (CLK), .D (signal_2370), .Q (signal_2371) ) ;
    buf_clk cell_1218 ( .C (CLK), .D (signal_2372), .Q (signal_2373) ) ;
    buf_clk cell_1220 ( .C (CLK), .D (signal_2374), .Q (signal_2375) ) ;
    buf_clk cell_1222 ( .C (CLK), .D (signal_2376), .Q (signal_2377) ) ;
    buf_clk cell_1224 ( .C (CLK), .D (signal_2378), .Q (signal_2379) ) ;
    buf_clk cell_1226 ( .C (CLK), .D (signal_2380), .Q (signal_2381) ) ;
    buf_clk cell_1228 ( .C (CLK), .D (signal_2382), .Q (signal_2383) ) ;
    buf_clk cell_1230 ( .C (CLK), .D (signal_2384), .Q (signal_2385) ) ;
    buf_clk cell_1232 ( .C (CLK), .D (signal_2386), .Q (signal_2387) ) ;
    buf_clk cell_1234 ( .C (CLK), .D (signal_2388), .Q (signal_2389) ) ;
    buf_clk cell_1236 ( .C (CLK), .D (signal_2390), .Q (signal_2391) ) ;
    buf_clk cell_1238 ( .C (CLK), .D (signal_2392), .Q (signal_2393) ) ;
    buf_clk cell_1240 ( .C (CLK), .D (signal_2394), .Q (signal_2395) ) ;
    buf_clk cell_1242 ( .C (CLK), .D (signal_2396), .Q (signal_2397) ) ;
    buf_clk cell_1244 ( .C (CLK), .D (signal_2398), .Q (signal_2399) ) ;
    buf_clk cell_1246 ( .C (CLK), .D (signal_2400), .Q (signal_2401) ) ;
    buf_clk cell_1248 ( .C (CLK), .D (signal_2402), .Q (signal_2403) ) ;
    buf_clk cell_1250 ( .C (CLK), .D (signal_2404), .Q (signal_2405) ) ;
    buf_clk cell_1252 ( .C (CLK), .D (signal_2406), .Q (signal_2407) ) ;
    buf_clk cell_1254 ( .C (CLK), .D (signal_2408), .Q (signal_2409) ) ;
    buf_clk cell_1256 ( .C (CLK), .D (signal_2410), .Q (signal_2411) ) ;
    buf_clk cell_1258 ( .C (CLK), .D (signal_2412), .Q (signal_2413) ) ;
    buf_clk cell_1260 ( .C (CLK), .D (signal_2414), .Q (signal_2415) ) ;
    buf_clk cell_1262 ( .C (CLK), .D (signal_2416), .Q (signal_2417) ) ;
    buf_clk cell_1264 ( .C (CLK), .D (signal_2418), .Q (signal_2419) ) ;
    buf_clk cell_1266 ( .C (CLK), .D (signal_2420), .Q (signal_2421) ) ;
    buf_clk cell_1268 ( .C (CLK), .D (signal_2422), .Q (signal_2423) ) ;
    buf_clk cell_1270 ( .C (CLK), .D (signal_2424), .Q (signal_2425) ) ;
    buf_clk cell_1272 ( .C (CLK), .D (signal_2426), .Q (signal_2427) ) ;
    buf_clk cell_1274 ( .C (CLK), .D (signal_2428), .Q (signal_2429) ) ;
    buf_clk cell_1276 ( .C (CLK), .D (signal_2430), .Q (signal_2431) ) ;
    buf_clk cell_1278 ( .C (CLK), .D (signal_2432), .Q (signal_2433) ) ;
    buf_clk cell_1280 ( .C (CLK), .D (signal_2434), .Q (signal_2435) ) ;
    buf_clk cell_1282 ( .C (CLK), .D (signal_2436), .Q (signal_2437) ) ;
    buf_clk cell_1284 ( .C (CLK), .D (signal_2438), .Q (signal_2439) ) ;
    buf_clk cell_1286 ( .C (CLK), .D (signal_2440), .Q (signal_2441) ) ;
    buf_clk cell_1288 ( .C (CLK), .D (signal_2442), .Q (signal_2443) ) ;
    buf_clk cell_1290 ( .C (CLK), .D (signal_2444), .Q (signal_2445) ) ;
    buf_clk cell_1292 ( .C (CLK), .D (signal_2446), .Q (signal_2447) ) ;
    buf_clk cell_1294 ( .C (CLK), .D (signal_2448), .Q (signal_2449) ) ;
    buf_clk cell_1296 ( .C (CLK), .D (signal_2450), .Q (signal_2451) ) ;
    buf_clk cell_1298 ( .C (CLK), .D (signal_2452), .Q (signal_2453) ) ;
    buf_clk cell_1300 ( .C (CLK), .D (signal_2454), .Q (signal_2455) ) ;
    buf_clk cell_1302 ( .C (CLK), .D (signal_2456), .Q (signal_2457) ) ;
    buf_clk cell_1304 ( .C (CLK), .D (signal_2458), .Q (signal_2459) ) ;
    buf_clk cell_1306 ( .C (CLK), .D (signal_2460), .Q (signal_2461) ) ;
    buf_clk cell_1308 ( .C (CLK), .D (signal_2462), .Q (signal_2463) ) ;
    buf_clk cell_1310 ( .C (CLK), .D (signal_2464), .Q (signal_2465) ) ;
    buf_clk cell_1312 ( .C (CLK), .D (signal_2466), .Q (signal_2467) ) ;
    buf_clk cell_1314 ( .C (CLK), .D (signal_2468), .Q (signal_2469) ) ;
    buf_clk cell_1316 ( .C (CLK), .D (signal_2470), .Q (signal_2471) ) ;
    buf_clk cell_1318 ( .C (CLK), .D (signal_2472), .Q (signal_2473) ) ;
    buf_clk cell_1320 ( .C (CLK), .D (signal_2474), .Q (signal_2475) ) ;
    buf_clk cell_1322 ( .C (CLK), .D (signal_2476), .Q (signal_2477) ) ;
    buf_clk cell_1324 ( .C (CLK), .D (signal_2478), .Q (signal_2479) ) ;
    buf_clk cell_1326 ( .C (CLK), .D (signal_2480), .Q (signal_2481) ) ;
    buf_clk cell_1328 ( .C (CLK), .D (signal_2482), .Q (signal_2483) ) ;
    buf_clk cell_1330 ( .C (CLK), .D (signal_2484), .Q (signal_2485) ) ;
    buf_clk cell_1332 ( .C (CLK), .D (signal_2486), .Q (signal_2487) ) ;
    buf_clk cell_1334 ( .C (CLK), .D (signal_2488), .Q (signal_2489) ) ;
    buf_clk cell_1336 ( .C (CLK), .D (signal_2490), .Q (signal_2491) ) ;
    buf_clk cell_1338 ( .C (CLK), .D (signal_2492), .Q (signal_2493) ) ;
    buf_clk cell_1340 ( .C (CLK), .D (signal_2494), .Q (signal_2495) ) ;
    buf_clk cell_1342 ( .C (CLK), .D (signal_2496), .Q (signal_2497) ) ;
    buf_clk cell_1344 ( .C (CLK), .D (signal_2498), .Q (signal_2499) ) ;
    buf_clk cell_1346 ( .C (CLK), .D (signal_2500), .Q (signal_2501) ) ;
    buf_clk cell_1348 ( .C (CLK), .D (signal_2502), .Q (signal_2503) ) ;
    buf_clk cell_1350 ( .C (CLK), .D (signal_2504), .Q (signal_2505) ) ;
    buf_clk cell_1352 ( .C (CLK), .D (signal_2506), .Q (signal_2507) ) ;
    buf_clk cell_1354 ( .C (CLK), .D (signal_2508), .Q (signal_2509) ) ;
    buf_clk cell_1356 ( .C (CLK), .D (signal_2510), .Q (signal_2511) ) ;
    buf_clk cell_1358 ( .C (CLK), .D (signal_2512), .Q (signal_2513) ) ;
    buf_clk cell_1360 ( .C (CLK), .D (signal_2514), .Q (signal_2515) ) ;
    buf_clk cell_1362 ( .C (CLK), .D (signal_2516), .Q (signal_2517) ) ;
    buf_clk cell_1364 ( .C (CLK), .D (signal_2518), .Q (signal_2519) ) ;
    buf_clk cell_1366 ( .C (CLK), .D (signal_2520), .Q (signal_2521) ) ;
    buf_clk cell_1368 ( .C (CLK), .D (signal_2522), .Q (signal_2523) ) ;
    buf_clk cell_1370 ( .C (CLK), .D (signal_2524), .Q (signal_2525) ) ;
    buf_clk cell_1372 ( .C (CLK), .D (signal_2526), .Q (signal_2527) ) ;
    buf_clk cell_1374 ( .C (CLK), .D (signal_2528), .Q (signal_2529) ) ;
    buf_clk cell_1376 ( .C (CLK), .D (signal_2530), .Q (signal_2531) ) ;
    buf_clk cell_1378 ( .C (CLK), .D (signal_2532), .Q (signal_2533) ) ;
    buf_clk cell_1380 ( .C (CLK), .D (signal_2534), .Q (signal_2535) ) ;
    buf_clk cell_1382 ( .C (CLK), .D (signal_2536), .Q (signal_2537) ) ;
    buf_clk cell_1384 ( .C (CLK), .D (signal_2538), .Q (signal_2539) ) ;
    buf_clk cell_1386 ( .C (CLK), .D (signal_2540), .Q (signal_2541) ) ;
    buf_clk cell_1388 ( .C (CLK), .D (signal_2542), .Q (signal_2543) ) ;
    buf_clk cell_1390 ( .C (CLK), .D (signal_2544), .Q (signal_2545) ) ;
    buf_clk cell_1392 ( .C (CLK), .D (signal_2546), .Q (signal_2547) ) ;
    buf_clk cell_1394 ( .C (CLK), .D (signal_2548), .Q (signal_2549) ) ;
    buf_clk cell_1396 ( .C (CLK), .D (signal_2550), .Q (signal_2551) ) ;
    buf_clk cell_1398 ( .C (CLK), .D (signal_2552), .Q (signal_2553) ) ;
    buf_clk cell_1400 ( .C (CLK), .D (signal_2554), .Q (signal_2555) ) ;
    buf_clk cell_1402 ( .C (CLK), .D (signal_2556), .Q (signal_2557) ) ;
    buf_clk cell_1404 ( .C (CLK), .D (signal_2558), .Q (signal_2559) ) ;
    buf_clk cell_1406 ( .C (CLK), .D (signal_2560), .Q (signal_2561) ) ;
    buf_clk cell_1408 ( .C (CLK), .D (signal_2562), .Q (signal_2563) ) ;
    buf_clk cell_1410 ( .C (CLK), .D (signal_2564), .Q (signal_2565) ) ;
    buf_clk cell_1412 ( .C (CLK), .D (signal_2566), .Q (signal_2567) ) ;
    buf_clk cell_1414 ( .C (CLK), .D (signal_2568), .Q (signal_2569) ) ;
    buf_clk cell_1416 ( .C (CLK), .D (signal_2570), .Q (signal_2571) ) ;
    buf_clk cell_1418 ( .C (CLK), .D (signal_2572), .Q (signal_2573) ) ;
    buf_clk cell_1420 ( .C (CLK), .D (signal_2574), .Q (signal_2575) ) ;
    buf_clk cell_1422 ( .C (CLK), .D (signal_2576), .Q (signal_2577) ) ;
    buf_clk cell_1424 ( .C (CLK), .D (signal_2578), .Q (signal_2579) ) ;
    buf_clk cell_1426 ( .C (CLK), .D (signal_2580), .Q (signal_2581) ) ;
    buf_clk cell_1428 ( .C (CLK), .D (signal_2582), .Q (signal_2583) ) ;
    buf_clk cell_1430 ( .C (CLK), .D (signal_2584), .Q (signal_2585) ) ;
    buf_clk cell_1432 ( .C (CLK), .D (signal_2586), .Q (signal_2587) ) ;
    buf_clk cell_1434 ( .C (CLK), .D (signal_2588), .Q (signal_2589) ) ;
    buf_clk cell_1436 ( .C (CLK), .D (signal_2590), .Q (signal_2591) ) ;
    buf_clk cell_1438 ( .C (CLK), .D (signal_2592), .Q (signal_2593) ) ;
    buf_clk cell_1440 ( .C (CLK), .D (signal_2594), .Q (signal_2595) ) ;
    buf_clk cell_1442 ( .C (CLK), .D (signal_2596), .Q (signal_2597) ) ;
    buf_clk cell_1444 ( .C (CLK), .D (signal_2598), .Q (signal_2599) ) ;
    buf_clk cell_1446 ( .C (CLK), .D (signal_2600), .Q (signal_2601) ) ;
    buf_clk cell_1448 ( .C (CLK), .D (signal_2602), .Q (signal_2603) ) ;
    buf_clk cell_1450 ( .C (CLK), .D (signal_2604), .Q (signal_2605) ) ;
    buf_clk cell_1452 ( .C (CLK), .D (signal_2606), .Q (signal_2607) ) ;
    buf_clk cell_1454 ( .C (CLK), .D (signal_2608), .Q (signal_2609) ) ;
    buf_clk cell_1456 ( .C (CLK), .D (signal_2610), .Q (signal_2611) ) ;
    buf_clk cell_1458 ( .C (CLK), .D (signal_2612), .Q (signal_2613) ) ;
    buf_clk cell_1460 ( .C (CLK), .D (signal_2614), .Q (signal_2615) ) ;
    buf_clk cell_1462 ( .C (CLK), .D (signal_2616), .Q (signal_2617) ) ;
    buf_clk cell_1464 ( .C (CLK), .D (signal_2618), .Q (signal_2619) ) ;
    buf_clk cell_1466 ( .C (CLK), .D (signal_2620), .Q (signal_2621) ) ;
    buf_clk cell_1468 ( .C (CLK), .D (signal_2622), .Q (signal_2623) ) ;
    buf_clk cell_1470 ( .C (CLK), .D (signal_2624), .Q (signal_2625) ) ;
    buf_clk cell_1472 ( .C (CLK), .D (signal_2626), .Q (signal_2627) ) ;
    buf_clk cell_1474 ( .C (CLK), .D (signal_2628), .Q (signal_2629) ) ;
    buf_clk cell_1476 ( .C (CLK), .D (signal_2630), .Q (signal_2631) ) ;
    buf_clk cell_1478 ( .C (CLK), .D (signal_2632), .Q (signal_2633) ) ;
    buf_clk cell_1480 ( .C (CLK), .D (signal_2634), .Q (signal_2635) ) ;
    buf_clk cell_1482 ( .C (CLK), .D (signal_2636), .Q (signal_2637) ) ;
    buf_clk cell_1484 ( .C (CLK), .D (signal_2638), .Q (signal_2639) ) ;
    buf_clk cell_1486 ( .C (CLK), .D (signal_2640), .Q (signal_2641) ) ;
    buf_clk cell_1488 ( .C (CLK), .D (signal_2642), .Q (signal_2643) ) ;
    buf_clk cell_1490 ( .C (CLK), .D (signal_2644), .Q (signal_2645) ) ;
    buf_clk cell_1492 ( .C (CLK), .D (signal_2646), .Q (signal_2647) ) ;
    buf_clk cell_1494 ( .C (CLK), .D (signal_2648), .Q (signal_2649) ) ;
    buf_clk cell_1496 ( .C (CLK), .D (signal_2650), .Q (signal_2651) ) ;
    buf_clk cell_1498 ( .C (CLK), .D (signal_2652), .Q (signal_2653) ) ;
    buf_clk cell_1500 ( .C (CLK), .D (signal_2654), .Q (signal_2655) ) ;
    buf_clk cell_1502 ( .C (CLK), .D (signal_2656), .Q (signal_2657) ) ;
    buf_clk cell_1504 ( .C (CLK), .D (signal_2658), .Q (signal_2659) ) ;
    buf_clk cell_1506 ( .C (CLK), .D (signal_2660), .Q (signal_2661) ) ;
    buf_clk cell_1508 ( .C (CLK), .D (signal_2662), .Q (signal_2663) ) ;
    buf_clk cell_1510 ( .C (CLK), .D (signal_2664), .Q (signal_2665) ) ;
    buf_clk cell_1512 ( .C (CLK), .D (signal_2666), .Q (signal_2667) ) ;
    buf_clk cell_1514 ( .C (CLK), .D (signal_2668), .Q (signal_2669) ) ;
    buf_clk cell_1516 ( .C (CLK), .D (signal_2670), .Q (signal_2671) ) ;
    buf_clk cell_1518 ( .C (CLK), .D (signal_2672), .Q (signal_2673) ) ;
    buf_clk cell_1520 ( .C (CLK), .D (signal_2674), .Q (signal_2675) ) ;
    buf_clk cell_1522 ( .C (CLK), .D (signal_2676), .Q (signal_2677) ) ;
    buf_clk cell_1524 ( .C (CLK), .D (signal_2678), .Q (signal_2679) ) ;
    buf_clk cell_1526 ( .C (CLK), .D (signal_2680), .Q (signal_2681) ) ;
    buf_clk cell_1528 ( .C (CLK), .D (signal_2682), .Q (signal_2683) ) ;
    buf_clk cell_1530 ( .C (CLK), .D (signal_2684), .Q (signal_2685) ) ;
    buf_clk cell_1532 ( .C (CLK), .D (signal_2686), .Q (signal_2687) ) ;
    buf_clk cell_1534 ( .C (CLK), .D (signal_2688), .Q (signal_2689) ) ;
    buf_clk cell_1536 ( .C (CLK), .D (signal_2690), .Q (signal_2691) ) ;
    buf_clk cell_1538 ( .C (CLK), .D (signal_2692), .Q (signal_2693) ) ;
    buf_clk cell_1540 ( .C (CLK), .D (signal_2694), .Q (signal_2695) ) ;
    buf_clk cell_1542 ( .C (CLK), .D (signal_2696), .Q (signal_2697) ) ;
    buf_clk cell_1544 ( .C (CLK), .D (signal_2698), .Q (signal_2699) ) ;
    buf_clk cell_1546 ( .C (CLK), .D (signal_2700), .Q (signal_2701) ) ;
    buf_clk cell_1548 ( .C (CLK), .D (signal_2702), .Q (signal_2703) ) ;
    buf_clk cell_1550 ( .C (CLK), .D (signal_2704), .Q (signal_2705) ) ;
    buf_clk cell_1552 ( .C (CLK), .D (signal_2706), .Q (signal_2707) ) ;
    buf_clk cell_1554 ( .C (CLK), .D (signal_2708), .Q (signal_2709) ) ;
    buf_clk cell_1556 ( .C (CLK), .D (signal_2710), .Q (signal_2711) ) ;
    buf_clk cell_1558 ( .C (CLK), .D (signal_2712), .Q (signal_2713) ) ;
    buf_clk cell_1560 ( .C (CLK), .D (signal_2714), .Q (signal_2715) ) ;
    buf_clk cell_1562 ( .C (CLK), .D (signal_2716), .Q (signal_2717) ) ;
    buf_clk cell_1564 ( .C (CLK), .D (signal_2718), .Q (signal_2719) ) ;
    buf_clk cell_1566 ( .C (CLK), .D (signal_2720), .Q (signal_2721) ) ;
    buf_clk cell_1568 ( .C (CLK), .D (signal_2722), .Q (signal_2723) ) ;
    buf_clk cell_1570 ( .C (CLK), .D (signal_2724), .Q (signal_2725) ) ;
    buf_clk cell_1572 ( .C (CLK), .D (signal_2726), .Q (signal_2727) ) ;
    buf_clk cell_1574 ( .C (CLK), .D (signal_2728), .Q (signal_2729) ) ;
    buf_clk cell_1576 ( .C (CLK), .D (signal_2730), .Q (signal_2731) ) ;
    buf_clk cell_1578 ( .C (CLK), .D (signal_2732), .Q (signal_2733) ) ;
    buf_clk cell_1580 ( .C (CLK), .D (signal_2734), .Q (signal_2735) ) ;
    buf_clk cell_1582 ( .C (CLK), .D (signal_2736), .Q (signal_2737) ) ;
    buf_clk cell_1584 ( .C (CLK), .D (signal_2738), .Q (signal_2739) ) ;
    buf_clk cell_1586 ( .C (CLK), .D (signal_2740), .Q (signal_2741) ) ;
    buf_clk cell_1588 ( .C (CLK), .D (signal_2742), .Q (signal_2743) ) ;
    buf_clk cell_1590 ( .C (CLK), .D (signal_2744), .Q (signal_2745) ) ;
    buf_clk cell_1592 ( .C (CLK), .D (signal_2746), .Q (signal_2747) ) ;
    buf_clk cell_1594 ( .C (CLK), .D (signal_2748), .Q (signal_2749) ) ;
    buf_clk cell_1596 ( .C (CLK), .D (signal_2750), .Q (signal_2751) ) ;
    buf_clk cell_1598 ( .C (CLK), .D (signal_2752), .Q (signal_2753) ) ;
    buf_clk cell_1600 ( .C (CLK), .D (signal_2754), .Q (signal_2755) ) ;
    buf_clk cell_1602 ( .C (CLK), .D (signal_2756), .Q (signal_2757) ) ;
    buf_clk cell_1604 ( .C (CLK), .D (signal_2758), .Q (signal_2759) ) ;
    buf_clk cell_1606 ( .C (CLK), .D (signal_2760), .Q (signal_2761) ) ;
    buf_clk cell_1608 ( .C (CLK), .D (signal_2762), .Q (signal_2763) ) ;
    buf_clk cell_1610 ( .C (CLK), .D (signal_2764), .Q (signal_2765) ) ;
    buf_clk cell_1612 ( .C (CLK), .D (signal_2766), .Q (signal_2767) ) ;
    buf_clk cell_1614 ( .C (CLK), .D (signal_2768), .Q (signal_2769) ) ;
    buf_clk cell_1616 ( .C (CLK), .D (signal_2770), .Q (signal_2771) ) ;
    buf_clk cell_1618 ( .C (CLK), .D (signal_2772), .Q (signal_2773) ) ;
    buf_clk cell_1620 ( .C (CLK), .D (signal_2774), .Q (signal_2775) ) ;
    buf_clk cell_1622 ( .C (CLK), .D (signal_2776), .Q (signal_2777) ) ;
    buf_clk cell_1624 ( .C (CLK), .D (signal_2778), .Q (signal_2779) ) ;
    buf_clk cell_1626 ( .C (CLK), .D (signal_2780), .Q (signal_2781) ) ;
    buf_clk cell_1628 ( .C (CLK), .D (signal_2782), .Q (signal_2783) ) ;
    buf_clk cell_1630 ( .C (CLK), .D (signal_2784), .Q (signal_2785) ) ;
    buf_clk cell_1632 ( .C (CLK), .D (signal_2786), .Q (signal_2787) ) ;
    buf_clk cell_1634 ( .C (CLK), .D (signal_2788), .Q (signal_2789) ) ;
    buf_clk cell_1636 ( .C (CLK), .D (signal_2790), .Q (signal_2791) ) ;
    buf_clk cell_1638 ( .C (CLK), .D (signal_2792), .Q (signal_2793) ) ;
    buf_clk cell_1640 ( .C (CLK), .D (signal_2794), .Q (signal_2795) ) ;
    buf_clk cell_1642 ( .C (CLK), .D (signal_2796), .Q (signal_2797) ) ;
    buf_clk cell_1644 ( .C (CLK), .D (signal_2798), .Q (signal_2799) ) ;
    buf_clk cell_1646 ( .C (CLK), .D (signal_2800), .Q (signal_2801) ) ;
    buf_clk cell_1648 ( .C (CLK), .D (signal_2802), .Q (signal_2803) ) ;
    buf_clk cell_1650 ( .C (CLK), .D (signal_2804), .Q (signal_2805) ) ;
    buf_clk cell_1652 ( .C (CLK), .D (signal_2806), .Q (signal_2807) ) ;
    buf_clk cell_1654 ( .C (CLK), .D (signal_2808), .Q (signal_2809) ) ;
    buf_clk cell_1656 ( .C (CLK), .D (signal_2810), .Q (signal_2811) ) ;
    buf_clk cell_1658 ( .C (CLK), .D (signal_2812), .Q (signal_2813) ) ;
    buf_clk cell_1660 ( .C (CLK), .D (signal_2814), .Q (signal_2815) ) ;
    buf_clk cell_1662 ( .C (CLK), .D (signal_2816), .Q (signal_2817) ) ;
    buf_clk cell_1664 ( .C (CLK), .D (signal_2818), .Q (signal_2819) ) ;
    buf_clk cell_1666 ( .C (CLK), .D (signal_2820), .Q (signal_2821) ) ;
    buf_clk cell_1668 ( .C (CLK), .D (signal_2822), .Q (signal_2823) ) ;
    buf_clk cell_1670 ( .C (CLK), .D (signal_2824), .Q (signal_2825) ) ;
    buf_clk cell_1672 ( .C (CLK), .D (signal_2826), .Q (signal_2827) ) ;
    buf_clk cell_1674 ( .C (CLK), .D (signal_2828), .Q (signal_2829) ) ;
    buf_clk cell_1676 ( .C (CLK), .D (signal_2830), .Q (signal_2831) ) ;
    buf_clk cell_1678 ( .C (CLK), .D (signal_2832), .Q (signal_2833) ) ;
    buf_clk cell_1680 ( .C (CLK), .D (signal_2834), .Q (signal_2835) ) ;
    buf_clk cell_1682 ( .C (CLK), .D (signal_2836), .Q (signal_2837) ) ;
    buf_clk cell_1684 ( .C (CLK), .D (signal_2838), .Q (signal_2839) ) ;
    buf_clk cell_1686 ( .C (CLK), .D (signal_2840), .Q (signal_2841) ) ;
    buf_clk cell_1688 ( .C (CLK), .D (signal_2842), .Q (signal_2843) ) ;
    buf_clk cell_1690 ( .C (CLK), .D (signal_2844), .Q (signal_2845) ) ;
    buf_clk cell_1692 ( .C (CLK), .D (signal_2846), .Q (signal_2847) ) ;
    buf_clk cell_1694 ( .C (CLK), .D (signal_2848), .Q (signal_2849) ) ;
    buf_clk cell_1696 ( .C (CLK), .D (signal_2850), .Q (signal_2851) ) ;
    buf_clk cell_1698 ( .C (CLK), .D (signal_2852), .Q (signal_2853) ) ;
    buf_clk cell_1700 ( .C (CLK), .D (signal_2854), .Q (signal_2855) ) ;
    buf_clk cell_1702 ( .C (CLK), .D (signal_2856), .Q (signal_2857) ) ;
    buf_clk cell_1704 ( .C (CLK), .D (signal_2858), .Q (signal_2859) ) ;

    /* register cells */
    DFF_X1 cell_979 ( .CK (CLK), .D (signal_2839), .Q (signal_808), .QN () ) ;
    DFF_X1 cell_981 ( .CK (CLK), .D (signal_2841), .Q (signal_307), .QN () ) ;
    DFF_X1 cell_983 ( .CK (CLK), .D (signal_2843), .Q (signal_304), .QN () ) ;
    DFF_X1 cell_985 ( .CK (CLK), .D (signal_2845), .Q (signal_288), .QN () ) ;
    DFF_X1 cell_987 ( .CK (CLK), .D (signal_2847), .Q (signal_879), .QN () ) ;
    DFF_X1 cell_989 ( .CK (CLK), .D (signal_2849), .Q (signal_878), .QN () ) ;
    DFF_X1 cell_991 ( .CK (CLK), .D (signal_2851), .Q (signal_877), .QN () ) ;
    DFF_X1 cell_993 ( .CK (CLK), .D (signal_2853), .Q (signal_876), .QN () ) ;
    DFF_X1 cell_995 ( .CK (CLK), .D (signal_2855), .Q (signal_875), .QN () ) ;
    DFF_X1 cell_997 ( .CK (CLK), .D (signal_2857), .Q (signal_874), .QN () ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_999 ( .clk (CLK), .D ({signal_1917, signal_1199}), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1001 ( .clk (CLK), .D ({signal_2001, signal_1198}), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1003 ( .clk (CLK), .D ({signal_1919, signal_1197}), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1005 ( .clk (CLK), .D ({signal_1965, signal_1196}), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1007 ( .clk (CLK), .D ({signal_1921, signal_1195}), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1009 ( .clk (CLK), .D ({signal_2003, signal_1194}), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1011 ( .clk (CLK), .D ({signal_1923, signal_1193}), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1013 ( .clk (CLK), .D ({signal_1967, signal_1192}), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1015 ( .clk (CLK), .D ({signal_1925, signal_1191}), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1017 ( .clk (CLK), .D ({signal_2005, signal_1190}), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1019 ( .clk (CLK), .D ({signal_1927, signal_1189}), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1021 ( .clk (CLK), .D ({signal_1969, signal_1188}), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1023 ( .clk (CLK), .D ({signal_1929, signal_1187}), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1025 ( .clk (CLK), .D ({signal_2007, signal_1186}), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1027 ( .clk (CLK), .D ({signal_1931, signal_1185}), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1029 ( .clk (CLK), .D ({signal_1971, signal_1184}), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1031 ( .clk (CLK), .D ({signal_2061, signal_1183}), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1033 ( .clk (CLK), .D ({signal_2085, signal_1182}), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1035 ( .clk (CLK), .D ({signal_2087, signal_1181}), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1037 ( .clk (CLK), .D ({signal_2009, signal_1180}), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1039 ( .clk (CLK), .D ({signal_2063, signal_1179}), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1041 ( .clk (CLK), .D ({signal_2089, signal_1178}), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1043 ( .clk (CLK), .D ({signal_2091, signal_1177}), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1045 ( .clk (CLK), .D ({signal_2011, signal_1176}), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1047 ( .clk (CLK), .D ({signal_2065, signal_1175}), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1049 ( .clk (CLK), .D ({signal_2093, signal_1174}), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1051 ( .clk (CLK), .D ({signal_2095, signal_1173}), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1053 ( .clk (CLK), .D ({signal_2013, signal_1172}), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1055 ( .clk (CLK), .D ({signal_2067, signal_1171}), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1057 ( .clk (CLK), .D ({signal_2097, signal_1170}), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1059 ( .clk (CLK), .D ({signal_2099, signal_1169}), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1061 ( .clk (CLK), .D ({signal_2015, signal_1168}), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1063 ( .clk (CLK), .D ({signal_2101, signal_1167}), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1065 ( .clk (CLK), .D ({signal_2141, signal_1166}), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1067 ( .clk (CLK), .D ({signal_2103, signal_1165}), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1069 ( .clk (CLK), .D ({signal_2153, signal_1164}), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1071 ( .clk (CLK), .D ({signal_2105, signal_1163}), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1073 ( .clk (CLK), .D ({signal_2143, signal_1162}), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1075 ( .clk (CLK), .D ({signal_2107, signal_1161}), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1077 ( .clk (CLK), .D ({signal_2155, signal_1160}), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1079 ( .clk (CLK), .D ({signal_2109, signal_1159}), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1081 ( .clk (CLK), .D ({signal_2145, signal_1158}), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1083 ( .clk (CLK), .D ({signal_2111, signal_1157}), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1085 ( .clk (CLK), .D ({signal_2157, signal_1156}), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1087 ( .clk (CLK), .D ({signal_2113, signal_1155}), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1089 ( .clk (CLK), .D ({signal_2147, signal_1154}), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1091 ( .clk (CLK), .D ({signal_2115, signal_1153}), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1093 ( .clk (CLK), .D ({signal_2159, signal_1152}), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1095 ( .clk (CLK), .D ({signal_2205, signal_1151}), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1097 ( .clk (CLK), .D ({signal_2213, signal_1150}), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1099 ( .clk (CLK), .D ({signal_2161, signal_1149}), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1101 ( .clk (CLK), .D ({signal_2163, signal_1148}), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1103 ( .clk (CLK), .D ({signal_2207, signal_1147}), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1105 ( .clk (CLK), .D ({signal_2215, signal_1146}), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1107 ( .clk (CLK), .D ({signal_2165, signal_1145}), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1109 ( .clk (CLK), .D ({signal_2167, signal_1144}), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1111 ( .clk (CLK), .D ({signal_2209, signal_1143}), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1113 ( .clk (CLK), .D ({signal_2217, signal_1142}), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1115 ( .clk (CLK), .D ({signal_2169, signal_1141}), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1117 ( .clk (CLK), .D ({signal_2171, signal_1140}), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1119 ( .clk (CLK), .D ({signal_2211, signal_1139}), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1121 ( .clk (CLK), .D ({signal_2219, signal_1138}), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1123 ( .clk (CLK), .D ({signal_2173, signal_1137}), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(1)) cell_1125 ( .clk (CLK), .D ({signal_2175, signal_1136}), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    DFF_X1 cell_1127 ( .CK (CLK), .D (signal_2859), .Q (OUT_done), .QN () ) ;
endmodule
