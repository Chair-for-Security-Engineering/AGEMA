/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 16 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 17 register stage(s) in total */

module sbox_HPC2_BDDcudd_Pipeline_d3 (X_s0, clk, X_s1, X_s2, X_s3, Fresh, Y_s0, Y_s1, Y_s2, Y_s3);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [7:0] X_s3 ;
    input [2465:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output [7:0] Y_s3 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_557 ;
    wire signal_558 ;
    wire signal_559 ;
    wire signal_563 ;
    wire signal_564 ;
    wire signal_565 ;
    wire signal_566 ;
    wire signal_567 ;
    wire signal_568 ;
    wire signal_572 ;
    wire signal_573 ;
    wire signal_574 ;
    wire signal_575 ;
    wire signal_576 ;
    wire signal_577 ;
    wire signal_578 ;
    wire signal_579 ;
    wire signal_580 ;
    wire signal_581 ;
    wire signal_582 ;
    wire signal_583 ;
    wire signal_584 ;
    wire signal_585 ;
    wire signal_586 ;
    wire signal_587 ;
    wire signal_588 ;
    wire signal_589 ;
    wire signal_590 ;
    wire signal_591 ;
    wire signal_592 ;
    wire signal_593 ;
    wire signal_594 ;
    wire signal_595 ;
    wire signal_596 ;
    wire signal_597 ;
    wire signal_598 ;
    wire signal_599 ;
    wire signal_600 ;
    wire signal_601 ;
    wire signal_602 ;
    wire signal_603 ;
    wire signal_604 ;
    wire signal_605 ;
    wire signal_606 ;
    wire signal_607 ;
    wire signal_608 ;
    wire signal_609 ;
    wire signal_610 ;
    wire signal_611 ;
    wire signal_612 ;
    wire signal_613 ;
    wire signal_614 ;
    wire signal_615 ;
    wire signal_616 ;
    wire signal_617 ;
    wire signal_618 ;
    wire signal_619 ;
    wire signal_620 ;
    wire signal_621 ;
    wire signal_622 ;
    wire signal_623 ;
    wire signal_624 ;
    wire signal_625 ;
    wire signal_626 ;
    wire signal_627 ;
    wire signal_628 ;
    wire signal_629 ;
    wire signal_630 ;
    wire signal_631 ;
    wire signal_632 ;
    wire signal_633 ;
    wire signal_634 ;
    wire signal_635 ;
    wire signal_636 ;
    wire signal_637 ;
    wire signal_638 ;
    wire signal_639 ;
    wire signal_640 ;
    wire signal_641 ;
    wire signal_642 ;
    wire signal_643 ;
    wire signal_644 ;
    wire signal_645 ;
    wire signal_646 ;
    wire signal_647 ;
    wire signal_648 ;
    wire signal_649 ;
    wire signal_650 ;
    wire signal_651 ;
    wire signal_652 ;
    wire signal_653 ;
    wire signal_654 ;
    wire signal_655 ;
    wire signal_656 ;
    wire signal_657 ;
    wire signal_658 ;
    wire signal_659 ;
    wire signal_660 ;
    wire signal_661 ;
    wire signal_662 ;
    wire signal_663 ;
    wire signal_664 ;
    wire signal_665 ;
    wire signal_666 ;
    wire signal_667 ;
    wire signal_668 ;
    wire signal_669 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;
    wire signal_4762 ;
    wire signal_4763 ;
    wire signal_4764 ;
    wire signal_4765 ;
    wire signal_4766 ;
    wire signal_4767 ;
    wire signal_4768 ;
    wire signal_4769 ;
    wire signal_4770 ;
    wire signal_4771 ;
    wire signal_4772 ;
    wire signal_4773 ;
    wire signal_4774 ;
    wire signal_4775 ;
    wire signal_4776 ;
    wire signal_4777 ;
    wire signal_4778 ;
    wire signal_4779 ;
    wire signal_4780 ;
    wire signal_4781 ;
    wire signal_4782 ;
    wire signal_4783 ;
    wire signal_4784 ;
    wire signal_4785 ;
    wire signal_4786 ;
    wire signal_4787 ;
    wire signal_4788 ;
    wire signal_4789 ;
    wire signal_4790 ;
    wire signal_4791 ;
    wire signal_4792 ;
    wire signal_4793 ;
    wire signal_4794 ;
    wire signal_4795 ;
    wire signal_4796 ;
    wire signal_4797 ;
    wire signal_4798 ;
    wire signal_4799 ;
    wire signal_4800 ;
    wire signal_4801 ;
    wire signal_4802 ;
    wire signal_4803 ;
    wire signal_4804 ;
    wire signal_4805 ;
    wire signal_4806 ;
    wire signal_4807 ;
    wire signal_4808 ;
    wire signal_4809 ;
    wire signal_4810 ;
    wire signal_4811 ;
    wire signal_4812 ;

    /* cells in depth 0 */

    /* cells in depth 1 */
    buf_clk cell_547 ( .C (clk), .D (X_s0[5]), .Q (signal_4301) ) ;
    buf_clk cell_549 ( .C (clk), .D (X_s1[5]), .Q (signal_4303) ) ;
    buf_clk cell_551 ( .C (clk), .D (X_s2[5]), .Q (signal_4305) ) ;
    buf_clk cell_553 ( .C (clk), .D (X_s3[5]), .Q (signal_4307) ) ;
    buf_clk cell_555 ( .C (clk), .D (X_s0[6]), .Q (signal_4309) ) ;
    buf_clk cell_557 ( .C (clk), .D (X_s1[6]), .Q (signal_4311) ) ;
    buf_clk cell_559 ( .C (clk), .D (X_s2[6]), .Q (signal_4313) ) ;
    buf_clk cell_561 ( .C (clk), .D (X_s3[6]), .Q (signal_4315) ) ;
    buf_clk cell_603 ( .C (clk), .D (X_s0[3]), .Q (signal_4357) ) ;
    buf_clk cell_607 ( .C (clk), .D (X_s1[3]), .Q (signal_4361) ) ;
    buf_clk cell_611 ( .C (clk), .D (X_s2[3]), .Q (signal_4365) ) ;
    buf_clk cell_615 ( .C (clk), .D (X_s3[3]), .Q (signal_4369) ) ;
    buf_clk cell_835 ( .C (clk), .D (X_s0[1]), .Q (signal_4589) ) ;
    buf_clk cell_843 ( .C (clk), .D (X_s1[1]), .Q (signal_4597) ) ;
    buf_clk cell_851 ( .C (clk), .D (X_s2[1]), .Q (signal_4605) ) ;
    buf_clk cell_859 ( .C (clk), .D (X_s3[1]), .Q (signal_4613) ) ;
    buf_clk cell_915 ( .C (clk), .D (X_s0[2]), .Q (signal_4669) ) ;
    buf_clk cell_925 ( .C (clk), .D (X_s1[2]), .Q (signal_4679) ) ;
    buf_clk cell_935 ( .C (clk), .D (X_s2[2]), .Q (signal_4689) ) ;
    buf_clk cell_945 ( .C (clk), .D (X_s3[2]), .Q (signal_4699) ) ;
    buf_clk cell_955 ( .C (clk), .D (X_s0[4]), .Q (signal_4709) ) ;
    buf_clk cell_967 ( .C (clk), .D (X_s1[4]), .Q (signal_4721) ) ;
    buf_clk cell_979 ( .C (clk), .D (X_s2[4]), .Q (signal_4733) ) ;
    buf_clk cell_991 ( .C (clk), .D (X_s3[4]), .Q (signal_4745) ) ;
    buf_clk cell_1003 ( .C (clk), .D (X_s0[7]), .Q (signal_4757) ) ;
    buf_clk cell_1017 ( .C (clk), .D (X_s1[7]), .Q (signal_4771) ) ;
    buf_clk cell_1031 ( .C (clk), .D (X_s2[7]), .Q (signal_4785) ) ;
    buf_clk cell_1045 ( .C (clk), .D (X_s3[7]), .Q (signal_4799) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_136 ( .s ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_559, signal_558, signal_557, signal_151}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_137 ( .s ({X_s3[6], X_s2[6], X_s1[6], X_s0[6]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_565, signal_564, signal_563, signal_152}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_138 ( .s ({X_s3[5], X_s2[5], X_s1[5], X_s0[5]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_568, signal_567, signal_566, signal_153}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_139 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_574, signal_573, signal_572, signal_154}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_140 ( .s ({X_s3[0], X_s2[0], X_s1[0], X_s0[0]}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_577, signal_576, signal_575, signal_155}) ) ;
    buf_clk cell_548 ( .C (clk), .D (signal_4301), .Q (signal_4302) ) ;
    buf_clk cell_550 ( .C (clk), .D (signal_4303), .Q (signal_4304) ) ;
    buf_clk cell_552 ( .C (clk), .D (signal_4305), .Q (signal_4306) ) ;
    buf_clk cell_554 ( .C (clk), .D (signal_4307), .Q (signal_4308) ) ;
    buf_clk cell_556 ( .C (clk), .D (signal_4309), .Q (signal_4310) ) ;
    buf_clk cell_558 ( .C (clk), .D (signal_4311), .Q (signal_4312) ) ;
    buf_clk cell_560 ( .C (clk), .D (signal_4313), .Q (signal_4314) ) ;
    buf_clk cell_562 ( .C (clk), .D (signal_4315), .Q (signal_4316) ) ;
    buf_clk cell_604 ( .C (clk), .D (signal_4357), .Q (signal_4358) ) ;
    buf_clk cell_608 ( .C (clk), .D (signal_4361), .Q (signal_4362) ) ;
    buf_clk cell_612 ( .C (clk), .D (signal_4365), .Q (signal_4366) ) ;
    buf_clk cell_616 ( .C (clk), .D (signal_4369), .Q (signal_4370) ) ;
    buf_clk cell_836 ( .C (clk), .D (signal_4589), .Q (signal_4590) ) ;
    buf_clk cell_844 ( .C (clk), .D (signal_4597), .Q (signal_4598) ) ;
    buf_clk cell_852 ( .C (clk), .D (signal_4605), .Q (signal_4606) ) ;
    buf_clk cell_860 ( .C (clk), .D (signal_4613), .Q (signal_4614) ) ;
    buf_clk cell_916 ( .C (clk), .D (signal_4669), .Q (signal_4670) ) ;
    buf_clk cell_926 ( .C (clk), .D (signal_4679), .Q (signal_4680) ) ;
    buf_clk cell_936 ( .C (clk), .D (signal_4689), .Q (signal_4690) ) ;
    buf_clk cell_946 ( .C (clk), .D (signal_4699), .Q (signal_4700) ) ;
    buf_clk cell_956 ( .C (clk), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_968 ( .C (clk), .D (signal_4721), .Q (signal_4722) ) ;
    buf_clk cell_980 ( .C (clk), .D (signal_4733), .Q (signal_4734) ) ;
    buf_clk cell_992 ( .C (clk), .D (signal_4745), .Q (signal_4746) ) ;
    buf_clk cell_1004 ( .C (clk), .D (signal_4757), .Q (signal_4758) ) ;
    buf_clk cell_1018 ( .C (clk), .D (signal_4771), .Q (signal_4772) ) ;
    buf_clk cell_1032 ( .C (clk), .D (signal_4785), .Q (signal_4786) ) ;
    buf_clk cell_1046 ( .C (clk), .D (signal_4799), .Q (signal_4800) ) ;

    /* cells in depth 3 */
    buf_clk cell_563 ( .C (clk), .D (signal_4310), .Q (signal_4317) ) ;
    buf_clk cell_565 ( .C (clk), .D (signal_4312), .Q (signal_4319) ) ;
    buf_clk cell_567 ( .C (clk), .D (signal_4314), .Q (signal_4321) ) ;
    buf_clk cell_569 ( .C (clk), .D (signal_4316), .Q (signal_4323) ) ;
    buf_clk cell_571 ( .C (clk), .D (signal_153), .Q (signal_4325) ) ;
    buf_clk cell_573 ( .C (clk), .D (signal_566), .Q (signal_4327) ) ;
    buf_clk cell_575 ( .C (clk), .D (signal_567), .Q (signal_4329) ) ;
    buf_clk cell_577 ( .C (clk), .D (signal_568), .Q (signal_4331) ) ;
    buf_clk cell_579 ( .C (clk), .D (signal_154), .Q (signal_4333) ) ;
    buf_clk cell_581 ( .C (clk), .D (signal_572), .Q (signal_4335) ) ;
    buf_clk cell_583 ( .C (clk), .D (signal_573), .Q (signal_4337) ) ;
    buf_clk cell_585 ( .C (clk), .D (signal_574), .Q (signal_4339) ) ;
    buf_clk cell_587 ( .C (clk), .D (signal_151), .Q (signal_4341) ) ;
    buf_clk cell_589 ( .C (clk), .D (signal_557), .Q (signal_4343) ) ;
    buf_clk cell_591 ( .C (clk), .D (signal_558), .Q (signal_4345) ) ;
    buf_clk cell_593 ( .C (clk), .D (signal_559), .Q (signal_4347) ) ;
    buf_clk cell_595 ( .C (clk), .D (signal_155), .Q (signal_4349) ) ;
    buf_clk cell_597 ( .C (clk), .D (signal_575), .Q (signal_4351) ) ;
    buf_clk cell_599 ( .C (clk), .D (signal_576), .Q (signal_4353) ) ;
    buf_clk cell_601 ( .C (clk), .D (signal_577), .Q (signal_4355) ) ;
    buf_clk cell_605 ( .C (clk), .D (signal_4358), .Q (signal_4359) ) ;
    buf_clk cell_609 ( .C (clk), .D (signal_4362), .Q (signal_4363) ) ;
    buf_clk cell_613 ( .C (clk), .D (signal_4366), .Q (signal_4367) ) ;
    buf_clk cell_617 ( .C (clk), .D (signal_4370), .Q (signal_4371) ) ;
    buf_clk cell_619 ( .C (clk), .D (signal_152), .Q (signal_4373) ) ;
    buf_clk cell_621 ( .C (clk), .D (signal_563), .Q (signal_4375) ) ;
    buf_clk cell_623 ( .C (clk), .D (signal_564), .Q (signal_4377) ) ;
    buf_clk cell_625 ( .C (clk), .D (signal_565), .Q (signal_4379) ) ;
    buf_clk cell_837 ( .C (clk), .D (signal_4590), .Q (signal_4591) ) ;
    buf_clk cell_845 ( .C (clk), .D (signal_4598), .Q (signal_4599) ) ;
    buf_clk cell_853 ( .C (clk), .D (signal_4606), .Q (signal_4607) ) ;
    buf_clk cell_861 ( .C (clk), .D (signal_4614), .Q (signal_4615) ) ;
    buf_clk cell_917 ( .C (clk), .D (signal_4670), .Q (signal_4671) ) ;
    buf_clk cell_927 ( .C (clk), .D (signal_4680), .Q (signal_4681) ) ;
    buf_clk cell_937 ( .C (clk), .D (signal_4690), .Q (signal_4691) ) ;
    buf_clk cell_947 ( .C (clk), .D (signal_4700), .Q (signal_4701) ) ;
    buf_clk cell_957 ( .C (clk), .D (signal_4710), .Q (signal_4711) ) ;
    buf_clk cell_969 ( .C (clk), .D (signal_4722), .Q (signal_4723) ) ;
    buf_clk cell_981 ( .C (clk), .D (signal_4734), .Q (signal_4735) ) ;
    buf_clk cell_993 ( .C (clk), .D (signal_4746), .Q (signal_4747) ) ;
    buf_clk cell_1005 ( .C (clk), .D (signal_4758), .Q (signal_4759) ) ;
    buf_clk cell_1019 ( .C (clk), .D (signal_4772), .Q (signal_4773) ) ;
    buf_clk cell_1033 ( .C (clk), .D (signal_4786), .Q (signal_4787) ) ;
    buf_clk cell_1047 ( .C (clk), .D (signal_4800), .Q (signal_4801) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_141 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({signal_577, signal_576, signal_575, signal_155}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_580, signal_579, signal_578, signal_156}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_142 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_577, signal_576, signal_575, signal_155}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_583, signal_582, signal_581, signal_157}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_143 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({signal_574, signal_573, signal_572, signal_154}), .a ({signal_577, signal_576, signal_575, signal_155}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_586, signal_585, signal_584, signal_158}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_144 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_568, signal_567, signal_566, signal_153}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_589, signal_588, signal_587, signal_159}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_145 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_577, signal_576, signal_575, signal_155}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_592, signal_591, signal_590, signal_160}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_146 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_568, signal_567, signal_566, signal_153}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_595, signal_594, signal_593, signal_161}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_147 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({signal_577, signal_576, signal_575, signal_155}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_598, signal_597, signal_596, signal_162}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_148 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_559, signal_558, signal_557, signal_151}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_601, signal_600, signal_599, signal_163}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_149 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_568, signal_567, signal_566, signal_153}), .a ({signal_577, signal_576, signal_575, signal_155}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_604, signal_603, signal_602, signal_164}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_150 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({signal_574, signal_573, signal_572, signal_154}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_607, signal_606, signal_605, signal_165}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_151 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_559, signal_558, signal_557, signal_151}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_610, signal_609, signal_608, signal_166}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_152 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_574, signal_573, signal_572, signal_154}), .a ({signal_559, signal_558, signal_557, signal_151}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_613, signal_612, signal_611, signal_167}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_153 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({signal_616, signal_615, signal_614, signal_168}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_154 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({signal_619, signal_618, signal_617, signal_169}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_155 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({signal_622, signal_621, signal_620, signal_170}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_156 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_559, signal_558, signal_557, signal_151}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({signal_625, signal_624, signal_623, signal_171}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_157 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({signal_628, signal_627, signal_626, signal_172}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_158 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_568, signal_567, signal_566, signal_153}), .a ({signal_559, signal_558, signal_557, signal_151}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({signal_631, signal_630, signal_629, signal_173}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_159 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({signal_574, signal_573, signal_572, signal_154}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({signal_634, signal_633, signal_632, signal_174}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_160 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_577, signal_576, signal_575, signal_155}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({signal_637, signal_636, signal_635, signal_175}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_161 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_568, signal_567, signal_566, signal_153}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({signal_640, signal_639, signal_638, signal_176}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_162 ( .s ({signal_4308, signal_4306, signal_4304, signal_4302}), .b ({signal_577, signal_576, signal_575, signal_155}), .a ({signal_574, signal_573, signal_572, signal_154}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({signal_643, signal_642, signal_641, signal_177}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_163 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_559, signal_558, signal_557, signal_151}), .a ({signal_568, signal_567, signal_566, signal_153}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({signal_646, signal_645, signal_644, signal_178}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_164 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_574, signal_573, signal_572, signal_154}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({signal_649, signal_648, signal_647, signal_179}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_165 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_577, signal_576, signal_575, signal_155}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({signal_652, signal_651, signal_650, signal_180}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_166 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_577, signal_576, signal_575, signal_155}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({signal_655, signal_654, signal_653, signal_181}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_167 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_577, signal_576, signal_575, signal_155}), .a ({signal_559, signal_558, signal_557, signal_151}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({signal_658, signal_657, signal_656, signal_182}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_168 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({signal_568, signal_567, signal_566, signal_153}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({signal_661, signal_660, signal_659, signal_183}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_169 ( .s ({signal_4316, signal_4314, signal_4312, signal_4310}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_559, signal_558, signal_557, signal_151}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({signal_664, signal_663, signal_662, signal_184}) ) ;
    buf_clk cell_564 ( .C (clk), .D (signal_4317), .Q (signal_4318) ) ;
    buf_clk cell_566 ( .C (clk), .D (signal_4319), .Q (signal_4320) ) ;
    buf_clk cell_568 ( .C (clk), .D (signal_4321), .Q (signal_4322) ) ;
    buf_clk cell_570 ( .C (clk), .D (signal_4323), .Q (signal_4324) ) ;
    buf_clk cell_572 ( .C (clk), .D (signal_4325), .Q (signal_4326) ) ;
    buf_clk cell_574 ( .C (clk), .D (signal_4327), .Q (signal_4328) ) ;
    buf_clk cell_576 ( .C (clk), .D (signal_4329), .Q (signal_4330) ) ;
    buf_clk cell_578 ( .C (clk), .D (signal_4331), .Q (signal_4332) ) ;
    buf_clk cell_580 ( .C (clk), .D (signal_4333), .Q (signal_4334) ) ;
    buf_clk cell_582 ( .C (clk), .D (signal_4335), .Q (signal_4336) ) ;
    buf_clk cell_584 ( .C (clk), .D (signal_4337), .Q (signal_4338) ) ;
    buf_clk cell_586 ( .C (clk), .D (signal_4339), .Q (signal_4340) ) ;
    buf_clk cell_588 ( .C (clk), .D (signal_4341), .Q (signal_4342) ) ;
    buf_clk cell_590 ( .C (clk), .D (signal_4343), .Q (signal_4344) ) ;
    buf_clk cell_592 ( .C (clk), .D (signal_4345), .Q (signal_4346) ) ;
    buf_clk cell_594 ( .C (clk), .D (signal_4347), .Q (signal_4348) ) ;
    buf_clk cell_596 ( .C (clk), .D (signal_4349), .Q (signal_4350) ) ;
    buf_clk cell_598 ( .C (clk), .D (signal_4351), .Q (signal_4352) ) ;
    buf_clk cell_600 ( .C (clk), .D (signal_4353), .Q (signal_4354) ) ;
    buf_clk cell_602 ( .C (clk), .D (signal_4355), .Q (signal_4356) ) ;
    buf_clk cell_606 ( .C (clk), .D (signal_4359), .Q (signal_4360) ) ;
    buf_clk cell_610 ( .C (clk), .D (signal_4363), .Q (signal_4364) ) ;
    buf_clk cell_614 ( .C (clk), .D (signal_4367), .Q (signal_4368) ) ;
    buf_clk cell_618 ( .C (clk), .D (signal_4371), .Q (signal_4372) ) ;
    buf_clk cell_620 ( .C (clk), .D (signal_4373), .Q (signal_4374) ) ;
    buf_clk cell_622 ( .C (clk), .D (signal_4375), .Q (signal_4376) ) ;
    buf_clk cell_624 ( .C (clk), .D (signal_4377), .Q (signal_4378) ) ;
    buf_clk cell_626 ( .C (clk), .D (signal_4379), .Q (signal_4380) ) ;
    buf_clk cell_838 ( .C (clk), .D (signal_4591), .Q (signal_4592) ) ;
    buf_clk cell_846 ( .C (clk), .D (signal_4599), .Q (signal_4600) ) ;
    buf_clk cell_854 ( .C (clk), .D (signal_4607), .Q (signal_4608) ) ;
    buf_clk cell_862 ( .C (clk), .D (signal_4615), .Q (signal_4616) ) ;
    buf_clk cell_918 ( .C (clk), .D (signal_4671), .Q (signal_4672) ) ;
    buf_clk cell_928 ( .C (clk), .D (signal_4681), .Q (signal_4682) ) ;
    buf_clk cell_938 ( .C (clk), .D (signal_4691), .Q (signal_4692) ) ;
    buf_clk cell_948 ( .C (clk), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_958 ( .C (clk), .D (signal_4711), .Q (signal_4712) ) ;
    buf_clk cell_970 ( .C (clk), .D (signal_4723), .Q (signal_4724) ) ;
    buf_clk cell_982 ( .C (clk), .D (signal_4735), .Q (signal_4736) ) ;
    buf_clk cell_994 ( .C (clk), .D (signal_4747), .Q (signal_4748) ) ;
    buf_clk cell_1006 ( .C (clk), .D (signal_4759), .Q (signal_4760) ) ;
    buf_clk cell_1020 ( .C (clk), .D (signal_4773), .Q (signal_4774) ) ;
    buf_clk cell_1034 ( .C (clk), .D (signal_4787), .Q (signal_4788) ) ;
    buf_clk cell_1048 ( .C (clk), .D (signal_4801), .Q (signal_4802) ) ;

    /* cells in depth 5 */
    buf_clk cell_627 ( .C (clk), .D (signal_4360), .Q (signal_4381) ) ;
    buf_clk cell_629 ( .C (clk), .D (signal_4364), .Q (signal_4383) ) ;
    buf_clk cell_631 ( .C (clk), .D (signal_4368), .Q (signal_4385) ) ;
    buf_clk cell_633 ( .C (clk), .D (signal_4372), .Q (signal_4387) ) ;
    buf_clk cell_635 ( .C (clk), .D (signal_4342), .Q (signal_4389) ) ;
    buf_clk cell_637 ( .C (clk), .D (signal_4344), .Q (signal_4391) ) ;
    buf_clk cell_639 ( .C (clk), .D (signal_4346), .Q (signal_4393) ) ;
    buf_clk cell_641 ( .C (clk), .D (signal_4348), .Q (signal_4395) ) ;
    buf_clk cell_643 ( .C (clk), .D (signal_4374), .Q (signal_4397) ) ;
    buf_clk cell_645 ( .C (clk), .D (signal_4376), .Q (signal_4399) ) ;
    buf_clk cell_647 ( .C (clk), .D (signal_4378), .Q (signal_4401) ) ;
    buf_clk cell_649 ( .C (clk), .D (signal_4380), .Q (signal_4403) ) ;
    buf_clk cell_651 ( .C (clk), .D (signal_182), .Q (signal_4405) ) ;
    buf_clk cell_653 ( .C (clk), .D (signal_656), .Q (signal_4407) ) ;
    buf_clk cell_655 ( .C (clk), .D (signal_657), .Q (signal_4409) ) ;
    buf_clk cell_657 ( .C (clk), .D (signal_658), .Q (signal_4411) ) ;
    buf_clk cell_659 ( .C (clk), .D (signal_175), .Q (signal_4413) ) ;
    buf_clk cell_661 ( .C (clk), .D (signal_635), .Q (signal_4415) ) ;
    buf_clk cell_663 ( .C (clk), .D (signal_636), .Q (signal_4417) ) ;
    buf_clk cell_665 ( .C (clk), .D (signal_637), .Q (signal_4419) ) ;
    buf_clk cell_667 ( .C (clk), .D (signal_177), .Q (signal_4421) ) ;
    buf_clk cell_669 ( .C (clk), .D (signal_641), .Q (signal_4423) ) ;
    buf_clk cell_671 ( .C (clk), .D (signal_642), .Q (signal_4425) ) ;
    buf_clk cell_673 ( .C (clk), .D (signal_643), .Q (signal_4427) ) ;
    buf_clk cell_675 ( .C (clk), .D (signal_169), .Q (signal_4429) ) ;
    buf_clk cell_677 ( .C (clk), .D (signal_617), .Q (signal_4431) ) ;
    buf_clk cell_679 ( .C (clk), .D (signal_618), .Q (signal_4433) ) ;
    buf_clk cell_681 ( .C (clk), .D (signal_619), .Q (signal_4435) ) ;
    buf_clk cell_683 ( .C (clk), .D (signal_178), .Q (signal_4437) ) ;
    buf_clk cell_685 ( .C (clk), .D (signal_644), .Q (signal_4439) ) ;
    buf_clk cell_687 ( .C (clk), .D (signal_645), .Q (signal_4441) ) ;
    buf_clk cell_689 ( .C (clk), .D (signal_646), .Q (signal_4443) ) ;
    buf_clk cell_691 ( .C (clk), .D (signal_167), .Q (signal_4445) ) ;
    buf_clk cell_693 ( .C (clk), .D (signal_611), .Q (signal_4447) ) ;
    buf_clk cell_695 ( .C (clk), .D (signal_612), .Q (signal_4449) ) ;
    buf_clk cell_697 ( .C (clk), .D (signal_613), .Q (signal_4451) ) ;
    buf_clk cell_699 ( .C (clk), .D (signal_171), .Q (signal_4453) ) ;
    buf_clk cell_701 ( .C (clk), .D (signal_623), .Q (signal_4455) ) ;
    buf_clk cell_703 ( .C (clk), .D (signal_624), .Q (signal_4457) ) ;
    buf_clk cell_705 ( .C (clk), .D (signal_625), .Q (signal_4459) ) ;
    buf_clk cell_707 ( .C (clk), .D (signal_183), .Q (signal_4461) ) ;
    buf_clk cell_709 ( .C (clk), .D (signal_659), .Q (signal_4463) ) ;
    buf_clk cell_711 ( .C (clk), .D (signal_660), .Q (signal_4465) ) ;
    buf_clk cell_713 ( .C (clk), .D (signal_661), .Q (signal_4467) ) ;
    buf_clk cell_715 ( .C (clk), .D (signal_184), .Q (signal_4469) ) ;
    buf_clk cell_717 ( .C (clk), .D (signal_662), .Q (signal_4471) ) ;
    buf_clk cell_719 ( .C (clk), .D (signal_663), .Q (signal_4473) ) ;
    buf_clk cell_721 ( .C (clk), .D (signal_664), .Q (signal_4475) ) ;
    buf_clk cell_723 ( .C (clk), .D (signal_180), .Q (signal_4477) ) ;
    buf_clk cell_725 ( .C (clk), .D (signal_650), .Q (signal_4479) ) ;
    buf_clk cell_727 ( .C (clk), .D (signal_651), .Q (signal_4481) ) ;
    buf_clk cell_729 ( .C (clk), .D (signal_652), .Q (signal_4483) ) ;
    buf_clk cell_731 ( .C (clk), .D (signal_172), .Q (signal_4485) ) ;
    buf_clk cell_733 ( .C (clk), .D (signal_626), .Q (signal_4487) ) ;
    buf_clk cell_735 ( .C (clk), .D (signal_627), .Q (signal_4489) ) ;
    buf_clk cell_737 ( .C (clk), .D (signal_628), .Q (signal_4491) ) ;
    buf_clk cell_739 ( .C (clk), .D (signal_163), .Q (signal_4493) ) ;
    buf_clk cell_741 ( .C (clk), .D (signal_599), .Q (signal_4495) ) ;
    buf_clk cell_743 ( .C (clk), .D (signal_600), .Q (signal_4497) ) ;
    buf_clk cell_745 ( .C (clk), .D (signal_601), .Q (signal_4499) ) ;
    buf_clk cell_747 ( .C (clk), .D (signal_168), .Q (signal_4501) ) ;
    buf_clk cell_749 ( .C (clk), .D (signal_614), .Q (signal_4503) ) ;
    buf_clk cell_751 ( .C (clk), .D (signal_615), .Q (signal_4505) ) ;
    buf_clk cell_753 ( .C (clk), .D (signal_616), .Q (signal_4507) ) ;
    buf_clk cell_755 ( .C (clk), .D (signal_170), .Q (signal_4509) ) ;
    buf_clk cell_757 ( .C (clk), .D (signal_620), .Q (signal_4511) ) ;
    buf_clk cell_759 ( .C (clk), .D (signal_621), .Q (signal_4513) ) ;
    buf_clk cell_761 ( .C (clk), .D (signal_622), .Q (signal_4515) ) ;
    buf_clk cell_763 ( .C (clk), .D (signal_161), .Q (signal_4517) ) ;
    buf_clk cell_765 ( .C (clk), .D (signal_593), .Q (signal_4519) ) ;
    buf_clk cell_767 ( .C (clk), .D (signal_594), .Q (signal_4521) ) ;
    buf_clk cell_769 ( .C (clk), .D (signal_595), .Q (signal_4523) ) ;
    buf_clk cell_771 ( .C (clk), .D (signal_164), .Q (signal_4525) ) ;
    buf_clk cell_773 ( .C (clk), .D (signal_602), .Q (signal_4527) ) ;
    buf_clk cell_775 ( .C (clk), .D (signal_603), .Q (signal_4529) ) ;
    buf_clk cell_777 ( .C (clk), .D (signal_604), .Q (signal_4531) ) ;
    buf_clk cell_779 ( .C (clk), .D (signal_162), .Q (signal_4533) ) ;
    buf_clk cell_781 ( .C (clk), .D (signal_596), .Q (signal_4535) ) ;
    buf_clk cell_783 ( .C (clk), .D (signal_597), .Q (signal_4537) ) ;
    buf_clk cell_785 ( .C (clk), .D (signal_598), .Q (signal_4539) ) ;
    buf_clk cell_787 ( .C (clk), .D (signal_173), .Q (signal_4541) ) ;
    buf_clk cell_789 ( .C (clk), .D (signal_629), .Q (signal_4543) ) ;
    buf_clk cell_791 ( .C (clk), .D (signal_630), .Q (signal_4545) ) ;
    buf_clk cell_793 ( .C (clk), .D (signal_631), .Q (signal_4547) ) ;
    buf_clk cell_795 ( .C (clk), .D (signal_158), .Q (signal_4549) ) ;
    buf_clk cell_797 ( .C (clk), .D (signal_584), .Q (signal_4551) ) ;
    buf_clk cell_799 ( .C (clk), .D (signal_585), .Q (signal_4553) ) ;
    buf_clk cell_801 ( .C (clk), .D (signal_586), .Q (signal_4555) ) ;
    buf_clk cell_803 ( .C (clk), .D (signal_181), .Q (signal_4557) ) ;
    buf_clk cell_805 ( .C (clk), .D (signal_653), .Q (signal_4559) ) ;
    buf_clk cell_807 ( .C (clk), .D (signal_654), .Q (signal_4561) ) ;
    buf_clk cell_809 ( .C (clk), .D (signal_655), .Q (signal_4563) ) ;
    buf_clk cell_811 ( .C (clk), .D (signal_176), .Q (signal_4565) ) ;
    buf_clk cell_813 ( .C (clk), .D (signal_638), .Q (signal_4567) ) ;
    buf_clk cell_815 ( .C (clk), .D (signal_639), .Q (signal_4569) ) ;
    buf_clk cell_817 ( .C (clk), .D (signal_640), .Q (signal_4571) ) ;
    buf_clk cell_819 ( .C (clk), .D (signal_157), .Q (signal_4573) ) ;
    buf_clk cell_821 ( .C (clk), .D (signal_581), .Q (signal_4575) ) ;
    buf_clk cell_823 ( .C (clk), .D (signal_582), .Q (signal_4577) ) ;
    buf_clk cell_825 ( .C (clk), .D (signal_583), .Q (signal_4579) ) ;
    buf_clk cell_827 ( .C (clk), .D (signal_166), .Q (signal_4581) ) ;
    buf_clk cell_829 ( .C (clk), .D (signal_608), .Q (signal_4583) ) ;
    buf_clk cell_831 ( .C (clk), .D (signal_609), .Q (signal_4585) ) ;
    buf_clk cell_833 ( .C (clk), .D (signal_610), .Q (signal_4587) ) ;
    buf_clk cell_839 ( .C (clk), .D (signal_4592), .Q (signal_4593) ) ;
    buf_clk cell_847 ( .C (clk), .D (signal_4600), .Q (signal_4601) ) ;
    buf_clk cell_855 ( .C (clk), .D (signal_4608), .Q (signal_4609) ) ;
    buf_clk cell_863 ( .C (clk), .D (signal_4616), .Q (signal_4617) ) ;
    buf_clk cell_919 ( .C (clk), .D (signal_4672), .Q (signal_4673) ) ;
    buf_clk cell_929 ( .C (clk), .D (signal_4682), .Q (signal_4683) ) ;
    buf_clk cell_939 ( .C (clk), .D (signal_4692), .Q (signal_4693) ) ;
    buf_clk cell_949 ( .C (clk), .D (signal_4702), .Q (signal_4703) ) ;
    buf_clk cell_959 ( .C (clk), .D (signal_4712), .Q (signal_4713) ) ;
    buf_clk cell_971 ( .C (clk), .D (signal_4724), .Q (signal_4725) ) ;
    buf_clk cell_983 ( .C (clk), .D (signal_4736), .Q (signal_4737) ) ;
    buf_clk cell_995 ( .C (clk), .D (signal_4748), .Q (signal_4749) ) ;
    buf_clk cell_1007 ( .C (clk), .D (signal_4760), .Q (signal_4761) ) ;
    buf_clk cell_1021 ( .C (clk), .D (signal_4774), .Q (signal_4775) ) ;
    buf_clk cell_1035 ( .C (clk), .D (signal_4788), .Q (signal_4789) ) ;
    buf_clk cell_1049 ( .C (clk), .D (signal_4802), .Q (signal_4803) ) ;

    /* cells in depth 6 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_170 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({signal_667, signal_666, signal_665, signal_185}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_171 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({signal_670, signal_669, signal_668, signal_186}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_172 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({signal_673, signal_672, signal_671, signal_187}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_173 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({signal_676, signal_675, signal_674, signal_188}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_174 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({signal_679, signal_678, signal_677, signal_189}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_175 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4340, signal_4338, signal_4336, signal_4334}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({signal_682, signal_681, signal_680, signal_190}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_176 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4332, signal_4330, signal_4328, signal_4326}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({signal_685, signal_684, signal_683, signal_191}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_177 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4332, signal_4330, signal_4328, signal_4326}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({signal_688, signal_687, signal_686, signal_192}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_178 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({signal_691, signal_690, signal_689, signal_193}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_179 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({signal_694, signal_693, signal_692, signal_194}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_180 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_4356, signal_4354, signal_4352, signal_4350}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({signal_697, signal_696, signal_695, signal_195}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_181 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({signal_700, signal_699, signal_698, signal_196}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_182 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({signal_703, signal_702, signal_701, signal_197}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_183 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({signal_706, signal_705, signal_704, signal_198}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_184 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({signal_709, signal_708, signal_707, signal_199}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_185 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({signal_712, signal_711, signal_710, signal_200}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_186 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4340, signal_4338, signal_4336, signal_4334}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({signal_715, signal_714, signal_713, signal_201}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_187 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_583, signal_582, signal_581, signal_157}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({signal_718, signal_717, signal_716, signal_202}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_188 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({signal_721, signal_720, signal_719, signal_203}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_189 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_4356, signal_4354, signal_4352, signal_4350}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({signal_724, signal_723, signal_722, signal_204}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_190 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4340, signal_4338, signal_4336, signal_4334}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({signal_727, signal_726, signal_725, signal_205}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_191 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_4348, signal_4346, signal_4344, signal_4342}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({signal_730, signal_729, signal_728, signal_206}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_192 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_4348, signal_4346, signal_4344, signal_4342}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({signal_733, signal_732, signal_731, signal_207}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_193 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({signal_736, signal_735, signal_734, signal_208}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_194 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({signal_739, signal_738, signal_737, signal_209}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_195 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({signal_742, signal_741, signal_740, signal_210}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_196 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({signal_745, signal_744, signal_743, signal_211}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_197 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({signal_748, signal_747, signal_746, signal_212}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_198 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({signal_751, signal_750, signal_749, signal_213}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_199 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({signal_754, signal_753, signal_752, signal_214}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_200 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({signal_757, signal_756, signal_755, signal_215}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_201 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({signal_760, signal_759, signal_758, signal_216}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_202 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_607, signal_606, signal_605, signal_165}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({signal_763, signal_762, signal_761, signal_217}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_203 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({signal_766, signal_765, signal_764, signal_218}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_204 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({signal_769, signal_768, signal_767, signal_219}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_205 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({signal_772, signal_771, signal_770, signal_220}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_206 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({signal_775, signal_774, signal_773, signal_221}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_207 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({signal_778, signal_777, signal_776, signal_222}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_208 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_4356, signal_4354, signal_4352, signal_4350}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({signal_781, signal_780, signal_779, signal_223}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_209 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({signal_784, signal_783, signal_782, signal_224}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_210 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({signal_787, signal_786, signal_785, signal_225}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_211 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({signal_790, signal_789, signal_788, signal_226}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_212 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({signal_793, signal_792, signal_791, signal_227}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_213 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4332, signal_4330, signal_4328, signal_4326}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({signal_796, signal_795, signal_794, signal_228}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_214 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_583, signal_582, signal_581, signal_157}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({signal_799, signal_798, signal_797, signal_229}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_215 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({signal_802, signal_801, signal_800, signal_230}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_216 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({signal_805, signal_804, signal_803, signal_231}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_217 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({signal_808, signal_807, signal_806, signal_232}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_218 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({signal_811, signal_810, signal_809, signal_233}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_219 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({signal_814, signal_813, signal_812, signal_234}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_220 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({signal_817, signal_816, signal_815, signal_235}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_221 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({signal_820, signal_819, signal_818, signal_236}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_222 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({signal_823, signal_822, signal_821, signal_237}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_223 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({signal_826, signal_825, signal_824, signal_238}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_224 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({signal_829, signal_828, signal_827, signal_239}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_225 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({signal_832, signal_831, signal_830, signal_240}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_226 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({signal_835, signal_834, signal_833, signal_241}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_227 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_607, signal_606, signal_605, signal_165}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({signal_838, signal_837, signal_836, signal_242}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_228 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_4348, signal_4346, signal_4344, signal_4342}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({signal_841, signal_840, signal_839, signal_243}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_229 ( .s ({signal_4372, signal_4368, signal_4364, signal_4360}), .b ({signal_592, signal_591, signal_590, signal_160}), .a ({signal_640, signal_639, signal_638, signal_176}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({signal_847, signal_846, signal_845, signal_244}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_230 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({signal_850, signal_849, signal_848, signal_245}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_231 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({signal_853, signal_852, signal_851, signal_246}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_232 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({signal_856, signal_855, signal_854, signal_247}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_233 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({signal_859, signal_858, signal_857, signal_248}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_234 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({signal_862, signal_861, signal_860, signal_249}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_235 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({signal_865, signal_864, signal_863, signal_250}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_236 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({signal_868, signal_867, signal_866, signal_251}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_237 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({signal_871, signal_870, signal_869, signal_252}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_238 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({signal_874, signal_873, signal_872, signal_253}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_239 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_583, signal_582, signal_581, signal_157}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({signal_877, signal_876, signal_875, signal_254}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_240 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({signal_880, signal_879, signal_878, signal_255}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_241 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4340, signal_4338, signal_4336, signal_4334}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({signal_883, signal_882, signal_881, signal_256}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_242 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({signal_886, signal_885, signal_884, signal_257}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_243 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({signal_889, signal_888, signal_887, signal_258}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_244 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({signal_892, signal_891, signal_890, signal_259}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_245 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_4356, signal_4354, signal_4352, signal_4350}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({signal_895, signal_894, signal_893, signal_260}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_246 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({signal_898, signal_897, signal_896, signal_261}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_247 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({signal_901, signal_900, signal_899, signal_262}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_248 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_607, signal_606, signal_605, signal_165}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({signal_904, signal_903, signal_902, signal_263}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_249 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_583, signal_582, signal_581, signal_157}), .a ({signal_4348, signal_4346, signal_4344, signal_4342}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({signal_907, signal_906, signal_905, signal_264}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_250 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({signal_910, signal_909, signal_908, signal_265}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_251 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4332, signal_4330, signal_4328, signal_4326}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({signal_913, signal_912, signal_911, signal_266}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_252 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({signal_916, signal_915, signal_914, signal_267}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_253 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({signal_919, signal_918, signal_917, signal_268}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_254 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({signal_922, signal_921, signal_920, signal_269}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_255 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_607, signal_606, signal_605, signal_165}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({signal_925, signal_924, signal_923, signal_270}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_256 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({signal_928, signal_927, signal_926, signal_271}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_257 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_4340, signal_4338, signal_4336, signal_4334}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({signal_931, signal_930, signal_929, signal_272}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_258 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({signal_934, signal_933, signal_932, signal_273}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_259 ( .s ({signal_4372, signal_4368, signal_4364, signal_4360}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_604, signal_603, signal_602, signal_164}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({signal_937, signal_936, signal_935, signal_274}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_260 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_583, signal_582, signal_581, signal_157}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({signal_940, signal_939, signal_938, signal_275}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_261 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({signal_943, signal_942, signal_941, signal_276}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_262 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({signal_946, signal_945, signal_944, signal_277}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_263 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({signal_949, signal_948, signal_947, signal_278}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_264 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({signal_952, signal_951, signal_950, signal_279}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_265 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({1'b0, 1'b0, 1'b0, 1'b1}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({signal_955, signal_954, signal_953, signal_280}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_266 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({signal_958, signal_957, signal_956, signal_281}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_267 ( .s ({signal_4372, signal_4368, signal_4364, signal_4360}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_4380, signal_4378, signal_4376, signal_4374}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({signal_961, signal_960, signal_959, signal_282}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_268 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_583, signal_582, signal_581, signal_157}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({signal_964, signal_963, signal_962, signal_283}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_269 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({signal_967, signal_966, signal_965, signal_284}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_270 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({signal_970, signal_969, signal_968, signal_285}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_271 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({signal_973, signal_972, signal_971, signal_286}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_272 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({signal_976, signal_975, signal_974, signal_287}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_273 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4340, signal_4338, signal_4336, signal_4334}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({signal_979, signal_978, signal_977, signal_288}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_274 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({signal_982, signal_981, signal_980, signal_289}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_275 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({signal_985, signal_984, signal_983, signal_290}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_276 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_580, signal_579, signal_578, signal_156}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({signal_988, signal_987, signal_986, signal_291}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_277 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_607, signal_606, signal_605, signal_165}), .a ({signal_4348, signal_4346, signal_4344, signal_4342}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({signal_991, signal_990, signal_989, signal_292}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_278 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_583, signal_582, signal_581, signal_157}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({signal_994, signal_993, signal_992, signal_293}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_279 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({signal_997, signal_996, signal_995, signal_294}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_280 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({signal_1000, signal_999, signal_998, signal_295}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_281 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({signal_1003, signal_1002, signal_1001, signal_296}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_282 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({1'b0, 1'b0, 1'b0, 1'b0}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({signal_1006, signal_1005, signal_1004, signal_297}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_283 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({signal_1009, signal_1008, signal_1007, signal_298}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_284 ( .s ({signal_4372, signal_4368, signal_4364, signal_4360}), .b ({signal_658, signal_657, signal_656, signal_182}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({signal_1012, signal_1011, signal_1010, signal_299}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_285 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_643, signal_642, signal_641, signal_177}), .a ({signal_637, signal_636, signal_635, signal_175}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({signal_1015, signal_1014, signal_1013, signal_300}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_286 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({signal_1018, signal_1017, signal_1016, signal_301}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_287 ( .s ({signal_4372, signal_4368, signal_4364, signal_4360}), .b ({signal_589, signal_588, signal_587, signal_159}), .a ({signal_595, signal_594, signal_593, signal_161}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({signal_1021, signal_1020, signal_1019, signal_302}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_288 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({signal_1024, signal_1023, signal_1022, signal_303}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_289 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4332, signal_4330, signal_4328, signal_4326}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({signal_1027, signal_1026, signal_1025, signal_304}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_290 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_619, signal_618, signal_617, signal_169}), .a ({signal_4356, signal_4354, signal_4352, signal_4350}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({signal_1030, signal_1029, signal_1028, signal_305}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_291 ( .s ({signal_4372, signal_4368, signal_4364, signal_4360}), .b ({signal_649, signal_648, signal_647, signal_179}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({signal_1033, signal_1032, signal_1031, signal_306}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_292 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4356, signal_4354, signal_4352, signal_4350}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({signal_1036, signal_1035, signal_1034, signal_307}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_293 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_607, signal_606, signal_605, signal_165}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({signal_1039, signal_1038, signal_1037, signal_308}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_294 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_643, signal_642, signal_641, signal_177}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({signal_1042, signal_1041, signal_1040, signal_309}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_295 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_616, signal_615, signal_614, signal_168}), .a ({signal_598, signal_597, signal_596, signal_162}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({signal_1045, signal_1044, signal_1043, signal_310}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_296 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4332, signal_4330, signal_4328, signal_4326}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({signal_1048, signal_1047, signal_1046, signal_311}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_297 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_598, signal_597, signal_596, signal_162}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({signal_1051, signal_1050, signal_1049, signal_312}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_298 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_586, signal_585, signal_584, signal_158}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({signal_1054, signal_1053, signal_1052, signal_313}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_299 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4340, signal_4338, signal_4336, signal_4334}), .a ({signal_580, signal_579, signal_578, signal_156}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({signal_1057, signal_1056, signal_1055, signal_314}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_300 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_4348, signal_4346, signal_4344, signal_4342}), .a ({signal_586, signal_585, signal_584, signal_158}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({signal_1060, signal_1059, signal_1058, signal_315}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_301 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_634, signal_633, signal_632, signal_174}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({signal_1063, signal_1062, signal_1061, signal_316}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_302 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_634, signal_633, signal_632, signal_174}), .a ({signal_616, signal_615, signal_614, signal_168}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({signal_1066, signal_1065, signal_1064, signal_317}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_303 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_607, signal_606, signal_605, signal_165}), .a ({signal_619, signal_618, signal_617, signal_169}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({signal_1069, signal_1068, signal_1067, signal_318}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_304 ( .s ({signal_4324, signal_4322, signal_4320, signal_4318}), .b ({signal_637, signal_636, signal_635, signal_175}), .a ({signal_4332, signal_4330, signal_4328, signal_4326}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({signal_1072, signal_1071, signal_1070, signal_319}) ) ;
    buf_clk cell_628 ( .C (clk), .D (signal_4381), .Q (signal_4382) ) ;
    buf_clk cell_630 ( .C (clk), .D (signal_4383), .Q (signal_4384) ) ;
    buf_clk cell_632 ( .C (clk), .D (signal_4385), .Q (signal_4386) ) ;
    buf_clk cell_634 ( .C (clk), .D (signal_4387), .Q (signal_4388) ) ;
    buf_clk cell_636 ( .C (clk), .D (signal_4389), .Q (signal_4390) ) ;
    buf_clk cell_638 ( .C (clk), .D (signal_4391), .Q (signal_4392) ) ;
    buf_clk cell_640 ( .C (clk), .D (signal_4393), .Q (signal_4394) ) ;
    buf_clk cell_642 ( .C (clk), .D (signal_4395), .Q (signal_4396) ) ;
    buf_clk cell_644 ( .C (clk), .D (signal_4397), .Q (signal_4398) ) ;
    buf_clk cell_646 ( .C (clk), .D (signal_4399), .Q (signal_4400) ) ;
    buf_clk cell_648 ( .C (clk), .D (signal_4401), .Q (signal_4402) ) ;
    buf_clk cell_650 ( .C (clk), .D (signal_4403), .Q (signal_4404) ) ;
    buf_clk cell_652 ( .C (clk), .D (signal_4405), .Q (signal_4406) ) ;
    buf_clk cell_654 ( .C (clk), .D (signal_4407), .Q (signal_4408) ) ;
    buf_clk cell_656 ( .C (clk), .D (signal_4409), .Q (signal_4410) ) ;
    buf_clk cell_658 ( .C (clk), .D (signal_4411), .Q (signal_4412) ) ;
    buf_clk cell_660 ( .C (clk), .D (signal_4413), .Q (signal_4414) ) ;
    buf_clk cell_662 ( .C (clk), .D (signal_4415), .Q (signal_4416) ) ;
    buf_clk cell_664 ( .C (clk), .D (signal_4417), .Q (signal_4418) ) ;
    buf_clk cell_666 ( .C (clk), .D (signal_4419), .Q (signal_4420) ) ;
    buf_clk cell_668 ( .C (clk), .D (signal_4421), .Q (signal_4422) ) ;
    buf_clk cell_670 ( .C (clk), .D (signal_4423), .Q (signal_4424) ) ;
    buf_clk cell_672 ( .C (clk), .D (signal_4425), .Q (signal_4426) ) ;
    buf_clk cell_674 ( .C (clk), .D (signal_4427), .Q (signal_4428) ) ;
    buf_clk cell_676 ( .C (clk), .D (signal_4429), .Q (signal_4430) ) ;
    buf_clk cell_678 ( .C (clk), .D (signal_4431), .Q (signal_4432) ) ;
    buf_clk cell_680 ( .C (clk), .D (signal_4433), .Q (signal_4434) ) ;
    buf_clk cell_682 ( .C (clk), .D (signal_4435), .Q (signal_4436) ) ;
    buf_clk cell_684 ( .C (clk), .D (signal_4437), .Q (signal_4438) ) ;
    buf_clk cell_686 ( .C (clk), .D (signal_4439), .Q (signal_4440) ) ;
    buf_clk cell_688 ( .C (clk), .D (signal_4441), .Q (signal_4442) ) ;
    buf_clk cell_690 ( .C (clk), .D (signal_4443), .Q (signal_4444) ) ;
    buf_clk cell_692 ( .C (clk), .D (signal_4445), .Q (signal_4446) ) ;
    buf_clk cell_694 ( .C (clk), .D (signal_4447), .Q (signal_4448) ) ;
    buf_clk cell_696 ( .C (clk), .D (signal_4449), .Q (signal_4450) ) ;
    buf_clk cell_698 ( .C (clk), .D (signal_4451), .Q (signal_4452) ) ;
    buf_clk cell_700 ( .C (clk), .D (signal_4453), .Q (signal_4454) ) ;
    buf_clk cell_702 ( .C (clk), .D (signal_4455), .Q (signal_4456) ) ;
    buf_clk cell_704 ( .C (clk), .D (signal_4457), .Q (signal_4458) ) ;
    buf_clk cell_706 ( .C (clk), .D (signal_4459), .Q (signal_4460) ) ;
    buf_clk cell_708 ( .C (clk), .D (signal_4461), .Q (signal_4462) ) ;
    buf_clk cell_710 ( .C (clk), .D (signal_4463), .Q (signal_4464) ) ;
    buf_clk cell_712 ( .C (clk), .D (signal_4465), .Q (signal_4466) ) ;
    buf_clk cell_714 ( .C (clk), .D (signal_4467), .Q (signal_4468) ) ;
    buf_clk cell_716 ( .C (clk), .D (signal_4469), .Q (signal_4470) ) ;
    buf_clk cell_718 ( .C (clk), .D (signal_4471), .Q (signal_4472) ) ;
    buf_clk cell_720 ( .C (clk), .D (signal_4473), .Q (signal_4474) ) ;
    buf_clk cell_722 ( .C (clk), .D (signal_4475), .Q (signal_4476) ) ;
    buf_clk cell_724 ( .C (clk), .D (signal_4477), .Q (signal_4478) ) ;
    buf_clk cell_726 ( .C (clk), .D (signal_4479), .Q (signal_4480) ) ;
    buf_clk cell_728 ( .C (clk), .D (signal_4481), .Q (signal_4482) ) ;
    buf_clk cell_730 ( .C (clk), .D (signal_4483), .Q (signal_4484) ) ;
    buf_clk cell_732 ( .C (clk), .D (signal_4485), .Q (signal_4486) ) ;
    buf_clk cell_734 ( .C (clk), .D (signal_4487), .Q (signal_4488) ) ;
    buf_clk cell_736 ( .C (clk), .D (signal_4489), .Q (signal_4490) ) ;
    buf_clk cell_738 ( .C (clk), .D (signal_4491), .Q (signal_4492) ) ;
    buf_clk cell_740 ( .C (clk), .D (signal_4493), .Q (signal_4494) ) ;
    buf_clk cell_742 ( .C (clk), .D (signal_4495), .Q (signal_4496) ) ;
    buf_clk cell_744 ( .C (clk), .D (signal_4497), .Q (signal_4498) ) ;
    buf_clk cell_746 ( .C (clk), .D (signal_4499), .Q (signal_4500) ) ;
    buf_clk cell_748 ( .C (clk), .D (signal_4501), .Q (signal_4502) ) ;
    buf_clk cell_750 ( .C (clk), .D (signal_4503), .Q (signal_4504) ) ;
    buf_clk cell_752 ( .C (clk), .D (signal_4505), .Q (signal_4506) ) ;
    buf_clk cell_754 ( .C (clk), .D (signal_4507), .Q (signal_4508) ) ;
    buf_clk cell_756 ( .C (clk), .D (signal_4509), .Q (signal_4510) ) ;
    buf_clk cell_758 ( .C (clk), .D (signal_4511), .Q (signal_4512) ) ;
    buf_clk cell_760 ( .C (clk), .D (signal_4513), .Q (signal_4514) ) ;
    buf_clk cell_762 ( .C (clk), .D (signal_4515), .Q (signal_4516) ) ;
    buf_clk cell_764 ( .C (clk), .D (signal_4517), .Q (signal_4518) ) ;
    buf_clk cell_766 ( .C (clk), .D (signal_4519), .Q (signal_4520) ) ;
    buf_clk cell_768 ( .C (clk), .D (signal_4521), .Q (signal_4522) ) ;
    buf_clk cell_770 ( .C (clk), .D (signal_4523), .Q (signal_4524) ) ;
    buf_clk cell_772 ( .C (clk), .D (signal_4525), .Q (signal_4526) ) ;
    buf_clk cell_774 ( .C (clk), .D (signal_4527), .Q (signal_4528) ) ;
    buf_clk cell_776 ( .C (clk), .D (signal_4529), .Q (signal_4530) ) ;
    buf_clk cell_778 ( .C (clk), .D (signal_4531), .Q (signal_4532) ) ;
    buf_clk cell_780 ( .C (clk), .D (signal_4533), .Q (signal_4534) ) ;
    buf_clk cell_782 ( .C (clk), .D (signal_4535), .Q (signal_4536) ) ;
    buf_clk cell_784 ( .C (clk), .D (signal_4537), .Q (signal_4538) ) ;
    buf_clk cell_786 ( .C (clk), .D (signal_4539), .Q (signal_4540) ) ;
    buf_clk cell_788 ( .C (clk), .D (signal_4541), .Q (signal_4542) ) ;
    buf_clk cell_790 ( .C (clk), .D (signal_4543), .Q (signal_4544) ) ;
    buf_clk cell_792 ( .C (clk), .D (signal_4545), .Q (signal_4546) ) ;
    buf_clk cell_794 ( .C (clk), .D (signal_4547), .Q (signal_4548) ) ;
    buf_clk cell_796 ( .C (clk), .D (signal_4549), .Q (signal_4550) ) ;
    buf_clk cell_798 ( .C (clk), .D (signal_4551), .Q (signal_4552) ) ;
    buf_clk cell_800 ( .C (clk), .D (signal_4553), .Q (signal_4554) ) ;
    buf_clk cell_802 ( .C (clk), .D (signal_4555), .Q (signal_4556) ) ;
    buf_clk cell_804 ( .C (clk), .D (signal_4557), .Q (signal_4558) ) ;
    buf_clk cell_806 ( .C (clk), .D (signal_4559), .Q (signal_4560) ) ;
    buf_clk cell_808 ( .C (clk), .D (signal_4561), .Q (signal_4562) ) ;
    buf_clk cell_810 ( .C (clk), .D (signal_4563), .Q (signal_4564) ) ;
    buf_clk cell_812 ( .C (clk), .D (signal_4565), .Q (signal_4566) ) ;
    buf_clk cell_814 ( .C (clk), .D (signal_4567), .Q (signal_4568) ) ;
    buf_clk cell_816 ( .C (clk), .D (signal_4569), .Q (signal_4570) ) ;
    buf_clk cell_818 ( .C (clk), .D (signal_4571), .Q (signal_4572) ) ;
    buf_clk cell_820 ( .C (clk), .D (signal_4573), .Q (signal_4574) ) ;
    buf_clk cell_822 ( .C (clk), .D (signal_4575), .Q (signal_4576) ) ;
    buf_clk cell_824 ( .C (clk), .D (signal_4577), .Q (signal_4578) ) ;
    buf_clk cell_826 ( .C (clk), .D (signal_4579), .Q (signal_4580) ) ;
    buf_clk cell_828 ( .C (clk), .D (signal_4581), .Q (signal_4582) ) ;
    buf_clk cell_830 ( .C (clk), .D (signal_4583), .Q (signal_4584) ) ;
    buf_clk cell_832 ( .C (clk), .D (signal_4585), .Q (signal_4586) ) ;
    buf_clk cell_834 ( .C (clk), .D (signal_4587), .Q (signal_4588) ) ;
    buf_clk cell_840 ( .C (clk), .D (signal_4593), .Q (signal_4594) ) ;
    buf_clk cell_848 ( .C (clk), .D (signal_4601), .Q (signal_4602) ) ;
    buf_clk cell_856 ( .C (clk), .D (signal_4609), .Q (signal_4610) ) ;
    buf_clk cell_864 ( .C (clk), .D (signal_4617), .Q (signal_4618) ) ;
    buf_clk cell_920 ( .C (clk), .D (signal_4673), .Q (signal_4674) ) ;
    buf_clk cell_930 ( .C (clk), .D (signal_4683), .Q (signal_4684) ) ;
    buf_clk cell_940 ( .C (clk), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_950 ( .C (clk), .D (signal_4703), .Q (signal_4704) ) ;
    buf_clk cell_960 ( .C (clk), .D (signal_4713), .Q (signal_4714) ) ;
    buf_clk cell_972 ( .C (clk), .D (signal_4725), .Q (signal_4726) ) ;
    buf_clk cell_984 ( .C (clk), .D (signal_4737), .Q (signal_4738) ) ;
    buf_clk cell_996 ( .C (clk), .D (signal_4749), .Q (signal_4750) ) ;
    buf_clk cell_1008 ( .C (clk), .D (signal_4761), .Q (signal_4762) ) ;
    buf_clk cell_1022 ( .C (clk), .D (signal_4775), .Q (signal_4776) ) ;
    buf_clk cell_1036 ( .C (clk), .D (signal_4789), .Q (signal_4790) ) ;
    buf_clk cell_1050 ( .C (clk), .D (signal_4803), .Q (signal_4804) ) ;

    /* cells in depth 7 */
    buf_clk cell_841 ( .C (clk), .D (signal_4594), .Q (signal_4595) ) ;
    buf_clk cell_849 ( .C (clk), .D (signal_4602), .Q (signal_4603) ) ;
    buf_clk cell_857 ( .C (clk), .D (signal_4610), .Q (signal_4611) ) ;
    buf_clk cell_865 ( .C (clk), .D (signal_4618), .Q (signal_4619) ) ;
    buf_clk cell_867 ( .C (clk), .D (signal_282), .Q (signal_4621) ) ;
    buf_clk cell_869 ( .C (clk), .D (signal_959), .Q (signal_4623) ) ;
    buf_clk cell_871 ( .C (clk), .D (signal_960), .Q (signal_4625) ) ;
    buf_clk cell_873 ( .C (clk), .D (signal_961), .Q (signal_4627) ) ;
    buf_clk cell_875 ( .C (clk), .D (signal_274), .Q (signal_4629) ) ;
    buf_clk cell_877 ( .C (clk), .D (signal_935), .Q (signal_4631) ) ;
    buf_clk cell_879 ( .C (clk), .D (signal_936), .Q (signal_4633) ) ;
    buf_clk cell_881 ( .C (clk), .D (signal_937), .Q (signal_4635) ) ;
    buf_clk cell_883 ( .C (clk), .D (signal_306), .Q (signal_4637) ) ;
    buf_clk cell_885 ( .C (clk), .D (signal_1031), .Q (signal_4639) ) ;
    buf_clk cell_887 ( .C (clk), .D (signal_1032), .Q (signal_4641) ) ;
    buf_clk cell_889 ( .C (clk), .D (signal_1033), .Q (signal_4643) ) ;
    buf_clk cell_891 ( .C (clk), .D (signal_299), .Q (signal_4645) ) ;
    buf_clk cell_893 ( .C (clk), .D (signal_1010), .Q (signal_4647) ) ;
    buf_clk cell_895 ( .C (clk), .D (signal_1011), .Q (signal_4649) ) ;
    buf_clk cell_897 ( .C (clk), .D (signal_1012), .Q (signal_4651) ) ;
    buf_clk cell_899 ( .C (clk), .D (signal_244), .Q (signal_4653) ) ;
    buf_clk cell_901 ( .C (clk), .D (signal_845), .Q (signal_4655) ) ;
    buf_clk cell_903 ( .C (clk), .D (signal_846), .Q (signal_4657) ) ;
    buf_clk cell_905 ( .C (clk), .D (signal_847), .Q (signal_4659) ) ;
    buf_clk cell_907 ( .C (clk), .D (signal_302), .Q (signal_4661) ) ;
    buf_clk cell_909 ( .C (clk), .D (signal_1019), .Q (signal_4663) ) ;
    buf_clk cell_911 ( .C (clk), .D (signal_1020), .Q (signal_4665) ) ;
    buf_clk cell_913 ( .C (clk), .D (signal_1021), .Q (signal_4667) ) ;
    buf_clk cell_921 ( .C (clk), .D (signal_4674), .Q (signal_4675) ) ;
    buf_clk cell_931 ( .C (clk), .D (signal_4684), .Q (signal_4685) ) ;
    buf_clk cell_941 ( .C (clk), .D (signal_4694), .Q (signal_4695) ) ;
    buf_clk cell_951 ( .C (clk), .D (signal_4704), .Q (signal_4705) ) ;
    buf_clk cell_961 ( .C (clk), .D (signal_4714), .Q (signal_4715) ) ;
    buf_clk cell_973 ( .C (clk), .D (signal_4726), .Q (signal_4727) ) ;
    buf_clk cell_985 ( .C (clk), .D (signal_4738), .Q (signal_4739) ) ;
    buf_clk cell_997 ( .C (clk), .D (signal_4750), .Q (signal_4751) ) ;
    buf_clk cell_1009 ( .C (clk), .D (signal_4762), .Q (signal_4763) ) ;
    buf_clk cell_1023 ( .C (clk), .D (signal_4776), .Q (signal_4777) ) ;
    buf_clk cell_1037 ( .C (clk), .D (signal_4790), .Q (signal_4791) ) ;
    buf_clk cell_1051 ( .C (clk), .D (signal_4804), .Q (signal_4805) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_305 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4396, signal_4394, signal_4392, signal_4390}), .a ({signal_799, signal_798, signal_797, signal_229}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({signal_1075, signal_1074, signal_1073, signal_320}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_306 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1066, signal_1065, signal_1064, signal_317}), .a ({signal_817, signal_816, signal_815, signal_235}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({signal_1078, signal_1077, signal_1076, signal_321}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_307 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1027, signal_1026, signal_1025, signal_304}), .a ({signal_988, signal_987, signal_986, signal_291}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({signal_1081, signal_1080, signal_1079, signal_322}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_308 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1048, signal_1047, signal_1046, signal_311}), .a ({signal_4404, signal_4402, signal_4400, signal_4398}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({signal_1084, signal_1083, signal_1082, signal_323}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_309 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_751, signal_750, signal_749, signal_213}), .a ({signal_874, signal_873, signal_872, signal_253}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({signal_1087, signal_1086, signal_1085, signal_324}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_310 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_850, signal_849, signal_848, signal_245}), .a ({signal_1006, signal_1005, signal_1004, signal_297}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({signal_1090, signal_1089, signal_1088, signal_325}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_311 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({1'b0, 1'b0, 1'b0, 1'b1}), .a ({signal_670, signal_669, signal_668, signal_186}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({signal_1093, signal_1092, signal_1091, signal_326}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_312 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4412, signal_4410, signal_4408, signal_4406}), .a ({signal_913, signal_912, signal_911, signal_266}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({signal_1096, signal_1095, signal_1094, signal_327}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_313 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_709, signal_708, signal_707, signal_199}), .a ({signal_790, signal_789, signal_788, signal_226}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({signal_1099, signal_1098, signal_1097, signal_328}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_314 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_892, signal_891, signal_890, signal_259}), .a ({signal_979, signal_978, signal_977, signal_288}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({signal_1102, signal_1101, signal_1100, signal_329}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_315 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_985, signal_984, signal_983, signal_290}), .a ({signal_904, signal_903, signal_902, signal_263}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({signal_1105, signal_1104, signal_1103, signal_330}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_316 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_991, signal_990, signal_989, signal_292}), .a ({signal_1066, signal_1065, signal_1064, signal_317}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({signal_1108, signal_1107, signal_1106, signal_331}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_317 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_757, signal_756, signal_755, signal_215}), .a ({signal_4420, signal_4418, signal_4416, signal_4414}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({signal_1111, signal_1110, signal_1109, signal_332}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_318 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_778, signal_777, signal_776, signal_222}), .a ({signal_889, signal_888, signal_887, signal_258}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({signal_1114, signal_1113, signal_1112, signal_333}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_319 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_727, signal_726, signal_725, signal_205}), .a ({signal_4428, signal_4426, signal_4424, signal_4422}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({signal_1117, signal_1116, signal_1115, signal_334}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_320 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_826, signal_825, signal_824, signal_238}), .a ({signal_814, signal_813, signal_812, signal_234}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({signal_1120, signal_1119, signal_1118, signal_335}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_321 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_769, signal_768, signal_767, signal_219}), .a ({signal_751, signal_750, signal_749, signal_213}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({signal_1123, signal_1122, signal_1121, signal_336}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_322 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1060, signal_1059, signal_1058, signal_315}), .a ({signal_958, signal_957, signal_956, signal_281}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({signal_1126, signal_1125, signal_1124, signal_337}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_323 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_994, signal_993, signal_992, signal_293}), .a ({signal_718, signal_717, signal_716, signal_202}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({signal_1129, signal_1128, signal_1127, signal_338}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_324 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1054, signal_1053, signal_1052, signal_313}), .a ({signal_4436, signal_4434, signal_4432, signal_4430}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({signal_1132, signal_1131, signal_1130, signal_339}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_325 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_772, signal_771, signal_770, signal_220}), .a ({signal_799, signal_798, signal_797, signal_229}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({signal_1135, signal_1134, signal_1133, signal_340}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_326 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_841, signal_840, signal_839, signal_243}), .a ({signal_823, signal_822, signal_821, signal_237}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({signal_1138, signal_1137, signal_1136, signal_341}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_327 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_838, signal_837, signal_836, signal_242}), .a ({signal_982, signal_981, signal_980, signal_289}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({signal_1141, signal_1140, signal_1139, signal_342}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_328 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_760, signal_759, signal_758, signal_216}), .a ({signal_1063, signal_1062, signal_1061, signal_316}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({signal_1144, signal_1143, signal_1142, signal_343}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_329 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_823, signal_822, signal_821, signal_237}), .a ({signal_964, signal_963, signal_962, signal_283}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({signal_1147, signal_1146, signal_1145, signal_344}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_330 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1072, signal_1071, signal_1070, signal_319}), .a ({signal_862, signal_861, signal_860, signal_249}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({signal_1150, signal_1149, signal_1148, signal_345}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_331 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_880, signal_879, signal_878, signal_255}), .a ({signal_841, signal_840, signal_839, signal_243}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({signal_1153, signal_1152, signal_1151, signal_346}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_332 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_733, signal_732, signal_731, signal_207}), .a ({signal_4444, signal_4442, signal_4440, signal_4438}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({signal_1156, signal_1155, signal_1154, signal_347}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_333 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_925, signal_924, signal_923, signal_270}), .a ({signal_877, signal_876, signal_875, signal_254}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({signal_1159, signal_1158, signal_1157, signal_348}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_334 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_898, signal_897, signal_896, signal_261}), .a ({signal_1060, signal_1059, signal_1058, signal_315}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({signal_1162, signal_1161, signal_1160, signal_349}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_335 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4404, signal_4402, signal_4400, signal_4398}), .a ({signal_862, signal_861, signal_860, signal_249}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({signal_1165, signal_1164, signal_1163, signal_350}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_336 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_880, signal_879, signal_878, signal_255}), .a ({signal_955, signal_954, signal_953, signal_280}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({signal_1168, signal_1167, signal_1166, signal_351}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_337 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_808, signal_807, signal_806, signal_232}), .a ({signal_685, signal_684, signal_683, signal_191}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({signal_1171, signal_1170, signal_1169, signal_352}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_338 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1045, signal_1044, signal_1043, signal_310}), .a ({signal_991, signal_990, signal_989, signal_292}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({signal_1174, signal_1173, signal_1172, signal_353}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_339 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_859, signal_858, signal_857, signal_248}), .a ({signal_805, signal_804, signal_803, signal_231}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({signal_1177, signal_1176, signal_1175, signal_354}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_340 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1015, signal_1014, signal_1013, signal_300}), .a ({signal_1042, signal_1041, signal_1040, signal_309}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({signal_1180, signal_1179, signal_1178, signal_355}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_341 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_781, signal_780, signal_779, signal_223}), .a ({signal_970, signal_969, signal_968, signal_285}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({signal_1183, signal_1182, signal_1181, signal_356}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_342 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_826, signal_825, signal_824, signal_238}), .a ({signal_865, signal_864, signal_863, signal_250}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({signal_1186, signal_1185, signal_1184, signal_357}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_343 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_820, signal_819, signal_818, signal_236}), .a ({signal_4452, signal_4450, signal_4448, signal_4446}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({signal_1189, signal_1188, signal_1187, signal_358}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_344 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_931, signal_930, signal_929, signal_272}), .a ({signal_808, signal_807, signal_806, signal_232}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({signal_1192, signal_1191, signal_1190, signal_359}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_345 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4460, signal_4458, signal_4456, signal_4454}), .a ({signal_1027, signal_1026, signal_1025, signal_304}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({signal_1195, signal_1194, signal_1193, signal_360}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_346 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_958, signal_957, signal_956, signal_281}), .a ({signal_970, signal_969, signal_968, signal_285}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({signal_1198, signal_1197, signal_1196, signal_361}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_347 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_688, signal_687, signal_686, signal_192}), .a ({signal_862, signal_861, signal_860, signal_249}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({signal_1201, signal_1200, signal_1199, signal_362}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_348 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1009, signal_1008, signal_1007, signal_298}), .a ({signal_4468, signal_4466, signal_4464, signal_4462}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({signal_1204, signal_1203, signal_1202, signal_363}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_349 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_787, signal_786, signal_785, signal_225}), .a ({signal_4476, signal_4474, signal_4472, signal_4470}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({signal_1207, signal_1206, signal_1205, signal_364}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_350 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4444, signal_4442, signal_4440, signal_4438}), .a ({signal_976, signal_975, signal_974, signal_287}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({signal_1210, signal_1209, signal_1208, signal_365}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_351 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_784, signal_783, signal_782, signal_224}), .a ({signal_4484, signal_4482, signal_4480, signal_4478}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({signal_1213, signal_1212, signal_1211, signal_366}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_352 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_682, signal_681, signal_680, signal_190}), .a ({signal_4492, signal_4490, signal_4488, signal_4486}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({signal_1216, signal_1215, signal_1214, signal_367}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_353 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_886, signal_885, signal_884, signal_257}), .a ({signal_703, signal_702, signal_701, signal_197}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({signal_1219, signal_1218, signal_1217, signal_368}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_354 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4500, signal_4498, signal_4496, signal_4494}), .a ({signal_907, signal_906, signal_905, signal_264}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({signal_1222, signal_1221, signal_1220, signal_369}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_355 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_901, signal_900, signal_899, signal_262}), .a ({signal_4508, signal_4506, signal_4504, signal_4502}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({signal_1225, signal_1224, signal_1223, signal_370}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_356 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_679, signal_678, signal_677, signal_189}), .a ({signal_1039, signal_1038, signal_1037, signal_308}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({signal_1228, signal_1227, signal_1226, signal_371}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_357 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4396, signal_4394, signal_4392, signal_4390}), .a ({signal_865, signal_864, signal_863, signal_250}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({signal_1231, signal_1230, signal_1229, signal_372}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_358 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_910, signal_909, signal_908, signal_265}), .a ({signal_904, signal_903, signal_902, signal_263}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({signal_1234, signal_1233, signal_1232, signal_373}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_359 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_949, signal_948, signal_947, signal_278}), .a ({signal_829, signal_828, signal_827, signal_239}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({signal_1237, signal_1236, signal_1235, signal_374}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_360 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_673, signal_672, signal_671, signal_187}), .a ({signal_754, signal_753, signal_752, signal_214}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({signal_1240, signal_1239, signal_1238, signal_375}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_361 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_682, signal_681, signal_680, signal_190}), .a ({signal_700, signal_699, signal_698, signal_196}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({signal_1243, signal_1242, signal_1241, signal_376}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_362 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_964, signal_963, signal_962, signal_283}), .a ({signal_4516, signal_4514, signal_4512, signal_4510}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({signal_1246, signal_1245, signal_1244, signal_377}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_363 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_898, signal_897, signal_896, signal_261}), .a ({signal_1000, signal_999, signal_998, signal_295}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({signal_1249, signal_1248, signal_1247, signal_378}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_364 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_766, signal_765, signal_764, signal_218}), .a ({signal_676, signal_675, signal_674, signal_188}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({signal_1252, signal_1251, signal_1250, signal_379}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_365 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_967, signal_966, signal_965, signal_284}), .a ({signal_715, signal_714, signal_713, signal_201}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({signal_1255, signal_1254, signal_1253, signal_380}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_366 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4524, signal_4522, signal_4520, signal_4518}), .a ({signal_934, signal_933, signal_932, signal_273}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({signal_1258, signal_1257, signal_1256, signal_381}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_367 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4524, signal_4522, signal_4520, signal_4518}), .a ({signal_703, signal_702, signal_701, signal_197}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({signal_1261, signal_1260, signal_1259, signal_382}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_368 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_712, signal_711, signal_710, signal_200}), .a ({signal_4532, signal_4530, signal_4528, signal_4526}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({signal_1264, signal_1263, signal_1262, signal_383}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_369 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1024, signal_1023, signal_1022, signal_303}), .a ({signal_922, signal_921, signal_920, signal_269}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({signal_1267, signal_1266, signal_1265, signal_384}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_370 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_859, signal_858, signal_857, signal_248}), .a ({signal_883, signal_882, signal_881, signal_256}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({signal_1270, signal_1269, signal_1268, signal_385}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_371 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4516, signal_4514, signal_4512, signal_4510}), .a ({signal_898, signal_897, signal_896, signal_261}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({signal_1273, signal_1272, signal_1271, signal_386}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_372 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_817, signal_816, signal_815, signal_235}), .a ({signal_1030, signal_1029, signal_1028, signal_305}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({signal_1276, signal_1275, signal_1274, signal_387}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_373 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_787, signal_786, signal_785, signal_225}), .a ({signal_4484, signal_4482, signal_4480, signal_4478}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({signal_1279, signal_1278, signal_1277, signal_388}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_374 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_757, signal_756, signal_755, signal_215}), .a ({signal_4516, signal_4514, signal_4512, signal_4510}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({signal_1282, signal_1281, signal_1280, signal_389}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_375 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_856, signal_855, signal_854, signal_247}), .a ({signal_943, signal_942, signal_941, signal_276}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({signal_1285, signal_1284, signal_1283, signal_390}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_376 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_763, signal_762, signal_761, signal_217}), .a ({signal_769, signal_768, signal_767, signal_219}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({signal_1288, signal_1287, signal_1286, signal_391}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_377 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_775, signal_774, signal_773, signal_221}), .a ({signal_748, signal_747, signal_746, signal_212}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({signal_1291, signal_1290, signal_1289, signal_392}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_378 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4540, signal_4538, signal_4536, signal_4534}), .a ({signal_871, signal_870, signal_869, signal_252}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({signal_1294, signal_1293, signal_1292, signal_393}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_379 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_685, signal_684, signal_683, signal_191}), .a ({signal_721, signal_720, signal_719, signal_203}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({signal_1297, signal_1296, signal_1295, signal_394}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_380 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1006, signal_1005, signal_1004, signal_297}), .a ({signal_820, signal_819, signal_818, signal_236}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({signal_1300, signal_1299, signal_1298, signal_395}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_381 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_754, signal_753, signal_752, signal_214}), .a ({signal_4404, signal_4402, signal_4400, signal_4398}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({signal_1303, signal_1302, signal_1301, signal_396}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_382 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_877, signal_876, signal_875, signal_254}), .a ({signal_679, signal_678, signal_677, signal_189}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({signal_1306, signal_1305, signal_1304, signal_397}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_383 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_877, signal_876, signal_875, signal_254}), .a ({signal_769, signal_768, signal_767, signal_219}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({signal_1309, signal_1308, signal_1307, signal_398}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_384 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_742, signal_741, signal_740, signal_210}), .a ({signal_688, signal_687, signal_686, signal_192}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({signal_1312, signal_1311, signal_1310, signal_399}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_385 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_949, signal_948, signal_947, signal_278}), .a ({signal_916, signal_915, signal_914, signal_267}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({signal_1315, signal_1314, signal_1313, signal_400}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_386 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_748, signal_747, signal_746, signal_212}), .a ({signal_757, signal_756, signal_755, signal_215}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({signal_1318, signal_1317, signal_1316, signal_401}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_387 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1003, signal_1002, signal_1001, signal_296}), .a ({signal_928, signal_927, signal_926, signal_271}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({signal_1321, signal_1320, signal_1319, signal_402}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_388 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4548, signal_4546, signal_4544, signal_4542}), .a ({signal_691, signal_690, signal_689, signal_193}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({signal_1324, signal_1323, signal_1322, signal_403}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_389 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_739, signal_738, signal_737, signal_209}), .a ({signal_952, signal_951, signal_950, signal_279}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({signal_1327, signal_1326, signal_1325, signal_404}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_390 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_868, signal_867, signal_866, signal_251}), .a ({signal_1006, signal_1005, signal_1004, signal_297}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({signal_1330, signal_1329, signal_1328, signal_405}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_391 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_721, signal_720, signal_719, signal_203}), .a ({signal_4556, signal_4554, signal_4552, signal_4550}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({signal_1333, signal_1332, signal_1331, signal_406}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_392 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_841, signal_840, signal_839, signal_243}), .a ({signal_973, signal_972, signal_971, signal_286}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({signal_1336, signal_1335, signal_1334, signal_407}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_393 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_814, signal_813, signal_812, signal_234}), .a ({signal_4564, signal_4562, signal_4560, signal_4558}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({signal_1339, signal_1338, signal_1337, signal_408}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_394 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_997, signal_996, signal_995, signal_294}), .a ({signal_880, signal_879, signal_878, signal_255}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({signal_1342, signal_1341, signal_1340, signal_409}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_395 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_814, signal_813, signal_812, signal_234}), .a ({signal_919, signal_918, signal_917, signal_268}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({signal_1345, signal_1344, signal_1343, signal_410}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_396 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_835, signal_834, signal_833, signal_241}), .a ({signal_4516, signal_4514, signal_4512, signal_4510}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({signal_1348, signal_1347, signal_1346, signal_411}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_397 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_685, signal_684, signal_683, signal_191}), .a ({signal_811, signal_810, signal_809, signal_233}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({signal_1351, signal_1350, signal_1349, signal_412}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_398 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_904, signal_903, signal_902, signal_263}), .a ({signal_691, signal_690, signal_689, signal_193}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({signal_1354, signal_1353, signal_1352, signal_413}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_399 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1063, signal_1062, signal_1061, signal_316}), .a ({signal_769, signal_768, signal_767, signal_219}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({signal_1357, signal_1356, signal_1355, signal_414}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_400 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_802, signal_801, signal_800, signal_230}), .a ({signal_1051, signal_1050, signal_1049, signal_312}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({signal_1360, signal_1359, signal_1358, signal_415}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_401 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_946, signal_945, signal_944, signal_277}), .a ({signal_763, signal_762, signal_761, signal_217}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({signal_1363, signal_1362, signal_1361, signal_416}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_402 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1006, signal_1005, signal_1004, signal_297}), .a ({signal_1024, signal_1023, signal_1022, signal_303}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({signal_1366, signal_1365, signal_1364, signal_417}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_403 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1018, signal_1017, signal_1016, signal_301}), .a ({signal_940, signal_939, signal_938, signal_275}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({signal_1369, signal_1368, signal_1367, signal_418}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_404 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_907, signal_906, signal_905, signal_264}), .a ({signal_724, signal_723, signal_722, signal_204}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({signal_1372, signal_1371, signal_1370, signal_419}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_405 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_697, signal_696, signal_695, signal_195}), .a ({signal_778, signal_777, signal_776, signal_222}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({signal_1375, signal_1374, signal_1373, signal_420}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_406 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_796, signal_795, signal_794, signal_228}), .a ({signal_838, signal_837, signal_836, signal_242}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({signal_1378, signal_1377, signal_1376, signal_421}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_407 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_871, signal_870, signal_869, signal_252}), .a ({signal_1066, signal_1065, signal_1064, signal_317}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({signal_1381, signal_1380, signal_1379, signal_422}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_408 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_769, signal_768, signal_767, signal_219}), .a ({signal_673, signal_672, signal_671, signal_187}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({signal_1384, signal_1383, signal_1382, signal_423}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_409 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1006, signal_1005, signal_1004, signal_297}), .a ({signal_4428, signal_4426, signal_4424, signal_4422}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({signal_1387, signal_1386, signal_1385, signal_424}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_410 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_673, signal_672, signal_671, signal_187}), .a ({signal_4572, signal_4570, signal_4568, signal_4566}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({signal_1390, signal_1389, signal_1388, signal_425}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_411 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_682, signal_681, signal_680, signal_190}), .a ({signal_793, signal_792, signal_791, signal_227}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({signal_1393, signal_1392, signal_1391, signal_426}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_412 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_943, signal_942, signal_941, signal_276}), .a ({signal_4580, signal_4578, signal_4576, signal_4574}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({signal_1396, signal_1395, signal_1394, signal_427}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_413 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_838, signal_837, signal_836, signal_242}), .a ({signal_742, signal_741, signal_740, signal_210}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({signal_1399, signal_1398, signal_1397, signal_428}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_414 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_706, signal_705, signal_704, signal_198}), .a ({signal_733, signal_732, signal_731, signal_207}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({signal_1402, signal_1401, signal_1400, signal_429}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_415 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_907, signal_906, signal_905, signal_264}), .a ({signal_1069, signal_1068, signal_1067, signal_318}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({signal_1405, signal_1404, signal_1403, signal_430}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_416 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4572, signal_4570, signal_4568, signal_4566}), .a ({signal_931, signal_930, signal_929, signal_272}), .clk (clk), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({signal_1408, signal_1407, signal_1406, signal_431}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_417 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1009, signal_1008, signal_1007, signal_298}), .a ({signal_730, signal_729, signal_728, signal_206}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({signal_1411, signal_1410, signal_1409, signal_432}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_418 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_832, signal_831, signal_830, signal_240}), .a ({signal_667, signal_666, signal_665, signal_185}), .clk (clk), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({signal_1414, signal_1413, signal_1412, signal_433}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_419 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_985, signal_984, signal_983, signal_290}), .a ({signal_832, signal_831, signal_830, signal_240}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({signal_1417, signal_1416, signal_1415, signal_434}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_420 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1057, signal_1056, signal_1055, signal_314}), .a ({signal_751, signal_750, signal_749, signal_213}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({signal_1420, signal_1419, signal_1418, signal_435}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_421 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_895, signal_894, signal_893, signal_260}), .a ({signal_763, signal_762, signal_761, signal_217}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({signal_1423, signal_1422, signal_1421, signal_436}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_422 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_694, signal_693, signal_692, signal_194}), .a ({signal_829, signal_828, signal_827, signal_239}), .clk (clk), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({signal_1426, signal_1425, signal_1424, signal_437}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_423 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_745, signal_744, signal_743, signal_211}), .a ({signal_736, signal_735, signal_734, signal_208}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({signal_1429, signal_1428, signal_1427, signal_438}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_424 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_886, signal_885, signal_884, signal_257}), .a ({signal_742, signal_741, signal_740, signal_210}), .clk (clk), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({signal_1432, signal_1431, signal_1430, signal_439}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_425 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_4588, signal_4586, signal_4584, signal_4582}), .a ({signal_1000, signal_999, signal_998, signal_295}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({signal_1435, signal_1434, signal_1433, signal_440}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_426 ( .s ({signal_4388, signal_4386, signal_4384, signal_4382}), .b ({signal_1036, signal_1035, signal_1034, signal_307}), .a ({signal_853, signal_852, signal_851, signal_246}), .clk (clk), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({signal_1438, signal_1437, signal_1436, signal_441}) ) ;
    buf_clk cell_842 ( .C (clk), .D (signal_4595), .Q (signal_4596) ) ;
    buf_clk cell_850 ( .C (clk), .D (signal_4603), .Q (signal_4604) ) ;
    buf_clk cell_858 ( .C (clk), .D (signal_4611), .Q (signal_4612) ) ;
    buf_clk cell_866 ( .C (clk), .D (signal_4619), .Q (signal_4620) ) ;
    buf_clk cell_868 ( .C (clk), .D (signal_4621), .Q (signal_4622) ) ;
    buf_clk cell_870 ( .C (clk), .D (signal_4623), .Q (signal_4624) ) ;
    buf_clk cell_872 ( .C (clk), .D (signal_4625), .Q (signal_4626) ) ;
    buf_clk cell_874 ( .C (clk), .D (signal_4627), .Q (signal_4628) ) ;
    buf_clk cell_876 ( .C (clk), .D (signal_4629), .Q (signal_4630) ) ;
    buf_clk cell_878 ( .C (clk), .D (signal_4631), .Q (signal_4632) ) ;
    buf_clk cell_880 ( .C (clk), .D (signal_4633), .Q (signal_4634) ) ;
    buf_clk cell_882 ( .C (clk), .D (signal_4635), .Q (signal_4636) ) ;
    buf_clk cell_884 ( .C (clk), .D (signal_4637), .Q (signal_4638) ) ;
    buf_clk cell_886 ( .C (clk), .D (signal_4639), .Q (signal_4640) ) ;
    buf_clk cell_888 ( .C (clk), .D (signal_4641), .Q (signal_4642) ) ;
    buf_clk cell_890 ( .C (clk), .D (signal_4643), .Q (signal_4644) ) ;
    buf_clk cell_892 ( .C (clk), .D (signal_4645), .Q (signal_4646) ) ;
    buf_clk cell_894 ( .C (clk), .D (signal_4647), .Q (signal_4648) ) ;
    buf_clk cell_896 ( .C (clk), .D (signal_4649), .Q (signal_4650) ) ;
    buf_clk cell_898 ( .C (clk), .D (signal_4651), .Q (signal_4652) ) ;
    buf_clk cell_900 ( .C (clk), .D (signal_4653), .Q (signal_4654) ) ;
    buf_clk cell_902 ( .C (clk), .D (signal_4655), .Q (signal_4656) ) ;
    buf_clk cell_904 ( .C (clk), .D (signal_4657), .Q (signal_4658) ) ;
    buf_clk cell_906 ( .C (clk), .D (signal_4659), .Q (signal_4660) ) ;
    buf_clk cell_908 ( .C (clk), .D (signal_4661), .Q (signal_4662) ) ;
    buf_clk cell_910 ( .C (clk), .D (signal_4663), .Q (signal_4664) ) ;
    buf_clk cell_912 ( .C (clk), .D (signal_4665), .Q (signal_4666) ) ;
    buf_clk cell_914 ( .C (clk), .D (signal_4667), .Q (signal_4668) ) ;
    buf_clk cell_922 ( .C (clk), .D (signal_4675), .Q (signal_4676) ) ;
    buf_clk cell_932 ( .C (clk), .D (signal_4685), .Q (signal_4686) ) ;
    buf_clk cell_942 ( .C (clk), .D (signal_4695), .Q (signal_4696) ) ;
    buf_clk cell_952 ( .C (clk), .D (signal_4705), .Q (signal_4706) ) ;
    buf_clk cell_962 ( .C (clk), .D (signal_4715), .Q (signal_4716) ) ;
    buf_clk cell_974 ( .C (clk), .D (signal_4727), .Q (signal_4728) ) ;
    buf_clk cell_986 ( .C (clk), .D (signal_4739), .Q (signal_4740) ) ;
    buf_clk cell_998 ( .C (clk), .D (signal_4751), .Q (signal_4752) ) ;
    buf_clk cell_1010 ( .C (clk), .D (signal_4763), .Q (signal_4764) ) ;
    buf_clk cell_1024 ( .C (clk), .D (signal_4777), .Q (signal_4778) ) ;
    buf_clk cell_1038 ( .C (clk), .D (signal_4791), .Q (signal_4792) ) ;
    buf_clk cell_1052 ( .C (clk), .D (signal_4805), .Q (signal_4806) ) ;

    /* cells in depth 9 */
    buf_clk cell_923 ( .C (clk), .D (signal_4676), .Q (signal_4677) ) ;
    buf_clk cell_933 ( .C (clk), .D (signal_4686), .Q (signal_4687) ) ;
    buf_clk cell_943 ( .C (clk), .D (signal_4696), .Q (signal_4697) ) ;
    buf_clk cell_953 ( .C (clk), .D (signal_4706), .Q (signal_4707) ) ;
    buf_clk cell_963 ( .C (clk), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_975 ( .C (clk), .D (signal_4728), .Q (signal_4729) ) ;
    buf_clk cell_987 ( .C (clk), .D (signal_4740), .Q (signal_4741) ) ;
    buf_clk cell_999 ( .C (clk), .D (signal_4752), .Q (signal_4753) ) ;
    buf_clk cell_1011 ( .C (clk), .D (signal_4764), .Q (signal_4765) ) ;
    buf_clk cell_1025 ( .C (clk), .D (signal_4778), .Q (signal_4779) ) ;
    buf_clk cell_1039 ( .C (clk), .D (signal_4792), .Q (signal_4793) ) ;
    buf_clk cell_1053 ( .C (clk), .D (signal_4806), .Q (signal_4807) ) ;

    /* cells in depth 10 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_427 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1153, signal_1152, signal_1151, signal_346}), .a ({signal_1294, signal_1293, signal_1292, signal_393}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({signal_1444, signal_1443, signal_1442, signal_442}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_428 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1147, signal_1146, signal_1145, signal_344}), .a ({signal_1393, signal_1392, signal_1391, signal_426}), .clk (clk), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({signal_1447, signal_1446, signal_1445, signal_443}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_429 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1282, signal_1281, signal_1280, signal_389}), .a ({signal_1330, signal_1329, signal_1328, signal_405}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({signal_1450, signal_1449, signal_1448, signal_444}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_430 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1207, signal_1206, signal_1205, signal_364}), .a ({signal_1423, signal_1422, signal_1421, signal_436}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({signal_1453, signal_1452, signal_1451, signal_445}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_431 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1414, signal_1413, signal_1412, signal_433}), .a ({signal_1387, signal_1386, signal_1385, signal_424}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({signal_1456, signal_1455, signal_1454, signal_446}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_432 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1126, signal_1125, signal_1124, signal_337}), .a ({signal_1264, signal_1263, signal_1262, signal_383}), .clk (clk), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({signal_1459, signal_1458, signal_1457, signal_447}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_433 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1216, signal_1215, signal_1214, signal_367}), .a ({signal_1381, signal_1380, signal_1379, signal_422}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({signal_1462, signal_1461, signal_1460, signal_448}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_434 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1144, signal_1143, signal_1142, signal_343}), .a ({signal_1321, signal_1320, signal_1319, signal_402}), .clk (clk), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({signal_1465, signal_1464, signal_1463, signal_449}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_435 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1435, signal_1434, signal_1433, signal_440}), .a ({signal_1087, signal_1086, signal_1085, signal_324}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({signal_1468, signal_1467, signal_1466, signal_450}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_436 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1192, signal_1191, signal_1190, signal_359}), .a ({signal_1438, signal_1437, signal_1436, signal_441}), .clk (clk), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({signal_1471, signal_1470, signal_1469, signal_451}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_437 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1186, signal_1185, signal_1184, signal_357}), .a ({signal_1261, signal_1260, signal_1259, signal_382}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({signal_1474, signal_1473, signal_1472, signal_452}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_438 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1291, signal_1290, signal_1289, signal_392}), .a ({signal_1273, signal_1272, signal_1271, signal_386}), .clk (clk), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({signal_1477, signal_1476, signal_1475, signal_453}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_439 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1108, signal_1107, signal_1106, signal_331}), .a ({signal_1375, signal_1374, signal_1373, signal_420}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({signal_1480, signal_1479, signal_1478, signal_454}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_440 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1360, signal_1359, signal_1358, signal_415}), .a ({signal_1363, signal_1362, signal_1361, signal_416}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({signal_1483, signal_1482, signal_1481, signal_455}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_441 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1303, signal_1302, signal_1301, signal_396}), .a ({signal_4628, signal_4626, signal_4624, signal_4622}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({signal_1486, signal_1485, signal_1484, signal_456}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_442 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1420, signal_1419, signal_1418, signal_435}), .a ({signal_1372, signal_1371, signal_1370, signal_419}), .clk (clk), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({signal_1489, signal_1488, signal_1487, signal_457}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_443 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1084, signal_1083, signal_1082, signal_323}), .a ({signal_1159, signal_1158, signal_1157, signal_348}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({signal_1492, signal_1491, signal_1490, signal_458}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_444 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1312, signal_1311, signal_1310, signal_399}), .a ({signal_4636, signal_4634, signal_4632, signal_4630}), .clk (clk), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({signal_1495, signal_1494, signal_1493, signal_459}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_445 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1411, signal_1410, signal_1409, signal_432}), .a ({signal_4644, signal_4642, signal_4640, signal_4638}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({signal_1498, signal_1497, signal_1496, signal_460}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_446 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1252, signal_1251, signal_1250, signal_379}), .a ({signal_1093, signal_1092, signal_1091, signal_326}), .clk (clk), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({signal_1501, signal_1500, signal_1499, signal_461}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_447 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1219, signal_1218, signal_1217, signal_368}), .a ({signal_1168, signal_1167, signal_1166, signal_351}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({signal_1504, signal_1503, signal_1502, signal_462}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_448 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1117, signal_1116, signal_1115, signal_334}), .a ({signal_1237, signal_1236, signal_1235, signal_374}), .clk (clk), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({signal_1507, signal_1506, signal_1505, signal_463}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_449 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1351, signal_1350, signal_1349, signal_412}), .a ({signal_1090, signal_1089, signal_1088, signal_325}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({signal_1510, signal_1509, signal_1508, signal_464}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_450 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1198, signal_1197, signal_1196, signal_361}), .a ({signal_1318, signal_1317, signal_1316, signal_401}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({signal_1513, signal_1512, signal_1511, signal_465}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_451 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1096, signal_1095, signal_1094, signal_327}), .a ({signal_1105, signal_1104, signal_1103, signal_330}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({signal_1516, signal_1515, signal_1514, signal_466}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_452 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1075, signal_1074, signal_1073, signal_320}), .a ({signal_1150, signal_1149, signal_1148, signal_345}), .clk (clk), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({signal_1519, signal_1518, signal_1517, signal_467}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_453 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1339, signal_1338, signal_1337, signal_408}), .a ({signal_1429, signal_1428, signal_1427, signal_438}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({signal_1522, signal_1521, signal_1520, signal_468}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_454 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1405, signal_1404, signal_1403, signal_430}), .a ({signal_1366, signal_1365, signal_1364, signal_417}), .clk (clk), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({signal_1525, signal_1524, signal_1523, signal_469}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_455 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1357, signal_1356, signal_1355, signal_414}), .a ({signal_1135, signal_1134, signal_1133, signal_340}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({signal_1528, signal_1527, signal_1526, signal_470}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_456 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1228, signal_1227, signal_1226, signal_371}), .a ({signal_4652, signal_4650, signal_4648, signal_4646}), .clk (clk), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({signal_1531, signal_1530, signal_1529, signal_471}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_457 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1162, signal_1161, signal_1160, signal_349}), .a ({signal_1165, signal_1164, signal_1163, signal_350}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({signal_1534, signal_1533, signal_1532, signal_472}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_458 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1267, signal_1266, signal_1265, signal_384}), .a ({signal_1276, signal_1275, signal_1274, signal_387}), .clk (clk), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({signal_1537, signal_1536, signal_1535, signal_473}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_459 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1240, signal_1239, signal_1238, signal_375}), .a ({signal_1138, signal_1137, signal_1136, signal_341}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({signal_1540, signal_1539, signal_1538, signal_474}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_460 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1279, signal_1278, signal_1277, signal_388}), .a ({signal_1345, signal_1344, signal_1343, signal_410}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({signal_1543, signal_1542, signal_1541, signal_475}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_461 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1195, signal_1194, signal_1193, signal_360}), .a ({signal_1270, signal_1269, signal_1268, signal_385}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({signal_1546, signal_1545, signal_1544, signal_476}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_462 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1426, signal_1425, signal_1424, signal_437}), .a ({signal_1132, signal_1131, signal_1130, signal_339}), .clk (clk), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({signal_1549, signal_1548, signal_1547, signal_477}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_463 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1324, signal_1323, signal_1322, signal_403}), .a ({signal_1111, signal_1110, signal_1109, signal_332}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({signal_1552, signal_1551, signal_1550, signal_478}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_464 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1120, signal_1119, signal_1118, signal_335}), .a ({signal_1141, signal_1140, signal_1139, signal_342}), .clk (clk), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({signal_1555, signal_1554, signal_1553, signal_479}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_465 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1123, signal_1122, signal_1121, signal_336}), .a ({signal_1210, signal_1209, signal_1208, signal_365}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({signal_1558, signal_1557, signal_1556, signal_480}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_466 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1183, signal_1182, signal_1181, signal_356}), .a ({signal_1399, signal_1398, signal_1397, signal_428}), .clk (clk), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({signal_1561, signal_1560, signal_1559, signal_481}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_467 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1222, signal_1221, signal_1220, signal_369}), .a ({signal_1249, signal_1248, signal_1247, signal_378}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({signal_1564, signal_1563, signal_1562, signal_482}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_468 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1288, signal_1287, signal_1286, signal_391}), .a ({signal_1306, signal_1305, signal_1304, signal_397}), .clk (clk), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({signal_1567, signal_1566, signal_1565, signal_483}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_469 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1234, signal_1233, signal_1232, signal_373}), .a ({signal_1099, signal_1098, signal_1097, signal_328}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({signal_1570, signal_1569, signal_1568, signal_484}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_470 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1378, signal_1377, signal_1376, signal_421}), .a ({signal_1243, signal_1242, signal_1241, signal_376}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({signal_1573, signal_1572, signal_1571, signal_485}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_471 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1171, signal_1170, signal_1169, signal_352}), .a ({signal_1213, signal_1212, signal_1211, signal_366}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({signal_1576, signal_1575, signal_1574, signal_486}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_472 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1408, signal_1407, signal_1406, signal_431}), .a ({signal_1369, signal_1368, signal_1367, signal_418}), .clk (clk), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({signal_1579, signal_1578, signal_1577, signal_487}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_473 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1309, signal_1308, signal_1307, signal_398}), .a ({signal_1390, signal_1389, signal_1388, signal_425}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({signal_1582, signal_1581, signal_1580, signal_488}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_474 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1177, signal_1176, signal_1175, signal_354}), .a ({signal_1348, signal_1347, signal_1346, signal_411}), .clk (clk), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({signal_1585, signal_1584, signal_1583, signal_489}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_475 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1174, signal_1173, signal_1172, signal_353}), .a ({signal_1114, signal_1113, signal_1112, signal_333}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({signal_1588, signal_1587, signal_1586, signal_490}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_476 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1201, signal_1200, signal_1199, signal_362}), .a ({signal_1258, signal_1257, signal_1256, signal_381}), .clk (clk), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({signal_1591, signal_1590, signal_1589, signal_491}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_477 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1255, signal_1254, signal_1253, signal_380}), .a ({signal_1327, signal_1326, signal_1325, signal_404}), .clk (clk), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({signal_1594, signal_1593, signal_1592, signal_492}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_478 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_4660, signal_4658, signal_4656, signal_4654}), .a ({signal_1204, signal_1203, signal_1202, signal_363}), .clk (clk), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({signal_1597, signal_1596, signal_1595, signal_493}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_479 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1189, signal_1188, signal_1187, signal_358}), .a ({signal_1300, signal_1299, signal_1298, signal_395}), .clk (clk), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({signal_1600, signal_1599, signal_1598, signal_494}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_480 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1432, signal_1431, signal_1430, signal_439}), .a ({signal_1402, signal_1401, signal_1400, signal_429}), .clk (clk), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({signal_1603, signal_1602, signal_1601, signal_495}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_481 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1336, signal_1335, signal_1334, signal_407}), .a ({signal_1081, signal_1080, signal_1079, signal_322}), .clk (clk), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({signal_1606, signal_1605, signal_1604, signal_496}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_482 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1180, signal_1179, signal_1178, signal_355}), .a ({signal_1417, signal_1416, signal_1415, signal_434}), .clk (clk), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({signal_1609, signal_1608, signal_1607, signal_497}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_483 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1285, signal_1284, signal_1283, signal_390}), .a ({signal_1342, signal_1341, signal_1340, signal_409}), .clk (clk), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({signal_1612, signal_1611, signal_1610, signal_498}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_484 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1102, signal_1101, signal_1100, signal_329}), .a ({signal_1246, signal_1245, signal_1244, signal_377}), .clk (clk), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({signal_1615, signal_1614, signal_1613, signal_499}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_485 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1078, signal_1077, signal_1076, signal_321}), .a ({signal_1384, signal_1383, signal_1382, signal_423}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({signal_1618, signal_1617, signal_1616, signal_500}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_486 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1354, signal_1353, signal_1352, signal_413}), .a ({signal_1315, signal_1314, signal_1313, signal_400}), .clk (clk), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({signal_1621, signal_1620, signal_1619, signal_501}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_487 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1231, signal_1230, signal_1229, signal_372}), .a ({signal_1333, signal_1332, signal_1331, signal_406}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({signal_1624, signal_1623, signal_1622, signal_502}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_488 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_4668, signal_4666, signal_4664, signal_4662}), .a ({signal_1396, signal_1395, signal_1394, signal_427}), .clk (clk), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({signal_1627, signal_1626, signal_1625, signal_503}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_489 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1225, signal_1224, signal_1223, signal_370}), .a ({signal_1156, signal_1155, signal_1154, signal_347}), .clk (clk), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({signal_1630, signal_1629, signal_1628, signal_504}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_490 ( .s ({signal_4620, signal_4612, signal_4604, signal_4596}), .b ({signal_1297, signal_1296, signal_1295, signal_394}), .a ({signal_1129, signal_1128, signal_1127, signal_338}), .clk (clk), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({signal_1633, signal_1632, signal_1631, signal_505}) ) ;
    buf_clk cell_924 ( .C (clk), .D (signal_4677), .Q (signal_4678) ) ;
    buf_clk cell_934 ( .C (clk), .D (signal_4687), .Q (signal_4688) ) ;
    buf_clk cell_944 ( .C (clk), .D (signal_4697), .Q (signal_4698) ) ;
    buf_clk cell_954 ( .C (clk), .D (signal_4707), .Q (signal_4708) ) ;
    buf_clk cell_964 ( .C (clk), .D (signal_4717), .Q (signal_4718) ) ;
    buf_clk cell_976 ( .C (clk), .D (signal_4729), .Q (signal_4730) ) ;
    buf_clk cell_988 ( .C (clk), .D (signal_4741), .Q (signal_4742) ) ;
    buf_clk cell_1000 ( .C (clk), .D (signal_4753), .Q (signal_4754) ) ;
    buf_clk cell_1012 ( .C (clk), .D (signal_4765), .Q (signal_4766) ) ;
    buf_clk cell_1026 ( .C (clk), .D (signal_4779), .Q (signal_4780) ) ;
    buf_clk cell_1040 ( .C (clk), .D (signal_4793), .Q (signal_4794) ) ;
    buf_clk cell_1054 ( .C (clk), .D (signal_4807), .Q (signal_4808) ) ;

    /* cells in depth 11 */
    buf_clk cell_965 ( .C (clk), .D (signal_4718), .Q (signal_4719) ) ;
    buf_clk cell_977 ( .C (clk), .D (signal_4730), .Q (signal_4731) ) ;
    buf_clk cell_989 ( .C (clk), .D (signal_4742), .Q (signal_4743) ) ;
    buf_clk cell_1001 ( .C (clk), .D (signal_4754), .Q (signal_4755) ) ;
    buf_clk cell_1013 ( .C (clk), .D (signal_4766), .Q (signal_4767) ) ;
    buf_clk cell_1027 ( .C (clk), .D (signal_4780), .Q (signal_4781) ) ;
    buf_clk cell_1041 ( .C (clk), .D (signal_4794), .Q (signal_4795) ) ;
    buf_clk cell_1055 ( .C (clk), .D (signal_4808), .Q (signal_4809) ) ;

    /* cells in depth 12 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_491 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1543, signal_1542, signal_1541, signal_475}), .a ({signal_1450, signal_1449, signal_1448, signal_444}), .clk (clk), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({signal_1639, signal_1638, signal_1637, signal_506}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_492 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1468, signal_1467, signal_1466, signal_450}), .a ({signal_1483, signal_1482, signal_1481, signal_455}), .clk (clk), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({signal_1642, signal_1641, signal_1640, signal_507}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_493 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1585, signal_1584, signal_1583, signal_489}), .a ({signal_1528, signal_1527, signal_1526, signal_470}), .clk (clk), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({signal_1645, signal_1644, signal_1643, signal_508}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_494 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1567, signal_1566, signal_1565, signal_483}), .a ({signal_1453, signal_1452, signal_1451, signal_445}), .clk (clk), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({signal_1648, signal_1647, signal_1646, signal_509}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_495 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1615, signal_1614, signal_1613, signal_499}), .a ({signal_1489, signal_1488, signal_1487, signal_457}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({signal_1651, signal_1650, signal_1649, signal_510}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_496 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1558, signal_1557, signal_1556, signal_480}), .a ({signal_1552, signal_1551, signal_1550, signal_478}), .clk (clk), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({signal_1654, signal_1653, signal_1652, signal_511}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_497 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1621, signal_1620, signal_1619, signal_501}), .a ({signal_1546, signal_1545, signal_1544, signal_476}), .clk (clk), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({signal_1657, signal_1656, signal_1655, signal_512}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_498 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1588, signal_1587, signal_1586, signal_490}), .a ({signal_1522, signal_1521, signal_1520, signal_468}), .clk (clk), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({signal_1660, signal_1659, signal_1658, signal_513}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_499 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1627, signal_1626, signal_1625, signal_503}), .a ({signal_1501, signal_1500, signal_1499, signal_461}), .clk (clk), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({signal_1663, signal_1662, signal_1661, signal_514}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_500 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1492, signal_1491, signal_1490, signal_458}), .a ({signal_1504, signal_1503, signal_1502, signal_462}), .clk (clk), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({signal_1666, signal_1665, signal_1664, signal_515}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_501 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1465, signal_1464, signal_1463, signal_449}), .a ({signal_1519, signal_1518, signal_1517, signal_467}), .clk (clk), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({signal_1669, signal_1668, signal_1667, signal_516}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_502 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1612, signal_1611, signal_1610, signal_498}), .a ({signal_1591, signal_1590, signal_1589, signal_491}), .clk (clk), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({signal_1672, signal_1671, signal_1670, signal_517}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_503 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1474, signal_1473, signal_1472, signal_452}), .a ({signal_1582, signal_1581, signal_1580, signal_488}), .clk (clk), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({signal_1675, signal_1674, signal_1673, signal_518}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_504 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1594, signal_1593, signal_1592, signal_492}), .a ({signal_1525, signal_1524, signal_1523, signal_469}), .clk (clk), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({signal_1678, signal_1677, signal_1676, signal_519}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_505 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1603, signal_1602, signal_1601, signal_495}), .a ({signal_1534, signal_1533, signal_1532, signal_472}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({signal_1681, signal_1680, signal_1679, signal_520}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_506 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1606, signal_1605, signal_1604, signal_496}), .a ({signal_1510, signal_1509, signal_1508, signal_464}), .clk (clk), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({signal_1684, signal_1683, signal_1682, signal_521}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_507 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1600, signal_1599, signal_1598, signal_494}), .a ({signal_1498, signal_1497, signal_1496, signal_460}), .clk (clk), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({signal_1687, signal_1686, signal_1685, signal_522}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_508 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1537, signal_1536, signal_1535, signal_473}), .a ({signal_1609, signal_1608, signal_1607, signal_497}), .clk (clk), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({signal_1690, signal_1689, signal_1688, signal_523}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_509 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1597, signal_1596, signal_1595, signal_493}), .a ({signal_1495, signal_1494, signal_1493, signal_459}), .clk (clk), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({signal_1693, signal_1692, signal_1691, signal_524}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_510 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1480, signal_1479, signal_1478, signal_454}), .a ({signal_1624, signal_1623, signal_1622, signal_502}), .clk (clk), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({signal_1696, signal_1695, signal_1694, signal_525}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_511 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1630, signal_1629, signal_1628, signal_504}), .a ({signal_1555, signal_1554, signal_1553, signal_479}), .clk (clk), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({signal_1699, signal_1698, signal_1697, signal_526}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_512 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1486, signal_1485, signal_1484, signal_456}), .a ({signal_1459, signal_1458, signal_1457, signal_447}), .clk (clk), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({signal_1702, signal_1701, signal_1700, signal_527}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_513 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1456, signal_1455, signal_1454, signal_446}), .a ({signal_1516, signal_1515, signal_1514, signal_466}), .clk (clk), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({signal_1705, signal_1704, signal_1703, signal_528}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_514 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1531, signal_1530, signal_1529, signal_471}), .a ({signal_1573, signal_1572, signal_1571, signal_485}), .clk (clk), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({signal_1708, signal_1707, signal_1706, signal_529}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_515 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1564, signal_1563, signal_1562, signal_482}), .a ({signal_1471, signal_1470, signal_1469, signal_451}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({signal_1711, signal_1710, signal_1709, signal_530}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_516 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1462, signal_1461, signal_1460, signal_448}), .a ({signal_1507, signal_1506, signal_1505, signal_463}), .clk (clk), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({signal_1714, signal_1713, signal_1712, signal_531}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_517 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1513, signal_1512, signal_1511, signal_465}), .a ({signal_1633, signal_1632, signal_1631, signal_505}), .clk (clk), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({signal_1717, signal_1716, signal_1715, signal_532}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_518 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1477, signal_1476, signal_1475, signal_453}), .a ({signal_1618, signal_1617, signal_1616, signal_500}), .clk (clk), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({signal_1720, signal_1719, signal_1718, signal_533}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_519 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1540, signal_1539, signal_1538, signal_474}), .a ({signal_1561, signal_1560, signal_1559, signal_481}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({signal_1723, signal_1722, signal_1721, signal_534}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_520 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1549, signal_1548, signal_1547, signal_477}), .a ({signal_1570, signal_1569, signal_1568, signal_484}), .clk (clk), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({signal_1726, signal_1725, signal_1724, signal_535}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_521 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1579, signal_1578, signal_1577, signal_487}), .a ({signal_1444, signal_1443, signal_1442, signal_442}), .clk (clk), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({signal_1729, signal_1728, signal_1727, signal_536}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_522 ( .s ({signal_4708, signal_4698, signal_4688, signal_4678}), .b ({signal_1576, signal_1575, signal_1574, signal_486}), .a ({signal_1447, signal_1446, signal_1445, signal_443}), .clk (clk), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({signal_1732, signal_1731, signal_1730, signal_537}) ) ;
    buf_clk cell_966 ( .C (clk), .D (signal_4719), .Q (signal_4720) ) ;
    buf_clk cell_978 ( .C (clk), .D (signal_4731), .Q (signal_4732) ) ;
    buf_clk cell_990 ( .C (clk), .D (signal_4743), .Q (signal_4744) ) ;
    buf_clk cell_1002 ( .C (clk), .D (signal_4755), .Q (signal_4756) ) ;
    buf_clk cell_1014 ( .C (clk), .D (signal_4767), .Q (signal_4768) ) ;
    buf_clk cell_1028 ( .C (clk), .D (signal_4781), .Q (signal_4782) ) ;
    buf_clk cell_1042 ( .C (clk), .D (signal_4795), .Q (signal_4796) ) ;
    buf_clk cell_1056 ( .C (clk), .D (signal_4809), .Q (signal_4810) ) ;

    /* cells in depth 13 */
    buf_clk cell_1015 ( .C (clk), .D (signal_4768), .Q (signal_4769) ) ;
    buf_clk cell_1029 ( .C (clk), .D (signal_4782), .Q (signal_4783) ) ;
    buf_clk cell_1043 ( .C (clk), .D (signal_4796), .Q (signal_4797) ) ;
    buf_clk cell_1057 ( .C (clk), .D (signal_4810), .Q (signal_4811) ) ;

    /* cells in depth 14 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_523 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1714, signal_1713, signal_1712, signal_531}), .a ({signal_1675, signal_1674, signal_1673, signal_518}), .clk (clk), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({signal_1738, signal_1737, signal_1736, signal_538}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_524 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1645, signal_1644, signal_1643, signal_508}), .a ({signal_1726, signal_1725, signal_1724, signal_535}), .clk (clk), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({signal_1741, signal_1740, signal_1739, signal_539}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_525 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1693, signal_1692, signal_1691, signal_524}), .a ({signal_1690, signal_1689, signal_1688, signal_523}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({signal_1744, signal_1743, signal_1742, signal_540}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_526 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1678, signal_1677, signal_1676, signal_519}), .a ({signal_1702, signal_1701, signal_1700, signal_527}), .clk (clk), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({signal_1747, signal_1746, signal_1745, signal_541}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_527 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1705, signal_1704, signal_1703, signal_528}), .a ({signal_1639, signal_1638, signal_1637, signal_506}), .clk (clk), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({signal_1750, signal_1749, signal_1748, signal_542}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_528 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1699, signal_1698, signal_1697, signal_526}), .a ({signal_1732, signal_1731, signal_1730, signal_537}), .clk (clk), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({signal_1753, signal_1752, signal_1751, signal_543}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_529 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1651, signal_1650, signal_1649, signal_510}), .a ({signal_1720, signal_1719, signal_1718, signal_533}), .clk (clk), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({signal_1756, signal_1755, signal_1754, signal_544}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_530 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1642, signal_1641, signal_1640, signal_507}), .a ({signal_1654, signal_1653, signal_1652, signal_511}), .clk (clk), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({signal_1759, signal_1758, signal_1757, signal_545}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_531 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1663, signal_1662, signal_1661, signal_514}), .a ({signal_1669, signal_1668, signal_1667, signal_516}), .clk (clk), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({signal_1762, signal_1761, signal_1760, signal_546}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_532 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1681, signal_1680, signal_1679, signal_520}), .a ({signal_1696, signal_1695, signal_1694, signal_525}), .clk (clk), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({signal_1765, signal_1764, signal_1763, signal_547}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_533 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1657, signal_1656, signal_1655, signal_512}), .a ({signal_1711, signal_1710, signal_1709, signal_530}), .clk (clk), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({signal_1768, signal_1767, signal_1766, signal_548}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_534 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1666, signal_1665, signal_1664, signal_515}), .a ({signal_1723, signal_1722, signal_1721, signal_534}), .clk (clk), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({signal_1771, signal_1770, signal_1769, signal_549}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_535 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1684, signal_1683, signal_1682, signal_521}), .a ({signal_1672, signal_1671, signal_1670, signal_517}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({signal_1774, signal_1773, signal_1772, signal_550}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_536 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1708, signal_1707, signal_1706, signal_529}), .a ({signal_1729, signal_1728, signal_1727, signal_536}), .clk (clk), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({signal_1777, signal_1776, signal_1775, signal_551}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_537 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1660, signal_1659, signal_1658, signal_513}), .a ({signal_1717, signal_1716, signal_1715, signal_532}), .clk (clk), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({signal_1780, signal_1779, signal_1778, signal_552}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_538 ( .s ({signal_4756, signal_4744, signal_4732, signal_4720}), .b ({signal_1648, signal_1647, signal_1646, signal_509}), .a ({signal_1687, signal_1686, signal_1685, signal_522}), .clk (clk), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({signal_1783, signal_1782, signal_1781, signal_553}) ) ;
    buf_clk cell_1016 ( .C (clk), .D (signal_4769), .Q (signal_4770) ) ;
    buf_clk cell_1030 ( .C (clk), .D (signal_4783), .Q (signal_4784) ) ;
    buf_clk cell_1044 ( .C (clk), .D (signal_4797), .Q (signal_4798) ) ;
    buf_clk cell_1058 ( .C (clk), .D (signal_4811), .Q (signal_4812) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_539 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1741, signal_1740, signal_1739, signal_539}), .a ({signal_1759, signal_1758, signal_1757, signal_545}), .clk (clk), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({signal_1789, signal_1788, signal_1787, signal_145}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_540 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1768, signal_1767, signal_1766, signal_548}), .a ({signal_1762, signal_1761, signal_1760, signal_546}), .clk (clk), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({signal_1792, signal_1791, signal_1790, signal_148}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_541 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1753, signal_1752, signal_1751, signal_543}), .a ({signal_1765, signal_1764, signal_1763, signal_547}), .clk (clk), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({signal_1795, signal_1794, signal_1793, signal_143}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_542 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1783, signal_1782, signal_1781, signal_553}), .a ({signal_1777, signal_1776, signal_1775, signal_551}), .clk (clk), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({signal_1798, signal_1797, signal_1796, signal_146}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_543 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1744, signal_1743, signal_1742, signal_540}), .a ({signal_1780, signal_1779, signal_1778, signal_552}), .clk (clk), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({signal_1801, signal_1800, signal_1799, signal_149}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_544 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1774, signal_1773, signal_1772, signal_550}), .a ({signal_1750, signal_1749, signal_1748, signal_542}), .clk (clk), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({signal_1804, signal_1803, signal_1802, signal_144}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_545 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1738, signal_1737, signal_1736, signal_538}), .a ({signal_1771, signal_1770, signal_1769, signal_549}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({signal_1807, signal_1806, signal_1805, signal_147}) ) ;
    mux2_HPC2 #(.security_order(3), .pipeline(1)) cell_546 ( .s ({signal_4812, signal_4798, signal_4784, signal_4770}), .b ({signal_1756, signal_1755, signal_1754, signal_544}), .a ({signal_1747, signal_1746, signal_1745, signal_541}), .clk (clk), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({signal_1810, signal_1809, signal_1808, signal_150}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_1795, signal_1794, signal_1793, signal_143}), .Q ({Y_s3[7], Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_1804, signal_1803, signal_1802, signal_144}), .Q ({Y_s3[6], Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_1789, signal_1788, signal_1787, signal_145}), .Q ({Y_s3[5], Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_1798, signal_1797, signal_1796, signal_146}), .Q ({Y_s3[4], Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_1807, signal_1806, signal_1805, signal_147}), .Q ({Y_s3[3], Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_1792, signal_1791, signal_1790, signal_148}), .Q ({Y_s3[2], Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_1801, signal_1800, signal_1799, signal_149}), .Q ({Y_s3[1], Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_1810, signal_1809, signal_1808, signal_150}), .Q ({Y_s3[0], Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
