module Reg1(x, y);
 input [215:0] x;
 output [214:0] y;

  assign y[0] = x[215];
  assign y[135] = x[45];
  assign y[136] = x[46];
  assign y[137] = x[47];
  assign y[138] = x[48];
  assign y[139] = x[6];
  assign y[140] = x[7];
  assign y[141] = x[8];
  assign y[142] = x[9];
  assign y[143] = x[50];
  assign y[144] = x[51];
  assign y[145] = x[52];
  assign y[146] = x[53];
  assign y[147] = x[10];
  assign y[148] = x[11];
  assign y[149] = x[12];
  assign y[150] = x[13];
  assign y[151] = x[54];
  assign y[152] = x[55];
  assign y[153] = x[56];
  assign y[154] = x[57];
  assign y[155] = x[14];
  assign y[156] = x[15];
  assign y[157] = x[16];
  assign y[158] = x[17];
  assign y[159] = x[58];
  assign y[160] = x[59];
  assign y[161] = x[61];
  assign y[162] = x[62];
  assign y[163] = x[18];
  assign y[164] = x[19];
  assign y[165] = x[20];
  assign y[166] = x[21];
  assign y[167] = x[63];
  assign y[168] = x[64];
  assign y[169] = x[65];
  assign y[170] = x[66];
  assign y[171] = x[67];
  assign y[172] = x[68];
  assign y[173] = x[69];
  assign y[174] = x[70];
  assign y[175] = x[72];
  assign y[176] = x[73];
  assign y[177] = x[74];
  assign y[178] = x[75];
  assign y[179] = x[76];
  assign y[180] = x[77];
  assign y[181] = x[78];
  assign y[182] = x[79];
  assign y[183] = x[22];
  assign y[184] = x[23];
  assign y[185] = x[24];
  assign y[186] = x[25];
  assign y[187] = x[26];
  assign y[188] = x[27];
  assign y[189] = x[28];
  assign y[190] = x[29];
  assign y[191] = x[30];
  assign y[192] = x[31];
  assign y[193] = x[32];
  assign y[194] = x[33];
  assign y[195] = x[34];
  assign y[196] = x[35];
  assign y[197] = x[36];
  assign y[198] = x[37];
  assign y[199] = x[38];
  assign y[200] = x[49];
  assign y[201] = x[60];
  assign y[202] = x[71];
  assign y[203] = x[80];
  assign y[204] = x[81];
  assign y[205] = x[82];
  assign y[206] = x[83];
  assign y[207] = x[84];
  assign y[208] = x[85];
  assign y[209] = x[39];
  assign y[210] = x[40];
  assign y[211] = x[41];
  assign y[212] = x[42];
  assign y[213] = x[43];
  assign y[214] = x[44];
  register_stage #(.WIDTH(134)) inst_0(.clk(x[214]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[86],x[97],x[108],x[119],x[130],x[141],x[146],x[147],x[148],x[149],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[142],x[143],x[144],x[145],x[150],x[161],x[172],x[183],x[194],x[205],x[210],x[211],x[212],x[213],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[206],x[207],x[208],x[209]}), .Q({y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134]}));
endmodule

module Reg2(x, y);
 input [295:0] x;
 output [294:0] y;

  assign y[0] = x[291];
  assign y[1] = x[292];
  assign y[2] = x[293];
  assign y[3] = x[294];
  assign y[4] = x[295];
  assign y[195] = x[80];
  assign y[196] = x[81];
  assign y[197] = x[82];
  assign y[198] = x[83];
  assign y[199] = x[84];
  assign y[200] = x[30];
  assign y[201] = x[31];
  assign y[202] = x[32];
  assign y[203] = x[33];
  assign y[204] = x[34];
  assign y[205] = x[85];
  assign y[206] = x[86];
  assign y[207] = x[87];
  assign y[208] = x[88];
  assign y[209] = x[89];
  assign y[210] = x[35];
  assign y[211] = x[36];
  assign y[212] = x[37];
  assign y[213] = x[38];
  assign y[214] = x[39];
  assign y[215] = x[90];
  assign y[216] = x[91];
  assign y[217] = x[92];
  assign y[218] = x[93];
  assign y[219] = x[94];
  assign y[220] = x[40];
  assign y[221] = x[41];
  assign y[222] = x[42];
  assign y[223] = x[43];
  assign y[224] = x[44];
  assign y[225] = x[95];
  assign y[226] = x[96];
  assign y[227] = x[97];
  assign y[228] = x[98];
  assign y[229] = x[99];
  assign y[230] = x[45];
  assign y[231] = x[46];
  assign y[232] = x[47];
  assign y[233] = x[48];
  assign y[234] = x[49];
  assign y[235] = x[100];
  assign y[236] = x[101];
  assign y[237] = x[102];
  assign y[238] = x[103];
  assign y[239] = x[104];
  assign y[240] = x[105];
  assign y[241] = x[106];
  assign y[242] = x[107];
  assign y[243] = x[108];
  assign y[244] = x[109];
  assign y[245] = x[110];
  assign y[246] = x[111];
  assign y[247] = x[112];
  assign y[248] = x[113];
  assign y[249] = x[114];
  assign y[250] = x[115];
  assign y[251] = x[116];
  assign y[252] = x[117];
  assign y[253] = x[118];
  assign y[254] = x[119];
  assign y[255] = x[50];
  assign y[256] = x[51];
  assign y[257] = x[52];
  assign y[258] = x[53];
  assign y[259] = x[54];
  assign y[260] = x[55];
  assign y[261] = x[56];
  assign y[262] = x[57];
  assign y[263] = x[58];
  assign y[264] = x[59];
  assign y[265] = x[60];
  assign y[266] = x[61];
  assign y[267] = x[62];
  assign y[268] = x[63];
  assign y[269] = x[64];
  assign y[270] = x[65];
  assign y[271] = x[66];
  assign y[272] = x[67];
  assign y[273] = x[68];
  assign y[274] = x[69];
  assign y[275] = x[70];
  assign y[276] = x[71];
  assign y[277] = x[72];
  assign y[278] = x[73];
  assign y[279] = x[74];
  assign y[280] = x[120];
  assign y[281] = x[121];
  assign y[282] = x[122];
  assign y[283] = x[123];
  assign y[284] = x[124];
  assign y[285] = x[125];
  assign y[286] = x[126];
  assign y[287] = x[127];
  assign y[288] = x[128];
  assign y[289] = x[129];
  assign y[290] = x[75];
  assign y[291] = x[76];
  assign y[292] = x[77];
  assign y[293] = x[78];
  assign y[294] = x[79];
  register_stage #(.WIDTH(190)) inst_0(.clk(x[290]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[130],x[131],x[132],x[133],x[134],x[185],x[186],x[187],x[188],x[189],x[205],x[206],x[207],x[208],x[209],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[190],x[191],x[192],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[210],x[211],x[212],x[213],x[214],x[265],x[266],x[267],x[268],x[269],x[285],x[286],x[287],x[288],x[289],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[264],x[270],x[271],x[272],x[273],x[274],x[275],x[276],x[277],x[278],x[279],x[280],x[281],x[282],x[283],x[284]}), .Q({y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194]}));
endmodule

module InF(x, y);
 input [128:0] x;
 output [164:0] y;

  assign y[0] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y[1] = (1'b0);
  assign y[2] = (1'b0);
  assign y[3] = (1'b0);
  assign y[4] = (x[0]);
  assign y[5] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign y[6] = (x[4]);
  assign y[7] = (x[3]);
  assign y[8] = (x[2]);
  assign y[9] = (x[1]);
  assign y[10] = (x[5] & ~x[6] & ~x[7] & ~x[8]) | (~x[5] & x[6] & ~x[7] & ~x[8]) | (~x[5] & ~x[6] & x[7] & ~x[8]) | (~x[5] & ~x[6] & ~x[7] & x[8]) | (x[5] & x[6] & x[7] & ~x[8]) | (x[5] & x[6] & ~x[7] & x[8]) | (x[5] & ~x[6] & x[7] & x[8]) | (~x[5] & x[6] & x[7] & x[8]);
  assign y[11] = (x[8]);
  assign y[12] = (x[7]);
  assign y[13] = (x[6]);
  assign y[14] = (x[5]);
  assign y[15] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign y[16] = (x[12]);
  assign y[17] = (x[11]);
  assign y[18] = (x[10]);
  assign y[19] = (x[9]);
  assign y[20] = (x[13] & ~x[14] & ~x[15] & ~x[16]) | (~x[13] & x[14] & ~x[15] & ~x[16]) | (~x[13] & ~x[14] & x[15] & ~x[16]) | (~x[13] & ~x[14] & ~x[15] & x[16]) | (x[13] & x[14] & x[15] & ~x[16]) | (x[13] & x[14] & ~x[15] & x[16]) | (x[13] & ~x[14] & x[15] & x[16]) | (~x[13] & x[14] & x[15] & x[16]);
  assign y[21] = (x[16]);
  assign y[22] = (x[15]);
  assign y[23] = (x[14]);
  assign y[24] = (x[13]);
  assign y[25] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign y[26] = (x[20]);
  assign y[27] = (x[19]);
  assign y[28] = (x[18]);
  assign y[29] = (x[17]);
  assign y[30] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign y[31] = (x[24]);
  assign y[32] = (x[23]);
  assign y[33] = (x[22]);
  assign y[34] = (x[21]);
  assign y[35] = (x[25] & ~x[26] & ~x[27] & ~x[28]) | (~x[25] & x[26] & ~x[27] & ~x[28]) | (~x[25] & ~x[26] & x[27] & ~x[28]) | (~x[25] & ~x[26] & ~x[27] & x[28]) | (x[25] & x[26] & x[27] & ~x[28]) | (x[25] & x[26] & ~x[27] & x[28]) | (x[25] & ~x[26] & x[27] & x[28]) | (~x[25] & x[26] & x[27] & x[28]);
  assign y[36] = (x[28]);
  assign y[37] = (x[27]);
  assign y[38] = (x[26]);
  assign y[39] = (x[25]);
  assign y[40] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign y[41] = (x[32]);
  assign y[42] = (x[31]);
  assign y[43] = (x[30]);
  assign y[44] = (x[29]);
  assign y[45] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign y[46] = (x[36]);
  assign y[47] = (x[35]);
  assign y[48] = (x[34]);
  assign y[49] = (x[33]);
  assign y[50] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign y[51] = (x[40]);
  assign y[52] = (x[39]);
  assign y[53] = (x[38]);
  assign y[54] = (x[37]);
  assign y[55] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign y[56] = (x[44]);
  assign y[57] = (x[43]);
  assign y[58] = (x[42]);
  assign y[59] = (x[41]);
  assign y[60] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign y[61] = (x[48]);
  assign y[62] = (x[47]);
  assign y[63] = (x[46]);
  assign y[64] = (x[45]);
  assign y[65] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign y[66] = (x[52]);
  assign y[67] = (x[51]);
  assign y[68] = (x[50]);
  assign y[69] = (x[49]);
  assign y[70] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign y[71] = (x[56]);
  assign y[72] = (x[55]);
  assign y[73] = (x[54]);
  assign y[74] = (x[53]);
  assign y[75] = (x[57] & ~x[58] & ~x[59] & ~x[60]) | (~x[57] & x[58] & ~x[59] & ~x[60]) | (~x[57] & ~x[58] & x[59] & ~x[60]) | (~x[57] & ~x[58] & ~x[59] & x[60]) | (x[57] & x[58] & x[59] & ~x[60]) | (x[57] & x[58] & ~x[59] & x[60]) | (x[57] & ~x[58] & x[59] & x[60]) | (~x[57] & x[58] & x[59] & x[60]);
  assign y[76] = (x[60]);
  assign y[77] = (x[59]);
  assign y[78] = (x[58]);
  assign y[79] = (x[57]);
  assign y[80] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign y[81] = (x[64]);
  assign y[82] = (x[63]);
  assign y[83] = (x[62]);
  assign y[84] = (x[61]);
  assign y[85] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign y[86] = (x[68]);
  assign y[87] = (x[67]);
  assign y[88] = (x[66]);
  assign y[89] = (x[65]);
  assign y[90] = (x[69] & ~x[70] & ~x[71] & ~x[72]) | (~x[69] & x[70] & ~x[71] & ~x[72]) | (~x[69] & ~x[70] & x[71] & ~x[72]) | (~x[69] & ~x[70] & ~x[71] & x[72]) | (x[69] & x[70] & x[71] & ~x[72]) | (x[69] & x[70] & ~x[71] & x[72]) | (x[69] & ~x[70] & x[71] & x[72]) | (~x[69] & x[70] & x[71] & x[72]);
  assign y[91] = (x[72]);
  assign y[92] = (x[71]);
  assign y[93] = (x[70]);
  assign y[94] = (x[69]);
  assign y[95] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign y[96] = (x[76]);
  assign y[97] = (x[75]);
  assign y[98] = (x[74]);
  assign y[99] = (x[73]);
  assign y[100] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign y[101] = (x[80]);
  assign y[102] = (x[79]);
  assign y[103] = (x[78]);
  assign y[104] = (x[77]);
  assign y[105] = (x[81] & ~x[82] & ~x[83] & ~x[84]) | (~x[81] & x[82] & ~x[83] & ~x[84]) | (~x[81] & ~x[82] & x[83] & ~x[84]) | (~x[81] & ~x[82] & ~x[83] & x[84]) | (x[81] & x[82] & x[83] & ~x[84]) | (x[81] & x[82] & ~x[83] & x[84]) | (x[81] & ~x[82] & x[83] & x[84]) | (~x[81] & x[82] & x[83] & x[84]);
  assign y[106] = (x[84]);
  assign y[107] = (x[83]);
  assign y[108] = (x[82]);
  assign y[109] = (x[81]);
  assign y[110] = (x[85] & ~x[86] & ~x[87] & ~x[88]) | (~x[85] & x[86] & ~x[87] & ~x[88]) | (~x[85] & ~x[86] & x[87] & ~x[88]) | (~x[85] & ~x[86] & ~x[87] & x[88]) | (x[85] & x[86] & x[87] & ~x[88]) | (x[85] & x[86] & ~x[87] & x[88]) | (x[85] & ~x[86] & x[87] & x[88]) | (~x[85] & x[86] & x[87] & x[88]);
  assign y[111] = (x[88]);
  assign y[112] = (x[87]);
  assign y[113] = (x[86]);
  assign y[114] = (x[85]);
  assign y[115] = (x[89] & ~x[90] & ~x[91] & ~x[92]) | (~x[89] & x[90] & ~x[91] & ~x[92]) | (~x[89] & ~x[90] & x[91] & ~x[92]) | (~x[89] & ~x[90] & ~x[91] & x[92]) | (x[89] & x[90] & x[91] & ~x[92]) | (x[89] & x[90] & ~x[91] & x[92]) | (x[89] & ~x[90] & x[91] & x[92]) | (~x[89] & x[90] & x[91] & x[92]);
  assign y[116] = (x[92]);
  assign y[117] = (x[91]);
  assign y[118] = (x[90]);
  assign y[119] = (x[89]);
  assign y[120] = (x[93] & ~x[94] & ~x[95] & ~x[96]) | (~x[93] & x[94] & ~x[95] & ~x[96]) | (~x[93] & ~x[94] & x[95] & ~x[96]) | (~x[93] & ~x[94] & ~x[95] & x[96]) | (x[93] & x[94] & x[95] & ~x[96]) | (x[93] & x[94] & ~x[95] & x[96]) | (x[93] & ~x[94] & x[95] & x[96]) | (~x[93] & x[94] & x[95] & x[96]);
  assign y[121] = (x[96]);
  assign y[122] = (x[95]);
  assign y[123] = (x[94]);
  assign y[124] = (x[93]);
  assign y[125] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign y[126] = (x[100]);
  assign y[127] = (x[99]);
  assign y[128] = (x[98]);
  assign y[129] = (x[97]);
  assign y[130] = (x[101] & ~x[102] & ~x[103] & ~x[104]) | (~x[101] & x[102] & ~x[103] & ~x[104]) | (~x[101] & ~x[102] & x[103] & ~x[104]) | (~x[101] & ~x[102] & ~x[103] & x[104]) | (x[101] & x[102] & x[103] & ~x[104]) | (x[101] & x[102] & ~x[103] & x[104]) | (x[101] & ~x[102] & x[103] & x[104]) | (~x[101] & x[102] & x[103] & x[104]);
  assign y[131] = (x[104]);
  assign y[132] = (x[103]);
  assign y[133] = (x[102]);
  assign y[134] = (x[101]);
  assign y[135] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign y[136] = (x[108]);
  assign y[137] = (x[107]);
  assign y[138] = (x[106]);
  assign y[139] = (x[105]);
  assign y[140] = (x[109] & ~x[110] & ~x[111] & ~x[112]) | (~x[109] & x[110] & ~x[111] & ~x[112]) | (~x[109] & ~x[110] & x[111] & ~x[112]) | (~x[109] & ~x[110] & ~x[111] & x[112]) | (x[109] & x[110] & x[111] & ~x[112]) | (x[109] & x[110] & ~x[111] & x[112]) | (x[109] & ~x[110] & x[111] & x[112]) | (~x[109] & x[110] & x[111] & x[112]);
  assign y[141] = (x[112]);
  assign y[142] = (x[111]);
  assign y[143] = (x[110]);
  assign y[144] = (x[109]);
  assign y[145] = (x[113] & ~x[114] & ~x[115] & ~x[116]) | (~x[113] & x[114] & ~x[115] & ~x[116]) | (~x[113] & ~x[114] & x[115] & ~x[116]) | (~x[113] & ~x[114] & ~x[115] & x[116]) | (x[113] & x[114] & x[115] & ~x[116]) | (x[113] & x[114] & ~x[115] & x[116]) | (x[113] & ~x[114] & x[115] & x[116]) | (~x[113] & x[114] & x[115] & x[116]);
  assign y[146] = (x[116]);
  assign y[147] = (x[115]);
  assign y[148] = (x[114]);
  assign y[149] = (x[113]);
  assign y[150] = (x[117] & ~x[118] & ~x[119] & ~x[120]) | (~x[117] & x[118] & ~x[119] & ~x[120]) | (~x[117] & ~x[118] & x[119] & ~x[120]) | (~x[117] & ~x[118] & ~x[119] & x[120]) | (x[117] & x[118] & x[119] & ~x[120]) | (x[117] & x[118] & ~x[119] & x[120]) | (x[117] & ~x[118] & x[119] & x[120]) | (~x[117] & x[118] & x[119] & x[120]);
  assign y[151] = (x[120]);
  assign y[152] = (x[119]);
  assign y[153] = (x[118]);
  assign y[154] = (x[117]);
  assign y[155] = (x[121] & ~x[122] & ~x[123] & ~x[124]) | (~x[121] & x[122] & ~x[123] & ~x[124]) | (~x[121] & ~x[122] & x[123] & ~x[124]) | (~x[121] & ~x[122] & ~x[123] & x[124]) | (x[121] & x[122] & x[123] & ~x[124]) | (x[121] & x[122] & ~x[123] & x[124]) | (x[121] & ~x[122] & x[123] & x[124]) | (~x[121] & x[122] & x[123] & x[124]);
  assign y[156] = (x[124]);
  assign y[157] = (x[123]);
  assign y[158] = (x[122]);
  assign y[159] = (x[121]);
  assign y[160] = (x[125] & ~x[126] & ~x[127] & ~x[128]) | (~x[125] & x[126] & ~x[127] & ~x[128]) | (~x[125] & ~x[126] & x[127] & ~x[128]) | (~x[125] & ~x[126] & ~x[127] & x[128]) | (x[125] & x[126] & x[127] & ~x[128]) | (x[125] & x[126] & ~x[127] & x[128]) | (x[125] & ~x[126] & x[127] & x[128]) | (~x[125] & x[126] & x[127] & x[128]);
  assign y[161] = (x[128]);
  assign y[162] = (x[127]);
  assign y[163] = (x[126]);
  assign y[164] = (x[125]);
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [308:0] x;
 output [173:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx29 Fx29_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx30 Fx30_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx34 Fx34_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx35 Fx35_inst(.x({x[25], x[24], x[23], x[22], x[21]}), .y(y[14]));
  Fx36 Fx36_inst(.x({x[26], x[24]}), .y(y[15]));
  Fx37 Fx37_inst(.x({x[27], x[23]}), .y(y[16]));
  Fx38 Fx38_inst(.x({x[28], x[22]}), .y(y[17]));
  Fx39 Fx39_inst(.x({x[29], x[21]}), .y(y[18]));
  Fx40 Fx40_inst(.x({x[34], x[33], x[32], x[31], x[30]}), .y(y[19]));
  Fx41 Fx41_inst(.x({x[35], x[33]}), .y(y[20]));
  Fx42 Fx42_inst(.x({x[36], x[32]}), .y(y[21]));
  Fx43 Fx43_inst(.x({x[37], x[31]}), .y(y[22]));
  Fx44 Fx44_inst(.x({x[38], x[30]}), .y(y[23]));
  Fx45 Fx45_inst(.x({x[43], x[42], x[41], x[40], x[39]}), .y(y[24]));
  Fx46 Fx46_inst(.x({x[44], x[42]}), .y(y[25]));
  Fx47 Fx47_inst(.x({x[45], x[41]}), .y(y[26]));
  Fx48 Fx48_inst(.x({x[46], x[40]}), .y(y[27]));
  Fx49 Fx49_inst(.x({x[47], x[39]}), .y(y[28]));
  Fx50 Fx50_inst(.x({x[52], x[51], x[50], x[49], x[48]}), .y(y[29]));
  Fx51 Fx51_inst(.x({x[53], x[51]}), .y(y[30]));
  Fx52 Fx52_inst(.x({x[54], x[50]}), .y(y[31]));
  Fx53 Fx53_inst(.x({x[55], x[49]}), .y(y[32]));
  Fx54 Fx54_inst(.x({x[56], x[48]}), .y(y[33]));
  Fx55 Fx55_inst(.x({x[61], x[60], x[59], x[58], x[57]}), .y(y[34]));
  Fx56 Fx56_inst(.x({x[62], x[60]}), .y(y[35]));
  Fx57 Fx57_inst(.x({x[63], x[59]}), .y(y[36]));
  Fx58 Fx58_inst(.x({x[64], x[58]}), .y(y[37]));
  Fx59 Fx59_inst(.x({x[65], x[57]}), .y(y[38]));
  Fx60 Fx60_inst(.x({x[70], x[69], x[68], x[67], x[66]}), .y(y[39]));
  Fx61 Fx61_inst(.x({x[71], x[69]}), .y(y[40]));
  Fx62 Fx62_inst(.x({x[72], x[68]}), .y(y[41]));
  Fx63 Fx63_inst(.x({x[73], x[67]}), .y(y[42]));
  Fx64 Fx64_inst(.x({x[74], x[66]}), .y(y[43]));
  Fx65 Fx65_inst(.x({x[79], x[78], x[77], x[76], x[75]}), .y(y[44]));
  Fx66 Fx66_inst(.x({x[80], x[78]}), .y(y[45]));
  Fx67 Fx67_inst(.x({x[81], x[77]}), .y(y[46]));
  Fx68 Fx68_inst(.x({x[82], x[76]}), .y(y[47]));
  Fx69 Fx69_inst(.x({x[83], x[75]}), .y(y[48]));
  Fx70 Fx70_inst(.x({x[88], x[87], x[86], x[85], x[84]}), .y(y[49]));
  Fx71 Fx71_inst(.x({x[89], x[87]}), .y(y[50]));
  Fx72 Fx72_inst(.x({x[90], x[86]}), .y(y[51]));
  Fx73 Fx73_inst(.x({x[91], x[85]}), .y(y[52]));
  Fx74 Fx74_inst(.x({x[92], x[84]}), .y(y[53]));
  Fx75 Fx75_inst(.x({x[97], x[96], x[95], x[94], x[93]}), .y(y[54]));
  Fx76 Fx76_inst(.x({x[98], x[96]}), .y(y[55]));
  Fx77 Fx77_inst(.x({x[99], x[95]}), .y(y[56]));
  Fx78 Fx78_inst(.x({x[100], x[94]}), .y(y[57]));
  Fx79 Fx79_inst(.x({x[101], x[93]}), .y(y[58]));
  Fx80 Fx80_inst(.x({x[106], x[105], x[104], x[103], x[102]}), .y(y[59]));
  Fx81 Fx81_inst(.x({x[107], x[105]}), .y(y[60]));
  Fx82 Fx82_inst(.x({x[108], x[104]}), .y(y[61]));
  Fx83 Fx83_inst(.x({x[109], x[103]}), .y(y[62]));
  Fx84 Fx84_inst(.x({x[110], x[102]}), .y(y[63]));
  Fx85 Fx85_inst(.x({x[115], x[114], x[113], x[112], x[111]}), .y(y[64]));
  Fx86 Fx86_inst(.x({x[116], x[114]}), .y(y[65]));
  Fx87 Fx87_inst(.x({x[117], x[113]}), .y(y[66]));
  Fx88 Fx88_inst(.x({x[118], x[112]}), .y(y[67]));
  Fx89 Fx89_inst(.x({x[119], x[111]}), .y(y[68]));
  Fx90 Fx90_inst(.x({x[124], x[123], x[122], x[121], x[120]}), .y(y[69]));
  Fx91 Fx91_inst(.x({x[125], x[123]}), .y(y[70]));
  Fx92 Fx92_inst(.x({x[126], x[122]}), .y(y[71]));
  Fx93 Fx93_inst(.x({x[127], x[121]}), .y(y[72]));
  Fx94 Fx94_inst(.x({x[128], x[120]}), .y(y[73]));
  Fx95 Fx95_inst(.x({x[133], x[132], x[131], x[130], x[129]}), .y(y[74]));
  Fx96 Fx96_inst(.x({x[134], x[132]}), .y(y[75]));
  Fx97 Fx97_inst(.x({x[135], x[131]}), .y(y[76]));
  Fx98 Fx98_inst(.x({x[136], x[130]}), .y(y[77]));
  Fx99 Fx99_inst(.x({x[137], x[129]}), .y(y[78]));
  Fx100 Fx100_inst(.x({x[142], x[141], x[140], x[139], x[138]}), .y(y[79]));
  Fx101 Fx101_inst(.x({x[143], x[141]}), .y(y[80]));
  Fx102 Fx102_inst(.x({x[144], x[140]}), .y(y[81]));
  Fx103 Fx103_inst(.x({x[145], x[139]}), .y(y[82]));
  Fx104 Fx104_inst(.x({x[146], x[138]}), .y(y[83]));
  Fx105 Fx105_inst(.x({x[151], x[150], x[149], x[148], x[147]}), .y(y[84]));
  Fx106 Fx106_inst(.x({x[152], x[150]}), .y(y[85]));
  Fx107 Fx107_inst(.x({x[153], x[149]}), .y(y[86]));
  Fx108 Fx108_inst(.x({x[154], x[148]}), .y(y[87]));
  Fx109 Fx109_inst(.x({x[155], x[147]}), .y(y[88]));
  Fx110 Fx110_inst(.x({x[160], x[159], x[158], x[157], x[156]}), .y(y[89]));
  Fx111 Fx111_inst(.x({x[161], x[159]}), .y(y[90]));
  Fx112 Fx112_inst(.x({x[162], x[158]}), .y(y[91]));
  Fx113 Fx113_inst(.x({x[163], x[157]}), .y(y[92]));
  Fx114 Fx114_inst(.x({x[164], x[156]}), .y(y[93]));
  Fx115 Fx115_inst(.x({x[169], x[168], x[167], x[166], x[165]}), .y(y[94]));
  Fx116 Fx116_inst(.x({x[170], x[168]}), .y(y[95]));
  Fx117 Fx117_inst(.x({x[171], x[167]}), .y(y[96]));
  Fx118 Fx118_inst(.x({x[172], x[166]}), .y(y[97]));
  Fx119 Fx119_inst(.x({x[173], x[165]}), .y(y[98]));
  Fx120 Fx120_inst(.x({x[178], x[177], x[176], x[175], x[174]}), .y(y[99]));
  Fx121 Fx121_inst(.x({x[179], x[177]}), .y(y[100]));
  Fx122 Fx122_inst(.x({x[180], x[176]}), .y(y[101]));
  Fx123 Fx123_inst(.x({x[181], x[175]}), .y(y[102]));
  Fx124 Fx124_inst(.x({x[182], x[174]}), .y(y[103]));
  Fx125 Fx125_inst(.x({x[187], x[186], x[185], x[184], x[183]}), .y(y[104]));
  Fx126 Fx126_inst(.x({x[188], x[186]}), .y(y[105]));
  Fx127 Fx127_inst(.x({x[189], x[185]}), .y(y[106]));
  Fx128 Fx128_inst(.x({x[190], x[184]}), .y(y[107]));
  Fx129 Fx129_inst(.x({x[191], x[183]}), .y(y[108]));
  Fx130 Fx130_inst(.x({x[196], x[195], x[194], x[193], x[192]}), .y(y[109]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[110]));
  Fx132 Fx132_inst(.x({x[198], x[194]}), .y(y[111]));
  Fx133 Fx133_inst(.x({x[199], x[193]}), .y(y[112]));
  Fx134 Fx134_inst(.x({x[200], x[192]}), .y(y[113]));
  Fx135 Fx135_inst(.x({x[205], x[204], x[203], x[202], x[201]}), .y(y[114]));
  Fx136 Fx136_inst(.x({x[206], x[204]}), .y(y[115]));
  Fx137 Fx137_inst(.x({x[207], x[203]}), .y(y[116]));
  Fx138 Fx138_inst(.x({x[208], x[202]}), .y(y[117]));
  Fx139 Fx139_inst(.x({x[209], x[201]}), .y(y[118]));
  Fx140 Fx140_inst(.x({x[214], x[213], x[212], x[211], x[210]}), .y(y[119]));
  Fx141 Fx141_inst(.x({x[215], x[213]}), .y(y[120]));
  Fx142 Fx142_inst(.x({x[216], x[212]}), .y(y[121]));
  Fx143 Fx143_inst(.x({x[217], x[211]}), .y(y[122]));
  Fx144 Fx144_inst(.x({x[218], x[210]}), .y(y[123]));
  Fx145 Fx145_inst(.x({x[223], x[222], x[221], x[220], x[219]}), .y(y[124]));
  Fx146 Fx146_inst(.x({x[224], x[222]}), .y(y[125]));
  Fx147 Fx147_inst(.x({x[225], x[221]}), .y(y[126]));
  Fx148 Fx148_inst(.x({x[226], x[220]}), .y(y[127]));
  Fx149 Fx149_inst(.x({x[227], x[219]}), .y(y[128]));
  Fx150 Fx150_inst(.x({x[232], x[231], x[230], x[229], x[228]}), .y(y[129]));
  Fx151 Fx151_inst(.x({x[233], x[231]}), .y(y[130]));
  Fx152 Fx152_inst(.x({x[234], x[230]}), .y(y[131]));
  Fx153 Fx153_inst(.x({x[235], x[229]}), .y(y[132]));
  Fx154 Fx154_inst(.x({x[236], x[228]}), .y(y[133]));
  Fx155 Fx155_inst(.x({x[241], x[240], x[239], x[238], x[237]}), .y(y[134]));
  Fx156 Fx156_inst(.x({x[242], x[240]}), .y(y[135]));
  Fx157 Fx157_inst(.x({x[243], x[239]}), .y(y[136]));
  Fx158 Fx158_inst(.x({x[244], x[238]}), .y(y[137]));
  Fx159 Fx159_inst(.x({x[245], x[237]}), .y(y[138]));
  Fx160 Fx160_inst(.x({x[250], x[249], x[248], x[247], x[246]}), .y(y[139]));
  Fx161 Fx161_inst(.x({x[251], x[249]}), .y(y[140]));
  Fx162 Fx162_inst(.x({x[252], x[248]}), .y(y[141]));
  Fx163 Fx163_inst(.x({x[253], x[247]}), .y(y[142]));
  Fx164 Fx164_inst(.x({x[254], x[246]}), .y(y[143]));
  Fx165 Fx165_inst(.x({x[259], x[258], x[257], x[256], x[255]}), .y(y[144]));
  Fx166 Fx166_inst(.x({x[260], x[258]}), .y(y[145]));
  Fx167 Fx167_inst(.x({x[261], x[257]}), .y(y[146]));
  Fx168 Fx168_inst(.x({x[262], x[256]}), .y(y[147]));
  Fx169 Fx169_inst(.x({x[263], x[255]}), .y(y[148]));
  Fx170 Fx170_inst(.x({x[268], x[267], x[266], x[265], x[264]}), .y(y[149]));
  Fx171 Fx171_inst(.x({x[269], x[267]}), .y(y[150]));
  Fx172 Fx172_inst(.x({x[270], x[266]}), .y(y[151]));
  Fx173 Fx173_inst(.x({x[271], x[265]}), .y(y[152]));
  Fx174 Fx174_inst(.x({x[272], x[264]}), .y(y[153]));
  Fx175 Fx175_inst(.x({x[277], x[276], x[275], x[274], x[273]}), .y(y[154]));
  Fx176 Fx176_inst(.x({x[278], x[276]}), .y(y[155]));
  Fx177 Fx177_inst(.x({x[279], x[275]}), .y(y[156]));
  Fx178 Fx178_inst(.x({x[280], x[274]}), .y(y[157]));
  Fx179 Fx179_inst(.x({x[281], x[273]}), .y(y[158]));
  Fx180 Fx180_inst(.x({x[286], x[285], x[284], x[283], x[282]}), .y(y[159]));
  Fx181 Fx181_inst(.x({x[287], x[285]}), .y(y[160]));
  Fx182 Fx182_inst(.x({x[288], x[284]}), .y(y[161]));
  Fx183 Fx183_inst(.x({x[289], x[283]}), .y(y[162]));
  Fx184 Fx184_inst(.x({x[290], x[282]}), .y(y[163]));
  Fx185 Fx185_inst(.x({x[295], x[294], x[293], x[292], x[291]}), .y(y[164]));
  Fx186 Fx186_inst(.x({x[296], x[294]}), .y(y[165]));
  Fx187 Fx187_inst(.x({x[297], x[293]}), .y(y[166]));
  Fx188 Fx188_inst(.x({x[298], x[292]}), .y(y[167]));
  Fx189 Fx189_inst(.x({x[299], x[291]}), .y(y[168]));
  Fx190 Fx190_inst(.x({x[304], x[303], x[302], x[301], x[300]}), .y(y[169]));
  Fx191 Fx191_inst(.x({x[305], x[303]}), .y(y[170]));
  Fx192 Fx192_inst(.x({x[306], x[302]}), .y(y[171]));
  Fx193 Fx193_inst(.x({x[307], x[301]}), .y(y[172]));
  Fx194 Fx194_inst(.x({x[308], x[300]}), .y(y[173]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [17:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[16] ^ x[17];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[6] & x[7]);
  assign t[14] = (x[9] & x[10]);
  assign t[15] = (x[12] & x[13]);
  assign t[16] = (x[15] & x[16]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[2] = ~(t[7] | t[8]);
  assign t[3] = ~(t[9] | t[4]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[11] ^ x[2];
  assign t[6] = t[12] ^ x[5];
  assign t[7] = t[13] ^ x[8];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[14];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind66(x, y);
 input [18:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] ? t[6] : t[1];
  assign t[10] = t[16] ^ x[18];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[15] = (x[13] & x[14]);
  assign t[16] = (x[16] & x[17]);
  assign t[1] = ~(t[6] & t[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = t[7] & t[8];
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[3];
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[9];
  assign t[8] = t[14] ^ x[12];
  assign t[9] = t[15] ^ x[15];
  assign y = ~(~x[0] & ~t[0]);
endmodule

module R1ind67(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind68(x, y);
 input [18:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] & t[5];
  assign t[10] = t[16] ^ x[18];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[15] = (x[13] & x[14]);
  assign t[16] = (x[16] & x[17]);
  assign t[1] = ~(t[2] & t[6]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[3];
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[9];
  assign t[8] = t[14] ^ x[12];
  assign t[9] = t[15] ^ x[15];
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind71(x, y);
 input [18:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] | t[1];
  assign t[10] = t[16] ^ x[18];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[15] = (x[13] & x[14]);
  assign t[16] = (x[16] & x[17]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[4] = ~(t[9] & t[10]);
  assign t[5] = t[11] ^ x[3];
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[9];
  assign t[8] = t[14] ^ x[12];
  assign t[9] = t[15] ^ x[15];
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind73(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind74(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind75(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind76(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind77(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind78(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind79(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind80(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind81(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind82(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind83(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind84(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind85(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind86(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind87(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind88(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind89(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind90(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind91(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind92(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind93(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind94(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind95(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind96(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind97(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind98(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind99(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind100(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind101(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind102(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind103(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind104(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind105(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind106(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind107(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind108(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind109(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind110(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind111(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind112(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind113(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind114(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind115(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind116(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind117(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind118(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind119(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind120(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind121(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind122(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind123(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind124(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind125(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind126(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind127(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind128(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind129(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind130(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind131(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind132(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind133(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind134(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind135(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = x[0] ? x[4] : t[0];
endmodule

module R1ind136(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind137(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind138(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind139(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind140(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind141(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind142(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind143(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind144(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind145(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind146(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind147(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind148(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind149(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind150(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind151(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind152(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind153(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind154(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind155(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind156(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind157(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind158(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind159(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind160(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind161(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind162(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind163(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind164(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind165(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind166(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind167(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[3];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind168(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind169(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind170(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind171(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind172(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind173(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind174(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind175(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind176(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind177(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind178(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind179(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind180(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind181(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind182(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind183(x, y);
 input [2:0] x;
 output y;

  assign y = x[0] ? x[2] : x[1];
endmodule

module R1ind184(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind185(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind186(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind187(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind188(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind189(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind190(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind191(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind192(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind193(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind194(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind195(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind196(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind197(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind198(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind199(x, y);
 input [4:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = ~(x[2] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[4]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind200(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind201(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind202(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind203(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind204(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind205(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind206(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind207(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind208(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind209(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind210(x, y);
 input [8:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = t[20] ^ x[2];
  assign t[17] = t[21] ^ x[4];
  assign t[18] = t[22] ^ x[6];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (x[0] & x[1]);
  assign t[21] = (x[0] & x[3]);
  assign t[22] = (x[0] & x[5]);
  assign t[23] = (x[0] & x[7]);
  assign t[2] = t[5] ^ t[6];
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = ~(t[0]);
endmodule

module R1ind211(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind212(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind213(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind214(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind215(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind216(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind217(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind218(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind219(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind220(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind221(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind222(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind223(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind224(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind225(x, y);
 input [14:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[22]);
  assign t[12] = ~(t[21] ^ t[11]);
  assign t[13] = t[23] ^ t[22];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[21] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[21] ^ t[18];
  assign t[18] = t[22] ^ t[24];
  assign t[19] = t[25] ^ x[2];
  assign t[1] = ~(t[2] ^ t[20]);
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[6] & x[9]);
  assign t[29] = (x[6] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & x[13]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[21] & t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = ~(t[0] ^ t[19]);
endmodule

module R1ind226(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind227(x, y);
 input [14:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[22] ^ t[23];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[21] ^ t[12]);
  assign t[14] = t[21] & t[16];
  assign t[15] = t[21] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[23] ^ t[24];
  assign t[18] = t[21] ^ t[10];
  assign t[19] = t[25] ^ x[2];
  assign t[1] = ~(t[2] ^ t[20]);
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[6] & x[9]);
  assign t[29] = (x[6] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & x[13]);
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] ^ t[9];
  assign t[6] = t[10] ^ t[11];
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[21] ^ t[12];
  assign y = ~(t[0] ^ t[19]);
endmodule

module R1ind228(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind229(x, y);
 input [12:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[10];
  assign t[13] = t[18] ^ x[12];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[6] & x[9]);
  assign t[18] = (x[6] & x[11]);
  assign t[1] = ~(t[2] ^ t[10]);
  assign t[2] = ~t[3];
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[13] ^ t[7]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] ^ t[9]);
endmodule

module R1ind230(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind231(x, y);
 input [14:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[17] ^ t[9]);
  assign t[11] = t[17] ^ t[12];
  assign t[12] = t[16] ^ t[18];
  assign t[13] = t[19] ^ x[2];
  assign t[14] = t[20] ^ x[5];
  assign t[15] = t[21] ^ x[8];
  assign t[16] = t[22] ^ x[10];
  assign t[17] = t[23] ^ x[12];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = ~(t[2] ^ t[14]);
  assign t[20] = (x[3] & x[4]);
  assign t[21] = (x[6] & x[7]);
  assign t[22] = (x[6] & x[9]);
  assign t[23] = (x[6] & x[11]);
  assign t[24] = (x[6] & x[13]);
  assign t[2] = ~t[3];
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[15] ^ t[16];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[13]);
endmodule

module R1ind232(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind233(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind234(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind235(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind236(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind237(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind238(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind239(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind240(x, y);
 input [14:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[22]);
  assign t[12] = ~(t[21] ^ t[11]);
  assign t[13] = t[23] ^ t[22];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[21] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[21] ^ t[18];
  assign t[18] = t[22] ^ t[24];
  assign t[19] = t[25] ^ x[2];
  assign t[1] = ~(t[2] ^ t[20]);
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[6] & x[9]);
  assign t[29] = (x[6] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & x[13]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[21] & t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = ~(t[0] ^ t[19]);
endmodule

module R1ind241(x, y);
 input [14:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[22] ^ t[23];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[21] ^ t[12]);
  assign t[14] = t[21] & t[16];
  assign t[15] = t[21] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[23] ^ t[24];
  assign t[18] = t[21] ^ t[10];
  assign t[19] = t[25] ^ x[2];
  assign t[1] = ~(t[2] ^ t[20]);
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[6] & x[9]);
  assign t[29] = (x[6] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & x[13]);
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] ^ t[9];
  assign t[6] = t[10] ^ t[11];
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[21] ^ t[12];
  assign y = ~(t[0] ^ t[19]);
endmodule

module R1ind242(x, y);
 input [9:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[7];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[3] & x[6]);
  assign t[16] = (x[3] & x[8]);
  assign t[1] = ~t[2];
  assign t[2] = ~t[3];
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[10] ^ t[11];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[12] ^ t[7]);
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0] ^ t[9]);
endmodule

module R1ind243(x, y);
 input [11:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] ^ t[12];
  assign t[12] = t[15] ^ t[17];
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[7];
  assign t[16] = t[21] ^ x[9];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = (x[0] & x[1]);
  assign t[19] = (x[3] & x[4]);
  assign t[1] = ~t[2];
  assign t[20] = (x[3] & x[6]);
  assign t[21] = (x[3] & x[8]);
  assign t[22] = (x[3] & x[10]);
  assign t[2] = ~t[3];
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[14] ^ t[15];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[13]);
endmodule

module R1ind244(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind245(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind246(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind247(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind248(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind249(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind250(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind251(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind252(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind253(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind254(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind255(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind256(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[18] ^ t[9]);
  assign t[11] = t[20] ^ t[19];
  assign t[12] = ~(t[15] ^ t[6]);
  assign t[13] = t[18] ^ t[11];
  assign t[14] = t[9] & t[15];
  assign t[15] = t[18] ^ t[16];
  assign t[16] = t[19] ^ t[21];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = t[2] ^ t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] & t[7];
  assign t[4] = t[18] & t[8];
  assign t[5] = t[9] & t[10];
  assign t[6] = t[11] ^ t[9];
  assign t[7] = t[12] ^ t[5];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = ~(t[19]);
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind257(x, y);
 input [11:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] & t[14];
  assign t[13] = t[18] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[20] ^ t[21];
  assign t[16] = t[18] ^ t[8];
  assign t[17] = t[22] ^ x[2];
  assign t[18] = t[23] ^ x[5];
  assign t[19] = t[24] ^ x[7];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[11];
  assign t[22] = (x[0] & x[1]);
  assign t[23] = (x[3] & x[4]);
  assign t[24] = (x[3] & x[6]);
  assign t[25] = (x[3] & x[8]);
  assign t[26] = (x[3] & x[10]);
  assign t[2] = t[4] ^ t[5];
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[18] ^ t[10];
  assign t[8] = t[19] ^ t[20];
  assign t[9] = t[10] & t[13];
  assign y = ~(t[0] ^ t[17]);
endmodule

module R1ind258(x, y);
 input [9:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[14] ^ x[9];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[3] & x[6]);
  assign t[14] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[8] ^ t[9];
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[10] ^ t[5]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[7];
  assign y = ~(t[0] ^ t[7]);
endmodule

module R1ind259(x, y);
 input [11:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[13] ^ t[15];
  assign t[11] = t[16] ^ x[2];
  assign t[12] = t[17] ^ x[5];
  assign t[13] = t[18] ^ x[7];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[11];
  assign t[16] = (x[0] & x[1]);
  assign t[17] = (x[3] & x[4]);
  assign t[18] = (x[3] & x[6]);
  assign t[19] = (x[3] & x[8]);
  assign t[1] = ~(t[2]);
  assign t[20] = (x[3] & x[10]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[12] ^ t[13];
  assign t[6] = t[7] & t[9];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14] ^ t[7]);
  assign t[9] = t[14] ^ t[10];
  assign y = ~(t[0] ^ t[11]);
endmodule

module R1ind260(x, y);
 input [14:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[22]);
  assign t[12] = ~(t[21] ^ t[11]);
  assign t[13] = t[23] ^ t[22];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[21] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[21] ^ t[18];
  assign t[18] = t[22] ^ t[24];
  assign t[19] = t[25] ^ x[2];
  assign t[1] = ~(t[2] ^ t[20]);
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[6] & x[9]);
  assign t[29] = (x[6] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & x[13]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[21] & t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = ~(t[0] ^ t[19]);
endmodule

module R1ind261(x, y);
 input [14:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[22] ^ t[23];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[21] ^ t[12]);
  assign t[14] = t[21] & t[16];
  assign t[15] = t[21] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[23] ^ t[24];
  assign t[18] = t[21] ^ t[10];
  assign t[19] = t[25] ^ x[2];
  assign t[1] = ~(t[2] ^ t[20]);
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[12];
  assign t[24] = t[30] ^ x[14];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[6] & x[9]);
  assign t[29] = (x[6] & x[11]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & x[13]);
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] ^ t[9];
  assign t[6] = t[10] ^ t[11];
  assign t[7] = t[12] & t[13];
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[21] ^ t[12];
  assign y = ~(t[0] ^ t[19]);
endmodule

module R1ind262(x, y);
 input [12:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = ~t[1];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[10];
  assign t[13] = t[18] ^ x[12];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[6] & x[9]);
  assign t[18] = (x[6] & x[11]);
  assign t[1] = ~(t[2] ^ t[10]);
  assign t[2] = ~t[3];
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[11] ^ t[12];
  assign t[6] = t[7] & t[8];
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[13] ^ t[7]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] ^ t[9]);
endmodule

module R1ind263(x, y);
 input [14:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = ~t[1];
  assign t[10] = ~(t[17] ^ t[9]);
  assign t[11] = t[17] ^ t[12];
  assign t[12] = t[16] ^ t[18];
  assign t[13] = t[19] ^ x[2];
  assign t[14] = t[20] ^ x[5];
  assign t[15] = t[21] ^ x[8];
  assign t[16] = t[22] ^ x[10];
  assign t[17] = t[23] ^ x[12];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = ~(t[2] ^ t[14]);
  assign t[20] = (x[3] & x[4]);
  assign t[21] = (x[6] & x[7]);
  assign t[22] = (x[6] & x[9]);
  assign t[23] = (x[6] & x[11]);
  assign t[24] = (x[6] & x[13]);
  assign t[2] = ~t[3];
  assign t[3] = ~(t[4]);
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[15] ^ t[16];
  assign t[8] = t[9] & t[11];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[13]);
endmodule

module R1ind264(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind265(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind266(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind267(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind268(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind269(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind270(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind271(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind272(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind273(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind274(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind275(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1ind276(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = ~(t[13] ^ t[4]);
  assign t[11] = t[15] ^ t[9];
  assign t[12] = t[7] & t[13];
  assign t[13] = t[15] ^ t[14];
  assign t[14] = t[16] ^ t[18];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] & t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[15] & t[6];
  assign t[3] = t[7] & t[8];
  assign t[4] = t[9] ^ t[7];
  assign t[5] = t[10] ^ t[3];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[16]);
  assign t[8] = ~(t[15] ^ t[7]);
  assign t[9] = t[17] ^ t[16];
  assign y = t[0] ^ t[1];
endmodule

module R1ind277(x, y);
 input [8:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = t[2] ^ t[3];
  assign t[10] = t[15] & t[12];
  assign t[11] = t[15] ^ t[13];
  assign t[12] = t[14] ^ t[7];
  assign t[13] = t[17] ^ t[18];
  assign t[14] = t[15] ^ t[6];
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[4];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[8];
  assign t[19] = (x[0] & x[1]);
  assign t[1] = t[4] ^ t[5];
  assign t[20] = (x[0] & x[3]);
  assign t[21] = (x[0] & x[5]);
  assign t[22] = (x[0] & x[7]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[8] & t[9];
  assign t[4] = t[10] ^ t[3];
  assign t[5] = t[15] ^ t[8];
  assign t[6] = t[16] ^ t[17];
  assign t[7] = t[8] & t[11];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind278(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (x[0] & x[5]);
  assign t[1] = t[5] ^ t[6];
  assign t[2] = t[3] & t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[7] ^ t[3]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0]);
endmodule

module R1ind279(x, y);
 input [8:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[0] & x[3]);
  assign t[15] = (x[0] & x[5]);
  assign t[16] = (x[0] & x[7]);
  assign t[1] = t[3] ^ t[4];
  assign t[2] = t[5] & t[6];
  assign t[3] = t[9] ^ t[10];
  assign t[4] = t[5] & t[7];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11] ^ t[5]);
  assign t[7] = t[11] ^ t[8];
  assign t[8] = t[10] ^ t[12];
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0]);
endmodule

module R1_ind(x, y);
 input [517:0] x;
 output [279:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[164], x[163], x[162], x[152], x[151], x[150], x[149], x[148], x[147], x[165]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[164], x[163], x[162], x[165]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[161], x[160], x[159], x[158], x[157], x[156], x[164], x[163], x[162], x[149], x[148], x[147], x[152], x[151], x[150], x[155], x[154], x[153], x[165]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[158], x[157], x[156], x[165]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[161], x[160], x[159], x[165]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[155], x[154], x[153], x[164], x[163], x[162], x[158], x[157], x[156], x[152], x[151], x[150], x[161], x[160], x[159], x[149], x[148], x[147], x[165]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[169], x[168], x[167], x[166], x[165]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[172], x[171], x[170], x[166], x[165]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[175], x[174], x[173], x[166], x[165]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[178], x[177], x[176], x[166], x[165]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[182], x[181], x[180], x[179], x[165]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[185], x[184], x[183], x[179], x[165]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[188], x[187], x[186], x[179], x[165]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[191], x[190], x[189], x[179], x[165]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[195], x[194], x[193], x[192], x[165]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[198], x[197], x[196], x[192], x[165]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[201], x[200], x[199], x[192], x[165]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[204], x[203], x[202], x[192], x[165]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[208], x[207], x[206], x[205], x[165]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[211], x[210], x[209], x[205], x[165]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[214], x[213], x[212], x[205], x[165]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[217], x[216], x[215], x[205], x[165]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[221], x[220], x[219], x[218], x[165]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[224], x[223], x[222], x[218], x[165]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[227], x[226], x[225], x[218], x[165]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[230], x[229], x[228], x[218], x[165]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[234], x[233], x[232], x[231], x[165]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[237], x[236], x[235], x[231], x[165]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[240], x[239], x[238], x[231], x[165]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[243], x[242], x[241], x[231], x[165]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[247], x[246], x[245], x[244], x[165]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[250], x[249], x[248], x[244], x[165]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[253], x[252], x[251], x[244], x[165]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[256], x[255], x[254], x[244], x[165]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[260], x[259], x[258], x[257], x[165]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[263], x[262], x[261], x[257], x[165]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[266], x[265], x[264], x[257], x[165]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[269], x[268], x[267], x[257], x[165]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[273], x[272], x[271], x[270], x[165]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[276], x[275], x[274], x[270], x[165]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[279], x[278], x[277], x[270], x[165]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[282], x[281], x[280], x[270], x[165]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[286], x[285], x[284], x[283], x[165]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[289], x[288], x[287], x[283], x[165]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[292], x[291], x[290], x[283], x[165]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[295], x[294], x[293], x[283], x[165]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[299], x[298], x[297], x[296], x[165]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[302], x[301], x[300], x[296], x[165]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[305], x[304], x[303], x[296], x[165]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[308], x[307], x[306], x[296], x[165]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[312], x[311], x[310], x[309], x[165]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[315], x[314], x[313], x[309], x[165]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[318], x[317], x[316], x[309], x[165]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[321], x[320], x[319], x[309], x[165]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[325], x[324], x[323], x[322], x[165]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[328], x[327], x[326], x[322], x[165]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[331], x[330], x[329], x[322], x[165]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[334], x[333], x[332], x[322], x[165]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[338], x[337], x[336], x[335], x[165]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[341], x[340], x[339], x[335], x[165]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[344], x[343], x[342], x[335], x[165]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[347], x[346], x[345], x[335], x[165]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[351], x[350], x[349], x[348], x[165]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[354], x[353], x[352], x[348], x[165]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[357], x[356], x[355], x[348], x[165]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[360], x[359], x[358], x[348], x[165]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[364], x[363], x[362], x[361], x[165]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[367], x[366], x[365], x[361], x[165]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[370], x[369], x[368], x[361], x[165]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[373], x[372], x[371], x[361], x[165]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[376], x[375], x[374], x[165]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[379], x[378], x[377], x[165]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[382], x[381], x[380], x[165]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[385], x[384], x[383], x[165]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[388], x[387], x[386], x[165]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[391], x[390], x[389], x[165]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[394], x[393], x[392], x[165]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[397], x[396], x[395], x[165]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[400], x[399], x[398], x[165]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[403], x[402], x[401], x[165]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[406], x[405], x[404], x[165]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[409], x[408], x[407], x[165]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[412], x[411], x[410], x[165]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[415], x[414], x[413], x[165]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[418], x[417], x[416], x[165]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[421], x[420], x[419], x[165]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[423], x[375], x[422], x[165]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[425], x[378], x[424], x[165]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[427], x[381], x[426], x[165]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[429], x[384], x[428], x[165]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[431], x[387], x[430], x[165]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[433], x[390], x[432], x[165]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[435], x[393], x[434], x[165]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[437], x[396], x[436], x[165]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[439], x[399], x[438], x[165]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[441], x[402], x[440], x[165]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[443], x[405], x[442], x[165]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[445], x[408], x[444], x[165]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[447], x[411], x[446], x[165]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[449], x[414], x[448], x[165]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[451], x[417], x[450], x[165]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[453], x[420], x[452], x[165]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[455], x[454], x[165]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[457], x[456], x[165]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[459], x[458], x[165]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[461], x[460], x[165]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[463], x[462], x[165]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[465], x[464], x[165]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[467], x[466], x[165]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[469], x[468], x[165]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[471], x[470], x[165]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[473], x[472], x[165]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[475], x[474], x[165]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[477], x[476], x[165]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[479], x[478], x[165]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[481], x[480], x[165]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[483], x[482], x[165]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[485], x[484], x[165]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[487], x[375], x[376], x[486], x[165]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[489], x[378], x[379], x[488], x[165]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[491], x[381], x[382], x[490], x[165]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[493], x[384], x[385], x[492], x[165]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[495], x[387], x[388], x[494], x[165]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[497], x[390], x[391], x[496], x[165]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[499], x[393], x[394], x[498], x[165]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[501], x[396], x[397], x[500], x[165]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[503], x[399], x[400], x[502], x[165]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[505], x[402], x[403], x[504], x[165]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[507], x[405], x[406], x[506], x[165]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[509], x[408], x[409], x[508], x[165]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[511], x[411], x[412], x[510], x[165]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[513], x[414], x[415], x[512], x[165]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[515], x[417], x[418], x[514], x[165]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[517], x[420], x[421], x[516], x[165]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[65], x[64], x[59], x[58], x[63], x[62], x[61], x[60], x[57]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[119], x[118], x[113], x[112], x[117], x[116], x[115], x[114], x[111], x[220], x[219], x[218]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[65], x[64], x[63], x[62], x[59], x[58], x[61], x[60], x[57]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[119], x[118], x[117], x[116], x[113], x[112], x[115], x[114], x[111], x[223], x[222], x[218]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[61], x[60], x[65], x[64], x[63], x[62], x[57]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[115], x[114], x[119], x[118], x[117], x[116], x[111], x[226], x[225], x[218]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[65], x[64], x[61], x[60], x[63], x[62], x[59], x[58], x[57]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[119], x[118], x[115], x[114], x[117], x[116], x[113], x[112], x[111], x[229], x[228], x[218]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[74], x[73], x[68], x[67], x[72], x[71], x[70], x[69], x[66]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[128], x[127], x[122], x[121], x[126], x[125], x[124], x[123], x[120], x[233], x[232], x[231]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[74], x[73], x[72], x[71], x[68], x[67], x[70], x[69], x[66]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[128], x[127], x[126], x[125], x[122], x[121], x[124], x[123], x[120], x[236], x[235], x[231]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[70], x[69], x[74], x[73], x[72], x[71], x[66]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[124], x[123], x[128], x[127], x[126], x[125], x[120], x[239], x[238], x[231]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[74], x[73], x[70], x[69], x[72], x[71], x[68], x[67], x[66]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[128], x[127], x[124], x[123], x[126], x[125], x[122], x[121], x[120], x[242], x[241], x[231]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[47], x[46], x[41], x[40], x[45], x[44], x[43], x[42], x[39]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[137], x[136], x[131], x[130], x[135], x[134], x[133], x[132], x[129], x[246], x[245], x[244]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[47], x[46], x[45], x[44], x[41], x[40], x[43], x[42], x[39]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[137], x[136], x[135], x[134], x[131], x[130], x[133], x[132], x[129], x[249], x[248], x[244]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[43], x[42], x[47], x[46], x[45], x[44], x[39]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[133], x[132], x[137], x[136], x[135], x[134], x[129], x[252], x[251], x[244]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[47], x[46], x[43], x[42], x[45], x[44], x[41], x[40], x[39]}), .y(y[222]));
  R1ind223 R1ind223_inst(.x({x[137], x[136], x[133], x[132], x[135], x[134], x[131], x[130], x[129], x[255], x[254], x[244]}), .y(y[223]));
  R1ind224 R1ind224_inst(.x({x[56], x[55], x[50], x[49], x[54], x[53], x[52], x[51], x[48]}), .y(y[224]));
  R1ind225 R1ind225_inst(.x({x[146], x[145], x[140], x[139], x[144], x[143], x[142], x[141], x[138], x[164], x[163], x[162], x[259], x[258], x[257]}), .y(y[225]));
  R1ind226 R1ind226_inst(.x({x[56], x[55], x[54], x[53], x[50], x[49], x[52], x[51], x[48]}), .y(y[226]));
  R1ind227 R1ind227_inst(.x({x[146], x[145], x[144], x[143], x[140], x[139], x[142], x[141], x[138], x[155], x[154], x[153], x[262], x[261], x[257]}), .y(y[227]));
  R1ind228 R1ind228_inst(.x({x[52], x[51], x[56], x[55], x[54], x[53], x[48]}), .y(y[228]));
  R1ind229 R1ind229_inst(.x({x[142], x[141], x[146], x[145], x[144], x[143], x[138], x[158], x[157], x[156], x[265], x[264], x[257]}), .y(y[229]));
  R1ind230 R1ind230_inst(.x({x[56], x[55], x[52], x[51], x[54], x[53], x[50], x[49], x[48]}), .y(y[230]));
  R1ind231 R1ind231_inst(.x({x[146], x[145], x[142], x[141], x[144], x[143], x[140], x[139], x[138], x[161], x[160], x[159], x[268], x[267], x[257]}), .y(y[231]));
  R1ind232 R1ind232_inst(.x({x[92], x[91], x[86], x[85], x[90], x[89], x[88], x[87], x[84], x[181], x[180], x[179]}), .y(y[232]));
  R1ind233 R1ind233_inst(.x({x[92], x[91], x[90], x[89], x[86], x[85], x[88], x[87], x[84], x[184], x[183], x[179]}), .y(y[233]));
  R1ind234 R1ind234_inst(.x({x[88], x[87], x[92], x[91], x[90], x[89], x[84], x[187], x[186], x[179]}), .y(y[234]));
  R1ind235 R1ind235_inst(.x({x[92], x[91], x[88], x[87], x[90], x[89], x[86], x[85], x[84], x[190], x[189], x[179]}), .y(y[235]));
  R1ind236 R1ind236_inst(.x({x[101], x[100], x[95], x[94], x[99], x[98], x[97], x[96], x[93], x[194], x[193], x[192]}), .y(y[236]));
  R1ind237 R1ind237_inst(.x({x[101], x[100], x[99], x[98], x[95], x[94], x[97], x[96], x[93], x[197], x[196], x[192]}), .y(y[237]));
  R1ind238 R1ind238_inst(.x({x[97], x[96], x[101], x[100], x[99], x[98], x[93], x[200], x[199], x[192]}), .y(y[238]));
  R1ind239 R1ind239_inst(.x({x[101], x[100], x[97], x[96], x[99], x[98], x[95], x[94], x[93], x[203], x[202], x[192]}), .y(y[239]));
  R1ind240 R1ind240_inst(.x({x[110], x[109], x[104], x[103], x[108], x[107], x[106], x[105], x[102], x[149], x[148], x[147], x[207], x[206], x[205]}), .y(y[240]));
  R1ind241 R1ind241_inst(.x({x[110], x[109], x[108], x[107], x[104], x[103], x[106], x[105], x[102], x[152], x[151], x[150], x[210], x[209], x[205]}), .y(y[241]));
  R1ind242 R1ind242_inst(.x({x[106], x[105], x[110], x[109], x[108], x[107], x[102], x[213], x[212], x[205]}), .y(y[242]));
  R1ind243 R1ind243_inst(.x({x[110], x[109], x[106], x[105], x[108], x[107], x[104], x[103], x[102], x[216], x[215], x[205]}), .y(y[243]));
  R1ind244 R1ind244_inst(.x({x[83], x[82], x[77], x[76], x[81], x[80], x[79], x[78], x[75], x[168], x[167], x[166]}), .y(y[244]));
  R1ind245 R1ind245_inst(.x({x[83], x[82], x[81], x[80], x[77], x[76], x[79], x[78], x[75], x[171], x[170], x[166]}), .y(y[245]));
  R1ind246 R1ind246_inst(.x({x[79], x[78], x[83], x[82], x[81], x[80], x[75], x[174], x[173], x[166]}), .y(y[246]));
  R1ind247 R1ind247_inst(.x({x[83], x[82], x[79], x[78], x[81], x[80], x[77], x[76], x[75], x[177], x[176], x[166]}), .y(y[247]));
  R1ind248 R1ind248_inst(.x({x[119], x[118], x[113], x[112], x[117], x[116], x[115], x[114], x[111], x[220], x[219], x[218]}), .y(y[248]));
  R1ind249 R1ind249_inst(.x({x[119], x[118], x[117], x[116], x[113], x[112], x[115], x[114], x[111], x[223], x[222], x[218]}), .y(y[249]));
  R1ind250 R1ind250_inst(.x({x[115], x[114], x[119], x[118], x[117], x[116], x[111], x[226], x[225], x[218]}), .y(y[250]));
  R1ind251 R1ind251_inst(.x({x[119], x[118], x[115], x[114], x[117], x[116], x[113], x[112], x[111], x[229], x[228], x[218]}), .y(y[251]));
  R1ind252 R1ind252_inst(.x({x[128], x[127], x[122], x[121], x[126], x[125], x[124], x[123], x[120], x[233], x[232], x[231]}), .y(y[252]));
  R1ind253 R1ind253_inst(.x({x[128], x[127], x[126], x[125], x[122], x[121], x[124], x[123], x[120], x[236], x[235], x[231]}), .y(y[253]));
  R1ind254 R1ind254_inst(.x({x[124], x[123], x[128], x[127], x[126], x[125], x[120], x[239], x[238], x[231]}), .y(y[254]));
  R1ind255 R1ind255_inst(.x({x[128], x[127], x[124], x[123], x[126], x[125], x[122], x[121], x[120], x[242], x[241], x[231]}), .y(y[255]));
  R1ind256 R1ind256_inst(.x({x[137], x[136], x[131], x[130], x[135], x[134], x[133], x[132], x[129], x[246], x[245], x[244]}), .y(y[256]));
  R1ind257 R1ind257_inst(.x({x[137], x[136], x[135], x[134], x[131], x[130], x[133], x[132], x[129], x[249], x[248], x[244]}), .y(y[257]));
  R1ind258 R1ind258_inst(.x({x[133], x[132], x[137], x[136], x[135], x[134], x[129], x[252], x[251], x[244]}), .y(y[258]));
  R1ind259 R1ind259_inst(.x({x[137], x[136], x[133], x[132], x[135], x[134], x[131], x[130], x[129], x[255], x[254], x[244]}), .y(y[259]));
  R1ind260 R1ind260_inst(.x({x[146], x[145], x[140], x[139], x[144], x[143], x[142], x[141], x[138], x[164], x[163], x[162], x[259], x[258], x[257]}), .y(y[260]));
  R1ind261 R1ind261_inst(.x({x[146], x[145], x[144], x[143], x[140], x[139], x[142], x[141], x[138], x[155], x[154], x[153], x[262], x[261], x[257]}), .y(y[261]));
  R1ind262 R1ind262_inst(.x({x[142], x[141], x[146], x[145], x[144], x[143], x[138], x[158], x[157], x[156], x[265], x[264], x[257]}), .y(y[262]));
  R1ind263 R1ind263_inst(.x({x[146], x[145], x[142], x[141], x[144], x[143], x[140], x[139], x[138], x[161], x[160], x[159], x[268], x[267], x[257]}), .y(y[263]));
  R1ind264 R1ind264_inst(.x({x[38], x[37], x[32], x[31], x[36], x[35], x[34], x[33], x[30]}), .y(y[264]));
  R1ind265 R1ind265_inst(.x({x[38], x[37], x[36], x[35], x[32], x[31], x[34], x[33], x[30]}), .y(y[265]));
  R1ind266 R1ind266_inst(.x({x[34], x[33], x[38], x[37], x[36], x[35], x[30]}), .y(y[266]));
  R1ind267 R1ind267_inst(.x({x[38], x[37], x[34], x[33], x[36], x[35], x[32], x[31], x[30]}), .y(y[267]));
  R1ind268 R1ind268_inst(.x({x[11], x[10], x[5], x[4], x[9], x[8], x[7], x[6], x[3]}), .y(y[268]));
  R1ind269 R1ind269_inst(.x({x[11], x[10], x[9], x[8], x[5], x[4], x[7], x[6], x[3]}), .y(y[269]));
  R1ind270 R1ind270_inst(.x({x[7], x[6], x[11], x[10], x[9], x[8], x[3]}), .y(y[270]));
  R1ind271 R1ind271_inst(.x({x[11], x[10], x[7], x[6], x[9], x[8], x[5], x[4], x[3]}), .y(y[271]));
  R1ind272 R1ind272_inst(.x({x[20], x[19], x[14], x[13], x[18], x[17], x[16], x[15], x[12]}), .y(y[272]));
  R1ind273 R1ind273_inst(.x({x[20], x[19], x[18], x[17], x[14], x[13], x[16], x[15], x[12]}), .y(y[273]));
  R1ind274 R1ind274_inst(.x({x[16], x[15], x[20], x[19], x[18], x[17], x[12]}), .y(y[274]));
  R1ind275 R1ind275_inst(.x({x[20], x[19], x[16], x[15], x[18], x[17], x[14], x[13], x[12]}), .y(y[275]));
  R1ind276 R1ind276_inst(.x({x[29], x[28], x[23], x[22], x[27], x[26], x[25], x[24], x[21]}), .y(y[276]));
  R1ind277 R1ind277_inst(.x({x[29], x[28], x[27], x[26], x[23], x[22], x[25], x[24], x[21]}), .y(y[277]));
  R1ind278 R1ind278_inst(.x({x[25], x[24], x[29], x[28], x[27], x[26], x[21]}), .y(y[278]));
  R1ind279 R1ind279_inst(.x({x[29], x[28], x[25], x[24], x[27], x[26], x[23], x[22], x[21]}), .y(y[279]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[2];
  assign t[13] = t[19] ^ x[5];
  assign t[14] = t[20] ^ x[8];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[14];
  assign t[17] = t[23] ^ x[17];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[1];
  assign t[25] = t[37] ^ x[2];
  assign t[26] = t[38] ^ x[4];
  assign t[27] = t[39] ^ x[5];
  assign t[28] = t[40] ^ x[7];
  assign t[29] = t[41] ^ x[8];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[0]);
  assign t[38] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[6]);
  assign t[42] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[9]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[5] = ~(t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[2];
  assign t[13] = t[19] ^ x[5];
  assign t[14] = t[20] ^ x[8];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[14];
  assign t[17] = t[23] ^ x[17];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[1];
  assign t[25] = t[37] ^ x[2];
  assign t[26] = t[38] ^ x[4];
  assign t[27] = t[39] ^ x[5];
  assign t[28] = t[40] ^ x[7];
  assign t[29] = t[41] ^ x[8];
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[42] ^ x[10];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[13];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[0]);
  assign t[38] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[6]);
  assign t[42] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[9]);
  assign t[44] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[12]);
  assign t[46] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[15]);
  assign t[4] = ~(t[10] | t[5]);
  assign t[5] = ~(t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = t[8] & t[9];
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = t[8] & t[9];
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[2] & t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] & t[5]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind31(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind34(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[3];
  assign t[6] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind36(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind37(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind38(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind39(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[3];
  assign t[13] = t[19] ^ x[6];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[12];
  assign t[16] = t[22] ^ x[15];
  assign t[17] = t[23] ^ x[18];
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[6] | t[2];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[32] & t[33]);
  assign t[23] = (~t[34] & t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[3];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[6];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[9];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[12];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[1]);
  assign t[38] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[39] = (x[4]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[41] = (x[7]);
  assign t[42] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = (x[10]);
  assign t[44] = (x[13] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0 & ~1'b0) | (x[13] & 1'b0 & ~1'b0 & 1'b0) | (x[13] & ~1'b0 & 1'b0 & 1'b0) | (~x[13] & 1'b0 & 1'b0 & 1'b0);
  assign t[45] = (x[13]);
  assign t[46] = (x[16] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0 & ~1'b0) | (x[16] & 1'b0 & ~1'b0 & 1'b0) | (x[16] & ~1'b0 & 1'b0 & 1'b0) | (~x[16] & 1'b0 & 1'b0 & 1'b0);
  assign t[47] = (x[16]);
  assign t[4] = ~(t[9] | t[5]);
  assign t[5] = ~(t[10] & t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind41(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind42(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind43(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind44(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind45(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind46(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind47(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind48(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind49(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind50(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind51(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind52(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind53(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind54(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind55(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind56(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind57(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind58(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind59(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[2]);
  assign t[1] = ~x[0];
  assign t[2] = x[3] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind60(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind61(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind62(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind63(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind64(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind65(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind66(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind67(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind68(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind69(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind70(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind71(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind72(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind73(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind74(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind75(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind76(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind77(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind78(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind79(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(t[1] ^ x[1]);
  assign t[1] = ~x[2];
  assign t[2] = x[3] ? x[0] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind80(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind81(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind82(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind83(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind84(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind85(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind86(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind87(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind88(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind89(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind90(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind91(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind92(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind93(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind94(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind95(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind96(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind97(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind98(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind99(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = x[2] ? x[1] : x[0];
  assign y = t ^ 1'b0 ^ 1'b0;
endmodule

module R2ind100(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind101(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind102(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind103(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind104(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind105(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind106(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind107(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind108(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind109(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind110(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind111(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind112(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind113(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind114(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[2] ^ x[3]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind115(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind116(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind117(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind118(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind119(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~(x[0] ^ t[1]);
  assign t[1] = ~(x[3] ^ x[2]);
  assign t[2] = x[4] ? x[1] : t[0];
  assign y = t[2] ^ 1'b0 ^ 1'b0;
endmodule

module R2ind120(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind121(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind126(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind131(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind136(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind141(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind146(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind151(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind156(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind161(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind166(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind171(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind176(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind181(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind186(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind191(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [13:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = x[0] ? x[7] : t[4];
  assign t[10] = t[14] ^ x[10];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (~t[16] & t[17]);
  assign t[13] = (~t[16] & t[18]);
  assign t[14] = (~t[16] & t[19]);
  assign t[15] = (~t[16] & t[20]);
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[10];
  assign t[1] = x[0] ? x[9] : t[5];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[22] = (x[1]);
  assign t[23] = (x[2]);
  assign t[24] = (x[3]);
  assign t[25] = (x[4]);
  assign t[2] = x[0] ? x[11] : t[6];
  assign t[3] = x[0] ? x[13] : t[7];
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind196(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[4]);
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [7:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = x[0] ? x[7] : t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[6];
  assign t[3] = (~t[4] & t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[6];
  assign t[6] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind201(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind206(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [8:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[27] ^ t[26];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[25] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[25] ^ t[15];
  assign t[15] = t[26] ^ t[28];
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[18] ^ t[19]);
  assign t[18] = t[20] ^ t[4];
  assign t[19] = t[1] ^ t[21];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[10] ^ t[13];
  assign t[21] = t[25] ^ t[8];
  assign t[22] = ~(t[23]);
  assign t[23] = t[15] ^ t[4];
  assign t[24] = ~(t[18]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = t[33] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[6];
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = (~t[37] & t[38]);
  assign t[34] = (~t[37] & t[39]);
  assign t[35] = (~t[37] & t[40]);
  assign t[36] = (~t[37] & t[41]);
  assign t[37] = t[42] ^ x[4];
  assign t[38] = t[43] ^ x[5];
  assign t[39] = t[44] ^ x[6];
  assign t[3] = t[25] & t[7];
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[43] = (x[1]);
  assign t[44] = (x[2]);
  assign t[45] = (x[0]);
  assign t[46] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[26]);
  assign t[9] = ~(t[25] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[22] & ~t[24]) | (~t[0] & t[16] & ~t[22] & ~t[24]) | (~t[0] & ~t[16] & t[22] & ~t[24]) | (~t[0] & ~t[16] & ~t[22] & t[24]) | (t[0] & t[16] & t[22] & ~t[24]) | (t[0] & t[16] & ~t[22] & t[24]) | (t[0] & ~t[16] & t[22] & t[24]) | (~t[0] & t[16] & t[22] & t[24]);
endmodule

module R2ind211(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [8:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = ~(t[19]);
  assign t[11] = ~(t[17] ^ t[10]);
  assign t[12] = t[17] & t[14];
  assign t[13] = t[17] ^ t[15];
  assign t[14] = t[16] ^ t[9];
  assign t[15] = t[19] ^ t[20];
  assign t[16] = t[17] ^ t[8];
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = (t[24]);
  assign t[21] = t[25] ^ x[5];
  assign t[22] = t[26] ^ x[6];
  assign t[23] = t[27] ^ x[7];
  assign t[24] = t[28] ^ x[8];
  assign t[25] = (~t[29] & t[30]);
  assign t[26] = (~t[29] & t[31]);
  assign t[27] = (~t[29] & t[32]);
  assign t[28] = (~t[29] & t[33]);
  assign t[29] = t[34] ^ x[4];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[35] ^ x[5];
  assign t[31] = t[36] ^ x[6];
  assign t[32] = t[37] ^ x[7];
  assign t[33] = t[38] ^ x[8];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[1]);
  assign t[36] = (x[0]);
  assign t[37] = (x[2]);
  assign t[38] = (x[3]);
  assign t[3] = t[6] ^ t[7];
  assign t[4] = t[8] ^ t[9];
  assign t[5] = t[10] & t[11];
  assign t[6] = t[12] ^ t[5];
  assign t[7] = t[17] ^ t[10];
  assign t[8] = t[18] ^ t[19];
  assign t[9] = t[10] & t[13];
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind216(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind221(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind226(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind231(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [29:0] x;
 output y;

 wire [111:0] t;
  assign t[0] = ~(t[1] ^ t[40]);
  assign t[100] = (x[11]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[1]);
  assign t[104] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[105] = (x[19]);
  assign t[106] = (x[2]);
  assign t[107] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[23]);
  assign t[109] = (x[3]);
  assign t[10] = t[15] ^ t[8];
  assign t[110] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[111] = (x[27]);
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[43]);
  assign t[13] = ~(t[42] ^ t[12]);
  assign t[14] = t[44] ^ t[43];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[42] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[42] ^ t[19];
  assign t[19] = t[43] ^ t[45];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[46]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[47]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27] ^ t[8];
  assign t[26] = t[5] ^ t[28];
  assign t[27] = t[14] ^ t[17];
  assign t[28] = t[42] ^ t[12];
  assign t[29] = ~(t[30] ^ t[48]);
  assign t[2] = ~(t[3] ^ t[41]);
  assign t[30] = ~t[31];
  assign t[31] = ~(t[32] ^ t[49]);
  assign t[32] = ~t[33];
  assign t[33] = ~(t[34]);
  assign t[34] = t[19] ^ t[8];
  assign t[35] = ~(t[36] ^ t[50]);
  assign t[36] = ~t[37];
  assign t[37] = ~(t[38] ^ t[51]);
  assign t[38] = ~t[39];
  assign t[39] = ~(t[25]);
  assign t[3] = ~t[4];
  assign t[40] = (t[52]);
  assign t[41] = (t[53]);
  assign t[42] = (t[54]);
  assign t[43] = (t[55]);
  assign t[44] = (t[56]);
  assign t[45] = (t[57]);
  assign t[46] = (t[58]);
  assign t[47] = (t[59]);
  assign t[48] = (t[60]);
  assign t[49] = (t[61]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (t[62]);
  assign t[51] = (t[63]);
  assign t[52] = t[64] ^ x[5];
  assign t[53] = t[65] ^ x[8];
  assign t[54] = t[66] ^ x[14];
  assign t[55] = t[67] ^ x[15];
  assign t[56] = t[68] ^ x[16];
  assign t[57] = t[69] ^ x[17];
  assign t[58] = t[70] ^ x[18];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[25];
  assign t[62] = t[74] ^ x[26];
  assign t[63] = t[75] ^ x[29];
  assign t[64] = (~t[76] & t[77]);
  assign t[65] = (~t[78] & t[79]);
  assign t[66] = (~t[80] & t[81]);
  assign t[67] = (~t[80] & t[82]);
  assign t[68] = (~t[80] & t[83]);
  assign t[69] = (~t[80] & t[84]);
  assign t[6] = t[9] & t[10];
  assign t[70] = (~t[76] & t[85]);
  assign t[71] = (~t[86] & t[87]);
  assign t[72] = (~t[76] & t[88]);
  assign t[73] = (~t[89] & t[90]);
  assign t[74] = (~t[76] & t[91]);
  assign t[75] = (~t[92] & t[93]);
  assign t[76] = t[94] ^ x[4];
  assign t[77] = t[95] ^ x[5];
  assign t[78] = t[96] ^ x[7];
  assign t[79] = t[97] ^ x[8];
  assign t[7] = t[42] & t[11];
  assign t[80] = t[98] ^ x[13];
  assign t[81] = t[99] ^ x[14];
  assign t[82] = t[100] ^ x[15];
  assign t[83] = t[101] ^ x[16];
  assign t[84] = t[102] ^ x[17];
  assign t[85] = t[103] ^ x[18];
  assign t[86] = t[104] ^ x[20];
  assign t[87] = t[105] ^ x[21];
  assign t[88] = t[106] ^ x[22];
  assign t[89] = t[107] ^ x[24];
  assign t[8] = t[12] & t[13];
  assign t[90] = t[108] ^ x[25];
  assign t[91] = t[109] ^ x[26];
  assign t[92] = t[110] ^ x[28];
  assign t[93] = t[111] ^ x[29];
  assign t[94] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[95] = (x[0]);
  assign t[96] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[6]);
  assign t[98] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[99] = (x[10]);
  assign t[9] = t[14] ^ t[12];
  assign y = (t[0] & ~t[20] & ~t[29] & ~t[35]) | (~t[0] & t[20] & ~t[29] & ~t[35]) | (~t[0] & ~t[20] & t[29] & ~t[35]) | (~t[0] & ~t[20] & ~t[29] & t[35]) | (t[0] & t[20] & t[29] & ~t[35]) | (t[0] & t[20] & ~t[29] & t[35]) | (t[0] & ~t[20] & t[29] & t[35]) | (~t[0] & t[20] & t[29] & t[35]);
endmodule

module R2ind236(x, y);
 input [17:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[14]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] ^ t[13];
  assign t[13] = t[17] ^ t[19];
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[14];
  assign t[23] = t[29] ^ x[15];
  assign t[24] = t[30] ^ x[16];
  assign t[25] = t[31] ^ x[17];
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[34] & t[35]);
  assign t[28] = (~t[36] & t[37]);
  assign t[29] = (~t[36] & t[38]);
  assign t[2] = ~(t[3] ^ t[15]);
  assign t[30] = (~t[36] & t[39]);
  assign t[31] = (~t[36] & t[40]);
  assign t[32] = t[41] ^ x[4];
  assign t[33] = t[42] ^ x[5];
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[8];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[14];
  assign t[38] = t[47] ^ x[15];
  assign t[39] = t[48] ^ x[16];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[17];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[3]);
  assign t[43] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[44] = (x[6]);
  assign t[45] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[46] = (x[9]);
  assign t[47] = (x[11]);
  assign t[48] = (x[10]);
  assign t[49] = (x[12]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[16] ^ t[17];
  assign t[9] = t[10] & t[12];
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[10]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = t[24] ^ x[16];
  assign t[1] = ~t[2];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[29] & t[31]);
  assign t[24] = (~t[29] & t[32]);
  assign t[25] = t[33] ^ x[4];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[7];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[13];
  assign t[2] = ~(t[3] ^ t[11]);
  assign t[30] = t[38] ^ x[14];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[16];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[2]);
  assign t[35] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[6]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[12]);
  assign t[3] = ~t[4];
  assign t[40] = (x[10]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[12] ^ t[13];
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[14] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [17:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[22] ^ t[13];
  assign t[11] = t[23] ^ t[24];
  assign t[12] = t[13] & t[16];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[22] ^ t[13]);
  assign t[15] = t[22] & t[17];
  assign t[16] = t[22] ^ t[18];
  assign t[17] = t[19] ^ t[12];
  assign t[18] = t[24] ^ t[25];
  assign t[19] = t[22] ^ t[11];
  assign t[1] = ~t[2];
  assign t[20] = (t[26]);
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[8];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = t[36] ^ x[16];
  assign t[31] = t[37] ^ x[17];
  assign t[32] = (~t[38] & t[39]);
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[42] & t[46]);
  assign t[38] = t[47] ^ x[4];
  assign t[39] = t[48] ^ x[5];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[8];
  assign t[42] = t[51] ^ x[13];
  assign t[43] = t[52] ^ x[14];
  assign t[44] = t[53] ^ x[15];
  assign t[45] = t[54] ^ x[16];
  assign t[46] = t[55] ^ x[17];
  assign t[47] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[48] = (x[1]);
  assign t[49] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[5] ^ t[6]);
  assign t[50] = (x[6]);
  assign t[51] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[52] = (x[10]);
  assign t[53] = (x[9]);
  assign t[54] = (x[11]);
  assign t[55] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[8];
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [17:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[22] ^ t[12]);
  assign t[14] = t[24] ^ t[23];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[22] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[22] ^ t[19];
  assign t[19] = t[23] ^ t[25];
  assign t[1] = ~t[2];
  assign t[20] = (t[26]);
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[8];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = t[36] ^ x[16];
  assign t[31] = t[37] ^ x[17];
  assign t[32] = (~t[38] & t[39]);
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[42] & t[46]);
  assign t[38] = t[47] ^ x[4];
  assign t[39] = t[48] ^ x[5];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[8];
  assign t[42] = t[51] ^ x[13];
  assign t[43] = t[52] ^ x[14];
  assign t[44] = t[53] ^ x[15];
  assign t[45] = t[54] ^ x[16];
  assign t[46] = t[55] ^ x[17];
  assign t[47] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[48] = (x[0]);
  assign t[49] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[6]);
  assign t[51] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[52] = (x[10]);
  assign t[53] = (x[11]);
  assign t[54] = (x[9]);
  assign t[55] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[22] & t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = t[14] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind241(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind246(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [23:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[40]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[43]);
  assign t[13] = ~(t[42] ^ t[12]);
  assign t[14] = t[44] ^ t[43];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[42] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[42] ^ t[19];
  assign t[19] = t[43] ^ t[45];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[46]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[47]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27] ^ t[8];
  assign t[26] = t[5] ^ t[28];
  assign t[27] = t[14] ^ t[17];
  assign t[28] = t[42] ^ t[12];
  assign t[29] = ~(t[30] ^ t[48]);
  assign t[2] = ~(t[3] ^ t[41]);
  assign t[30] = ~t[31];
  assign t[31] = ~t[32];
  assign t[32] = ~t[33];
  assign t[33] = ~(t[34]);
  assign t[34] = t[19] ^ t[8];
  assign t[35] = ~(t[36] ^ t[49]);
  assign t[36] = ~t[37];
  assign t[37] = ~t[38];
  assign t[38] = ~t[39];
  assign t[39] = ~(t[25]);
  assign t[3] = ~t[4];
  assign t[40] = (t[50]);
  assign t[41] = (t[51]);
  assign t[42] = (t[52]);
  assign t[43] = (t[53]);
  assign t[44] = (t[54]);
  assign t[45] = (t[55]);
  assign t[46] = (t[56]);
  assign t[47] = (t[57]);
  assign t[48] = (t[58]);
  assign t[49] = (t[59]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = t[60] ^ x[5];
  assign t[51] = t[61] ^ x[8];
  assign t[52] = t[62] ^ x[14];
  assign t[53] = t[63] ^ x[15];
  assign t[54] = t[64] ^ x[16];
  assign t[55] = t[65] ^ x[17];
  assign t[56] = t[66] ^ x[18];
  assign t[57] = t[67] ^ x[21];
  assign t[58] = t[68] ^ x[22];
  assign t[59] = t[69] ^ x[23];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = (~t[70] & t[71]);
  assign t[61] = (~t[72] & t[73]);
  assign t[62] = (~t[74] & t[75]);
  assign t[63] = (~t[74] & t[76]);
  assign t[64] = (~t[74] & t[77]);
  assign t[65] = (~t[74] & t[78]);
  assign t[66] = (~t[70] & t[79]);
  assign t[67] = (~t[80] & t[81]);
  assign t[68] = (~t[70] & t[82]);
  assign t[69] = (~t[70] & t[83]);
  assign t[6] = t[9] & t[10];
  assign t[70] = t[84] ^ x[4];
  assign t[71] = t[85] ^ x[5];
  assign t[72] = t[86] ^ x[7];
  assign t[73] = t[87] ^ x[8];
  assign t[74] = t[88] ^ x[13];
  assign t[75] = t[89] ^ x[14];
  assign t[76] = t[90] ^ x[15];
  assign t[77] = t[91] ^ x[16];
  assign t[78] = t[92] ^ x[17];
  assign t[79] = t[93] ^ x[18];
  assign t[7] = t[42] & t[11];
  assign t[80] = t[94] ^ x[20];
  assign t[81] = t[95] ^ x[21];
  assign t[82] = t[96] ^ x[22];
  assign t[83] = t[97] ^ x[23];
  assign t[84] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[85] = (x[0]);
  assign t[86] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[6]);
  assign t[88] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[89] = (x[10]);
  assign t[8] = t[12] & t[13];
  assign t[90] = (x[11]);
  assign t[91] = (x[9]);
  assign t[92] = (x[12]);
  assign t[93] = (x[1]);
  assign t[94] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[19]);
  assign t[96] = (x[2]);
  assign t[97] = (x[3]);
  assign t[9] = t[14] ^ t[12];
  assign y = (t[0] & ~t[20] & ~t[29] & ~t[35]) | (~t[0] & t[20] & ~t[29] & ~t[35]) | (~t[0] & ~t[20] & t[29] & ~t[35]) | (~t[0] & ~t[20] & ~t[29] & t[35]) | (t[0] & t[20] & t[29] & ~t[35]) | (t[0] & t[20] & ~t[29] & t[35]) | (t[0] & ~t[20] & t[29] & t[35]) | (~t[0] & t[20] & t[29] & t[35]);
endmodule

module R2ind251(x, y);
 input [14:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[14]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17] ^ t[10]);
  assign t[12] = t[17] ^ t[13];
  assign t[13] = t[16] ^ t[18];
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[5];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[11];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[13];
  assign t[23] = t[28] ^ x[14];
  assign t[24] = (~t[29] & t[30]);
  assign t[25] = (~t[31] & t[32]);
  assign t[26] = (~t[31] & t[33]);
  assign t[27] = (~t[31] & t[34]);
  assign t[28] = (~t[31] & t[35]);
  assign t[29] = t[36] ^ x[4];
  assign t[2] = ~t[3];
  assign t[30] = t[37] ^ x[5];
  assign t[31] = t[38] ^ x[10];
  assign t[32] = t[39] ^ x[11];
  assign t[33] = t[40] ^ x[12];
  assign t[34] = t[41] ^ x[13];
  assign t[35] = t[42] ^ x[14];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[39] = (x[6]);
  assign t[3] = ~t[4];
  assign t[40] = (x[8]);
  assign t[41] = (x[7]);
  assign t[42] = (x[9]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[10] & t[12];
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [13:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = ~(t[1] ^ t[10]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[11];
  assign t[16] = t[20] ^ x[12];
  assign t[17] = t[21] ^ x[13];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = (~t[24] & t[26]);
  assign t[21] = (~t[24] & t[27]);
  assign t[22] = t[28] ^ x[4];
  assign t[23] = t[29] ^ x[5];
  assign t[24] = t[30] ^ x[10];
  assign t[25] = t[31] ^ x[11];
  assign t[26] = t[32] ^ x[12];
  assign t[27] = t[33] ^ x[13];
  assign t[28] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[29] = (x[2]);
  assign t[2] = ~t[3];
  assign t[30] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[31] = (x[8]);
  assign t[32] = (x[9]);
  assign t[33] = (x[7]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[11] ^ t[12];
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[13] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [17:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[22] ^ t[13];
  assign t[11] = t[23] ^ t[24];
  assign t[12] = t[13] & t[16];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[22] ^ t[13]);
  assign t[15] = t[22] & t[17];
  assign t[16] = t[22] ^ t[18];
  assign t[17] = t[19] ^ t[12];
  assign t[18] = t[24] ^ t[25];
  assign t[19] = t[22] ^ t[11];
  assign t[1] = ~t[2];
  assign t[20] = (t[26]);
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[8];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = t[36] ^ x[16];
  assign t[31] = t[37] ^ x[17];
  assign t[32] = (~t[38] & t[39]);
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[42] & t[46]);
  assign t[38] = t[47] ^ x[4];
  assign t[39] = t[48] ^ x[5];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[8];
  assign t[42] = t[51] ^ x[13];
  assign t[43] = t[52] ^ x[14];
  assign t[44] = t[53] ^ x[15];
  assign t[45] = t[54] ^ x[16];
  assign t[46] = t[55] ^ x[17];
  assign t[47] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[48] = (x[1]);
  assign t[49] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[5] ^ t[6]);
  assign t[50] = (x[6]);
  assign t[51] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[52] = (x[10]);
  assign t[53] = (x[9]);
  assign t[54] = (x[11]);
  assign t[55] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[8];
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [17:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[22] ^ t[12]);
  assign t[14] = t[24] ^ t[23];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[22] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[22] ^ t[19];
  assign t[19] = t[23] ^ t[25];
  assign t[1] = ~t[2];
  assign t[20] = (t[26]);
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[8];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = t[36] ^ x[16];
  assign t[31] = t[37] ^ x[17];
  assign t[32] = (~t[38] & t[39]);
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[42] & t[46]);
  assign t[38] = t[47] ^ x[4];
  assign t[39] = t[48] ^ x[5];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[8];
  assign t[42] = t[51] ^ x[13];
  assign t[43] = t[52] ^ x[14];
  assign t[44] = t[53] ^ x[15];
  assign t[45] = t[54] ^ x[16];
  assign t[46] = t[55] ^ x[17];
  assign t[47] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[48] = (x[0]);
  assign t[49] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[6]);
  assign t[51] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[52] = (x[10]);
  assign t[53] = (x[11]);
  assign t[54] = (x[9]);
  assign t[55] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[22] & t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = t[14] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind256(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind261(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind266(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [17:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] ^ t[32]);
  assign t[10] = ~(t[34]);
  assign t[11] = ~(t[33] ^ t[10]);
  assign t[12] = t[35] ^ t[34];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[33] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[33] ^ t[17];
  assign t[17] = t[34] ^ t[36];
  assign t[18] = ~(t[19] ^ t[37]);
  assign t[19] = ~t[20];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = t[23] ^ t[6];
  assign t[22] = t[3] ^ t[24];
  assign t[23] = t[12] ^ t[15];
  assign t[24] = t[33] ^ t[10];
  assign t[25] = ~(t[26] ^ t[38]);
  assign t[26] = ~t[27];
  assign t[27] = ~(t[28]);
  assign t[28] = t[17] ^ t[6];
  assign t[29] = ~(t[30] ^ t[39]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = ~t[31];
  assign t[31] = ~(t[21]);
  assign t[32] = (t[40]);
  assign t[33] = (t[41]);
  assign t[34] = (t[42]);
  assign t[35] = (t[43]);
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] ^ t[6];
  assign t[40] = t[48] ^ x[5];
  assign t[41] = t[49] ^ x[11];
  assign t[42] = t[50] ^ x[12];
  assign t[43] = t[51] ^ x[13];
  assign t[44] = t[52] ^ x[14];
  assign t[45] = t[53] ^ x[15];
  assign t[46] = t[54] ^ x[16];
  assign t[47] = t[55] ^ x[17];
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = t[7] & t[8];
  assign t[50] = (~t[58] & t[60]);
  assign t[51] = (~t[58] & t[61]);
  assign t[52] = (~t[58] & t[62]);
  assign t[53] = (~t[56] & t[63]);
  assign t[54] = (~t[56] & t[64]);
  assign t[55] = (~t[56] & t[65]);
  assign t[56] = t[66] ^ x[4];
  assign t[57] = t[67] ^ x[5];
  assign t[58] = t[68] ^ x[10];
  assign t[59] = t[69] ^ x[11];
  assign t[5] = t[33] & t[9];
  assign t[60] = t[70] ^ x[12];
  assign t[61] = t[71] ^ x[13];
  assign t[62] = t[72] ^ x[14];
  assign t[63] = t[73] ^ x[15];
  assign t[64] = t[74] ^ x[16];
  assign t[65] = t[75] ^ x[17];
  assign t[66] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[67] = (x[0]);
  assign t[68] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[69] = (x[7]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (x[8]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[1]);
  assign t[74] = (x[2]);
  assign t[75] = (x[3]);
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0] & ~t[18] & ~t[25] & ~t[29]) | (~t[0] & t[18] & ~t[25] & ~t[29]) | (~t[0] & ~t[18] & t[25] & ~t[29]) | (~t[0] & ~t[18] & ~t[25] & t[29]) | (t[0] & t[18] & t[25] & ~t[29]) | (t[0] & t[18] & ~t[25] & t[29]) | (t[0] & ~t[18] & t[25] & t[29]) | (~t[0] & t[18] & t[25] & t[29]);
endmodule

module R2ind271(x, y);
 input [14:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[13];
  assign t[21] = t[26] ^ x[14];
  assign t[22] = (~t[27] & t[28]);
  assign t[23] = (~t[29] & t[30]);
  assign t[24] = (~t[29] & t[31]);
  assign t[25] = (~t[29] & t[32]);
  assign t[26] = (~t[29] & t[33]);
  assign t[27] = t[34] ^ x[4];
  assign t[28] = t[35] ^ x[5];
  assign t[29] = t[36] ^ x[10];
  assign t[2] = ~(t[3]);
  assign t[30] = t[37] ^ x[11];
  assign t[31] = t[38] ^ x[12];
  assign t[32] = t[39] ^ x[13];
  assign t[33] = t[40] ^ x[14];
  assign t[34] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[35] = (x[3]);
  assign t[36] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[37] = (x[6]);
  assign t[38] = (x[8]);
  assign t[39] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[40] = (x[9]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [13:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[13];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[22] & t[24]);
  assign t[19] = (~t[22] & t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[4];
  assign t[21] = t[27] ^ x[5];
  assign t[22] = t[28] ^ x[10];
  assign t[23] = t[29] ^ x[11];
  assign t[24] = t[30] ^ x[12];
  assign t[25] = t[31] ^ x[13];
  assign t[26] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[27] = (x[2]);
  assign t[28] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[29] = (x[8]);
  assign t[2] = ~(t[3]);
  assign t[30] = (x[9]);
  assign t[31] = (x[7]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[1]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[6]);
  assign t[45] = (x[8]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [14:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[2];
  assign t[20] = (t[25]);
  assign t[21] = (t[26]);
  assign t[22] = (t[27]);
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[11];
  assign t[25] = t[30] ^ x[12];
  assign t[26] = t[31] ^ x[13];
  assign t[27] = t[32] ^ x[14];
  assign t[28] = (~t[33] & t[34]);
  assign t[29] = (~t[35] & t[36]);
  assign t[2] = t[3] ^ t[4];
  assign t[30] = (~t[35] & t[37]);
  assign t[31] = (~t[35] & t[38]);
  assign t[32] = (~t[35] & t[39]);
  assign t[33] = t[40] ^ x[4];
  assign t[34] = t[41] ^ x[5];
  assign t[35] = t[42] ^ x[10];
  assign t[36] = t[43] ^ x[11];
  assign t[37] = t[44] ^ x[12];
  assign t[38] = t[45] ^ x[13];
  assign t[39] = t[46] ^ x[14];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[41] = (x[0]);
  assign t[42] = (x[6] & ~x[7] & ~x[8] & ~x[9]) | (~x[6] & x[7] & ~x[8] & ~x[9]) | (~x[6] & ~x[7] & x[8] & ~x[9]) | (~x[6] & ~x[7] & ~x[8] & x[9]) | (x[6] & x[7] & x[8] & ~x[9]) | (x[6] & x[7] & ~x[8] & x[9]) | (x[6] & ~x[7] & x[8] & x[9]) | (~x[6] & x[7] & x[8] & x[9]);
  assign t[43] = (x[7]);
  assign t[44] = (x[8]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [29:0] x;
 output y;

 wire [111:0] t;
  assign t[0] = ~(t[1] ^ t[40]);
  assign t[100] = (x[11]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[1]);
  assign t[104] = (x[19] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[19] & 1'b0 & ~1'b0 & ~1'b0) | (~x[19] & ~1'b0 & 1'b0 & ~1'b0) | (~x[19] & ~1'b0 & ~1'b0 & 1'b0) | (x[19] & 1'b0 & 1'b0 & ~1'b0) | (x[19] & 1'b0 & ~1'b0 & 1'b0) | (x[19] & ~1'b0 & 1'b0 & 1'b0) | (~x[19] & 1'b0 & 1'b0 & 1'b0);
  assign t[105] = (x[19]);
  assign t[106] = (x[2]);
  assign t[107] = (x[23] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0 & ~1'b0) | (x[23] & 1'b0 & ~1'b0 & 1'b0) | (x[23] & ~1'b0 & 1'b0 & 1'b0) | (~x[23] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[23]);
  assign t[109] = (x[3]);
  assign t[10] = t[15] ^ t[8];
  assign t[110] = (x[27] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[27] & 1'b0 & ~1'b0 & ~1'b0) | (~x[27] & ~1'b0 & 1'b0 & ~1'b0) | (~x[27] & ~1'b0 & ~1'b0 & 1'b0) | (x[27] & 1'b0 & 1'b0 & ~1'b0) | (x[27] & 1'b0 & ~1'b0 & 1'b0) | (x[27] & ~1'b0 & 1'b0 & 1'b0) | (~x[27] & 1'b0 & 1'b0 & 1'b0);
  assign t[111] = (x[27]);
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[43]);
  assign t[13] = ~(t[42] ^ t[12]);
  assign t[14] = t[44] ^ t[43];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[42] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[42] ^ t[19];
  assign t[19] = t[43] ^ t[45];
  assign t[1] = ~t[2];
  assign t[20] = ~(t[21] ^ t[46]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[47]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = t[27] ^ t[8];
  assign t[26] = t[5] ^ t[28];
  assign t[27] = t[14] ^ t[17];
  assign t[28] = t[42] ^ t[12];
  assign t[29] = ~(t[30] ^ t[48]);
  assign t[2] = ~(t[3] ^ t[41]);
  assign t[30] = ~t[31];
  assign t[31] = ~(t[32] ^ t[49]);
  assign t[32] = ~t[33];
  assign t[33] = ~(t[34]);
  assign t[34] = t[19] ^ t[8];
  assign t[35] = ~(t[36] ^ t[50]);
  assign t[36] = ~t[37];
  assign t[37] = ~(t[38] ^ t[51]);
  assign t[38] = ~t[39];
  assign t[39] = ~(t[25]);
  assign t[3] = ~t[4];
  assign t[40] = (t[52]);
  assign t[41] = (t[53]);
  assign t[42] = (t[54]);
  assign t[43] = (t[55]);
  assign t[44] = (t[56]);
  assign t[45] = (t[57]);
  assign t[46] = (t[58]);
  assign t[47] = (t[59]);
  assign t[48] = (t[60]);
  assign t[49] = (t[61]);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (t[62]);
  assign t[51] = (t[63]);
  assign t[52] = t[64] ^ x[5];
  assign t[53] = t[65] ^ x[8];
  assign t[54] = t[66] ^ x[14];
  assign t[55] = t[67] ^ x[15];
  assign t[56] = t[68] ^ x[16];
  assign t[57] = t[69] ^ x[17];
  assign t[58] = t[70] ^ x[18];
  assign t[59] = t[71] ^ x[21];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[72] ^ x[22];
  assign t[61] = t[73] ^ x[25];
  assign t[62] = t[74] ^ x[26];
  assign t[63] = t[75] ^ x[29];
  assign t[64] = (~t[76] & t[77]);
  assign t[65] = (~t[78] & t[79]);
  assign t[66] = (~t[80] & t[81]);
  assign t[67] = (~t[80] & t[82]);
  assign t[68] = (~t[80] & t[83]);
  assign t[69] = (~t[80] & t[84]);
  assign t[6] = t[9] & t[10];
  assign t[70] = (~t[76] & t[85]);
  assign t[71] = (~t[86] & t[87]);
  assign t[72] = (~t[76] & t[88]);
  assign t[73] = (~t[89] & t[90]);
  assign t[74] = (~t[76] & t[91]);
  assign t[75] = (~t[92] & t[93]);
  assign t[76] = t[94] ^ x[4];
  assign t[77] = t[95] ^ x[5];
  assign t[78] = t[96] ^ x[7];
  assign t[79] = t[97] ^ x[8];
  assign t[7] = t[42] & t[11];
  assign t[80] = t[98] ^ x[13];
  assign t[81] = t[99] ^ x[14];
  assign t[82] = t[100] ^ x[15];
  assign t[83] = t[101] ^ x[16];
  assign t[84] = t[102] ^ x[17];
  assign t[85] = t[103] ^ x[18];
  assign t[86] = t[104] ^ x[20];
  assign t[87] = t[105] ^ x[21];
  assign t[88] = t[106] ^ x[22];
  assign t[89] = t[107] ^ x[24];
  assign t[8] = t[12] & t[13];
  assign t[90] = t[108] ^ x[25];
  assign t[91] = t[109] ^ x[26];
  assign t[92] = t[110] ^ x[28];
  assign t[93] = t[111] ^ x[29];
  assign t[94] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[95] = (x[0]);
  assign t[96] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[6]);
  assign t[98] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[99] = (x[10]);
  assign t[9] = t[14] ^ t[12];
  assign y = (t[0] & ~t[20] & ~t[29] & ~t[35]) | (~t[0] & t[20] & ~t[29] & ~t[35]) | (~t[0] & ~t[20] & t[29] & ~t[35]) | (~t[0] & ~t[20] & ~t[29] & t[35]) | (t[0] & t[20] & t[29] & ~t[35]) | (t[0] & t[20] & ~t[29] & t[35]) | (t[0] & ~t[20] & t[29] & t[35]) | (~t[0] & t[20] & t[29] & t[35]);
endmodule

module R2ind276(x, y);
 input [17:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[14]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] ^ t[13];
  assign t[13] = t[17] ^ t[19];
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = (t[22]);
  assign t[17] = (t[23]);
  assign t[18] = (t[24]);
  assign t[19] = (t[25]);
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[5];
  assign t[21] = t[27] ^ x[8];
  assign t[22] = t[28] ^ x[14];
  assign t[23] = t[29] ^ x[15];
  assign t[24] = t[30] ^ x[16];
  assign t[25] = t[31] ^ x[17];
  assign t[26] = (~t[32] & t[33]);
  assign t[27] = (~t[34] & t[35]);
  assign t[28] = (~t[36] & t[37]);
  assign t[29] = (~t[36] & t[38]);
  assign t[2] = ~(t[3] ^ t[15]);
  assign t[30] = (~t[36] & t[39]);
  assign t[31] = (~t[36] & t[40]);
  assign t[32] = t[41] ^ x[4];
  assign t[33] = t[42] ^ x[5];
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[8];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[14];
  assign t[38] = t[47] ^ x[15];
  assign t[39] = t[48] ^ x[16];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[17];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[3]);
  assign t[43] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[44] = (x[6]);
  assign t[45] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[46] = (x[9]);
  assign t[47] = (x[11]);
  assign t[48] = (x[10]);
  assign t[49] = (x[12]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[16] ^ t[17];
  assign t[9] = t[10] & t[12];
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [16:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[10]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[14];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = t[24] ^ x[16];
  assign t[1] = ~t[2];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = (~t[29] & t[31]);
  assign t[24] = (~t[29] & t[32]);
  assign t[25] = t[33] ^ x[4];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[7];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[13];
  assign t[2] = ~(t[3] ^ t[11]);
  assign t[30] = t[38] ^ x[14];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[16];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[2]);
  assign t[35] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[6]);
  assign t[37] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[38] = (x[11]);
  assign t[39] = (x[12]);
  assign t[3] = ~t[4];
  assign t[40] = (x[10]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[12] ^ t[13];
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[14] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [17:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[22] ^ t[13];
  assign t[11] = t[23] ^ t[24];
  assign t[12] = t[13] & t[16];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[22] ^ t[13]);
  assign t[15] = t[22] & t[17];
  assign t[16] = t[22] ^ t[18];
  assign t[17] = t[19] ^ t[12];
  assign t[18] = t[24] ^ t[25];
  assign t[19] = t[22] ^ t[11];
  assign t[1] = ~t[2];
  assign t[20] = (t[26]);
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[8];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = t[36] ^ x[16];
  assign t[31] = t[37] ^ x[17];
  assign t[32] = (~t[38] & t[39]);
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[42] & t[46]);
  assign t[38] = t[47] ^ x[4];
  assign t[39] = t[48] ^ x[5];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[8];
  assign t[42] = t[51] ^ x[13];
  assign t[43] = t[52] ^ x[14];
  assign t[44] = t[53] ^ x[15];
  assign t[45] = t[54] ^ x[16];
  assign t[46] = t[55] ^ x[17];
  assign t[47] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[48] = (x[1]);
  assign t[49] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = ~(t[5] ^ t[6]);
  assign t[50] = (x[6]);
  assign t[51] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[52] = (x[10]);
  assign t[53] = (x[9]);
  assign t[54] = (x[11]);
  assign t[55] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[8];
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [17:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[22] ^ t[12]);
  assign t[14] = t[24] ^ t[23];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[22] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[22] ^ t[19];
  assign t[19] = t[23] ^ t[25];
  assign t[1] = ~t[2];
  assign t[20] = (t[26]);
  assign t[21] = (t[27]);
  assign t[22] = (t[28]);
  assign t[23] = (t[29]);
  assign t[24] = (t[30]);
  assign t[25] = (t[31]);
  assign t[26] = t[32] ^ x[5];
  assign t[27] = t[33] ^ x[8];
  assign t[28] = t[34] ^ x[14];
  assign t[29] = t[35] ^ x[15];
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = t[36] ^ x[16];
  assign t[31] = t[37] ^ x[17];
  assign t[32] = (~t[38] & t[39]);
  assign t[33] = (~t[40] & t[41]);
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[42] & t[44]);
  assign t[36] = (~t[42] & t[45]);
  assign t[37] = (~t[42] & t[46]);
  assign t[38] = t[47] ^ x[4];
  assign t[39] = t[48] ^ x[5];
  assign t[3] = ~t[4];
  assign t[40] = t[49] ^ x[7];
  assign t[41] = t[50] ^ x[8];
  assign t[42] = t[51] ^ x[13];
  assign t[43] = t[52] ^ x[14];
  assign t[44] = t[53] ^ x[15];
  assign t[45] = t[54] ^ x[16];
  assign t[46] = t[55] ^ x[17];
  assign t[47] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[48] = (x[0]);
  assign t[49] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[4] = t[5] ^ t[6];
  assign t[50] = (x[6]);
  assign t[51] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[52] = (x[10]);
  assign t[53] = (x[11]);
  assign t[54] = (x[9]);
  assign t[55] = (x[12]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[22] & t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = t[14] ^ t[12];
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind281(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind286(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind291(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [8:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[26] ^ t[25];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[24] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[24] ^ t[15];
  assign t[15] = t[25] ^ t[27];
  assign t[16] = ~(t[17] ^ t[18]);
  assign t[17] = t[19] ^ t[4];
  assign t[18] = t[1] ^ t[20];
  assign t[19] = t[10] ^ t[13];
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ t[8];
  assign t[21] = ~(t[22]);
  assign t[22] = t[15] ^ t[4];
  assign t[23] = ~(t[17]);
  assign t[24] = (t[28]);
  assign t[25] = (t[29]);
  assign t[26] = (t[30]);
  assign t[27] = (t[31]);
  assign t[28] = t[32] ^ x[5];
  assign t[29] = t[33] ^ x[6];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[34] ^ x[7];
  assign t[31] = t[35] ^ x[8];
  assign t[32] = (~t[36] & t[37]);
  assign t[33] = (~t[36] & t[38]);
  assign t[34] = (~t[36] & t[39]);
  assign t[35] = (~t[36] & t[40]);
  assign t[36] = t[41] ^ x[4];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[6];
  assign t[39] = t[44] ^ x[7];
  assign t[3] = t[24] & t[7];
  assign t[40] = t[45] ^ x[8];
  assign t[41] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[42] = (x[1]);
  assign t[43] = (x[2]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[25]);
  assign t[9] = ~(t[24] ^ t[8]);
  assign y = (t[0] & ~t[16] & ~t[21] & ~t[23]) | (~t[0] & t[16] & ~t[21] & ~t[23]) | (~t[0] & ~t[16] & t[21] & ~t[23]) | (~t[0] & ~t[16] & ~t[21] & t[23]) | (t[0] & t[16] & t[21] & ~t[23]) | (t[0] & t[16] & ~t[21] & t[23]) | (t[0] & ~t[16] & t[21] & t[23]) | (~t[0] & t[16] & t[21] & t[23]);
endmodule

module R2ind296(x, y);
 input [8:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[5];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[7];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[4];
  assign t[23] = t[28] ^ x[5];
  assign t[24] = t[29] ^ x[6];
  assign t[25] = t[30] ^ x[7];
  assign t[26] = t[31] ^ x[8];
  assign t[27] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (x[1]);
  assign t[31] = (x[3]);
  assign t[3] = t[6] & t[7];
  assign t[4] = t[10] ^ t[11];
  assign t[5] = t[6] & t[8];
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[12] ^ t[6]);
  assign t[8] = t[12] ^ t[9];
  assign t[9] = t[11] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = t[2] ^ t[3];
  assign t[20] = (x[2]);
  assign t[21] = (x[3]);
  assign t[22] = (x[1]);
  assign t[2] = t[6] ^ t[7];
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[8] ^ t[4]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] ^ t[9]);
  assign t[11] = t[16] & t[13];
  assign t[12] = t[16] ^ t[14];
  assign t[13] = t[15] ^ t[8];
  assign t[14] = t[18] ^ t[19];
  assign t[15] = t[16] ^ t[7];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[0]);
  assign t[36] = (x[2]);
  assign t[37] = (x[3]);
  assign t[3] = t[7] ^ t[8];
  assign t[4] = t[9] & t[10];
  assign t[5] = t[11] ^ t[4];
  assign t[6] = t[16] ^ t[9];
  assign t[7] = t[17] ^ t[18];
  assign t[8] = t[9] & t[12];
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [8:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[18] ^ t[17];
  assign t[11] = ~(t[14] ^ t[5]);
  assign t[12] = t[16] ^ t[10];
  assign t[13] = t[8] & t[14];
  assign t[14] = t[16] ^ t[15];
  assign t[15] = t[17] ^ t[19];
  assign t[16] = (t[20]);
  assign t[17] = (t[21]);
  assign t[18] = (t[22]);
  assign t[19] = (t[23]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = t[24] ^ x[5];
  assign t[21] = t[25] ^ x[6];
  assign t[22] = t[26] ^ x[7];
  assign t[23] = t[27] ^ x[8];
  assign t[24] = (~t[28] & t[29]);
  assign t[25] = (~t[28] & t[30]);
  assign t[26] = (~t[28] & t[31]);
  assign t[27] = (~t[28] & t[32]);
  assign t[28] = t[33] ^ x[4];
  assign t[29] = t[34] ^ x[5];
  assign t[2] = t[5] & t[6];
  assign t[30] = t[35] ^ x[6];
  assign t[31] = t[36] ^ x[7];
  assign t[32] = t[37] ^ x[8];
  assign t[33] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[34] = (x[1]);
  assign t[35] = (x[2]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[3] = t[16] & t[7];
  assign t[4] = t[8] & t[9];
  assign t[5] = t[10] ^ t[8];
  assign t[6] = t[11] ^ t[4];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[17]);
  assign t[9] = ~(t[16] ^ t[8]);
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [556:0] x;
 output [299:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[23], x[22], x[21], x[11], x[10], x[9], x[8], x[7], x[6], x[24]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[23], x[22], x[21], x[11], x[10], x[9], x[8], x[7], x[6], x[24]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[23], x[22], x[21], x[24]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[23], x[22], x[21], x[24]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[23], x[22], x[21], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[24]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[20], x[19], x[18], x[17], x[16], x[15], x[23], x[22], x[21], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[24]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[17], x[16], x[15], x[24]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[17], x[16], x[15], x[24]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[20], x[19], x[18], x[24]}), .y(y[30]));
  R2ind31 R2ind31_inst(.y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.x({x[20], x[19], x[18], x[24]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[14], x[13], x[12], x[23], x[22], x[21], x[17], x[16], x[15], x[11], x[10], x[9], x[20], x[19], x[18], x[8], x[7], x[6], x[24]}), .y(y[35]));
  R2ind36 R2ind36_inst(.y(y[36]));
  R2ind37 R2ind37_inst(.y(y[37]));
  R2ind38 R2ind38_inst(.y(y[38]));
  R2ind39 R2ind39_inst(.x({x[14], x[13], x[12], x[23], x[22], x[21], x[17], x[16], x[15], x[11], x[10], x[9], x[20], x[19], x[18], x[8], x[7], x[6], x[24]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[24], x[27], x[26], x[25]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[24], x[30], x[29], x[28]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[24], x[33], x[32], x[31]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[24], x[36], x[35], x[34]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[24], x[39], x[38], x[37]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[24], x[42], x[41], x[40]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[24], x[45], x[44], x[43]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[24], x[48], x[47], x[46]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[24], x[51], x[50], x[49]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[24], x[54], x[53], x[52]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[24], x[57], x[56], x[55]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[24], x[60], x[59], x[58]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[24], x[63], x[62], x[61]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[24], x[66], x[65], x[64]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[24], x[69], x[68], x[67]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[24], x[72], x[71], x[70]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[24], x[75], x[74], x[73]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[24], x[78], x[77], x[76]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[24], x[81], x[80], x[79]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[24], x[84], x[83], x[82]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[24], x[86], x[27], x[85]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[24], x[88], x[30], x[87]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[24], x[90], x[33], x[89]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[24], x[92], x[36], x[91]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[24], x[94], x[39], x[93]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[24], x[96], x[42], x[95]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[24], x[98], x[45], x[97]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[24], x[100], x[48], x[99]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[24], x[102], x[51], x[101]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[24], x[104], x[54], x[103]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[24], x[106], x[57], x[105]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[24], x[108], x[60], x[107]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[24], x[110], x[63], x[109]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[24], x[112], x[66], x[111]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[24], x[114], x[69], x[113]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[24], x[116], x[72], x[115]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[24], x[118], x[75], x[117]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[24], x[120], x[78], x[119]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[24], x[122], x[81], x[121]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[24], x[124], x[84], x[123]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[24], x[126], x[125]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[24], x[128], x[127]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[24], x[130], x[129]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[24], x[132], x[131]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[24], x[134], x[133]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[24], x[136], x[135]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[24], x[138], x[137]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[24], x[140], x[139]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[24], x[142], x[141]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[24], x[144], x[143]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[24], x[146], x[145]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[24], x[148], x[147]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[24], x[150], x[149]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[24], x[152], x[151]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[24], x[154], x[153]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[24], x[156], x[155]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[24], x[158], x[157]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[24], x[160], x[159]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[24], x[162], x[161]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[24], x[164], x[163]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[24], x[27], x[166], x[165], x[25]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[24], x[30], x[168], x[167], x[28]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[24], x[33], x[170], x[169], x[31]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[24], x[36], x[172], x[171], x[34]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[24], x[39], x[174], x[173], x[37]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[24], x[176], x[42], x[175], x[40]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[24], x[178], x[45], x[177], x[43]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[24], x[180], x[48], x[179], x[46]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[24], x[182], x[51], x[181], x[49]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[24], x[184], x[54], x[183], x[52]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[24], x[186], x[57], x[185], x[55]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[24], x[188], x[60], x[187], x[58]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[24], x[190], x[63], x[189], x[61]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[24], x[192], x[66], x[191], x[64]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[24], x[194], x[69], x[193], x[67]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[24], x[72], x[196], x[195], x[70]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[24], x[75], x[198], x[197], x[73]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[24], x[78], x[200], x[199], x[76]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[24], x[81], x[202], x[201], x[79]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[24], x[84], x[204], x[203], x[82]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[24]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[217], x[216], x[209], x[208], x[207], x[206], x[205], x[24]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[215], x[214], x[209], x[208], x[207], x[206], x[205], x[24]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[213], x[212], x[209], x[208], x[207], x[206], x[205], x[24]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[24]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[24]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[230], x[229], x[222], x[221], x[220], x[219], x[218], x[24]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[228], x[227], x[222], x[221], x[220], x[219], x[218], x[24]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[226], x[225], x[222], x[221], x[220], x[219], x[218], x[24]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[24]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[24]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[243], x[242], x[235], x[234], x[233], x[232], x[231], x[24]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[241], x[240], x[235], x[234], x[233], x[232], x[231], x[24]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[239], x[238], x[235], x[234], x[233], x[232], x[231], x[24]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[24]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[24]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[256], x[255], x[248], x[247], x[246], x[245], x[244], x[24]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[254], x[253], x[248], x[247], x[246], x[245], x[244], x[24]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[252], x[251], x[248], x[247], x[246], x[245], x[244], x[24]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[24]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[24]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[269], x[268], x[261], x[260], x[259], x[258], x[257], x[24]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[267], x[266], x[261], x[260], x[259], x[258], x[257], x[24]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[265], x[264], x[261], x[260], x[259], x[258], x[257], x[24]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[24]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[24]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[282], x[281], x[274], x[273], x[272], x[271], x[270], x[24]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[280], x[279], x[274], x[273], x[272], x[271], x[270], x[24]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[278], x[277], x[274], x[273], x[272], x[271], x[270], x[24]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[24]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[295], x[294], x[293], x[292], x[291], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[24]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[295], x[294], x[287], x[286], x[285], x[284], x[283], x[24]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[293], x[292], x[287], x[286], x[285], x[284], x[283], x[24]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[291], x[290], x[287], x[286], x[285], x[284], x[283], x[24]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[24]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[24]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[308], x[307], x[300], x[299], x[298], x[297], x[296], x[24]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[306], x[305], x[300], x[299], x[298], x[297], x[296], x[24]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[304], x[303], x[300], x[299], x[298], x[297], x[296], x[24]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[24]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[24]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[321], x[320], x[313], x[312], x[311], x[310], x[309], x[24]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[319], x[318], x[313], x[312], x[311], x[310], x[309], x[24]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[317], x[316], x[313], x[312], x[311], x[310], x[309], x[24]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[24]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[24]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[334], x[333], x[326], x[325], x[324], x[323], x[322], x[24]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[332], x[331], x[326], x[325], x[324], x[323], x[322], x[24]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[330], x[329], x[326], x[325], x[324], x[323], x[322], x[24]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[328], x[327], x[326], x[325], x[324], x[323], x[322], x[24]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[24]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[347], x[346], x[339], x[338], x[337], x[336], x[335], x[24]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[345], x[344], x[339], x[338], x[337], x[336], x[335], x[24]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[343], x[342], x[339], x[338], x[337], x[336], x[335], x[24]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[24]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[24]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[360], x[359], x[352], x[351], x[350], x[349], x[348], x[24]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[358], x[357], x[352], x[351], x[350], x[349], x[348], x[24]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[356], x[355], x[352], x[351], x[350], x[349], x[348], x[24]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[354], x[353], x[352], x[351], x[350], x[349], x[348], x[24]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[373], x[372], x[371], x[370], x[369], x[368], x[367], x[366], x[365], x[364], x[363], x[362], x[361], x[24]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[373], x[372], x[365], x[364], x[363], x[362], x[361], x[24]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[371], x[370], x[365], x[364], x[363], x[362], x[361], x[24]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[369], x[368], x[365], x[364], x[363], x[362], x[361], x[24]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[367], x[366], x[365], x[364], x[363], x[362], x[361], x[24]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[377], x[376], x[375], x[374], x[24]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[386], x[385], x[378], x[377], x[376], x[375], x[374], x[24]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[384], x[383], x[378], x[377], x[376], x[375], x[374], x[24]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[382], x[381], x[378], x[377], x[376], x[375], x[374], x[24]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[380], x[379], x[378], x[377], x[376], x[375], x[374], x[24]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[24]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[399], x[398], x[391], x[390], x[389], x[388], x[387], x[24]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[397], x[396], x[391], x[390], x[389], x[388], x[387], x[24]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[395], x[394], x[391], x[390], x[389], x[388], x[387], x[24]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[24]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[24]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[24]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[410], x[409], x[404], x[403], x[402], x[401], x[400], x[24]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[408], x[407], x[404], x[403], x[402], x[401], x[400], x[24]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[24]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[421], x[418], x[419], x[420], x[417], x[416], x[415], x[414], x[413]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[418], x[421], x[419], x[417], x[416], x[415], x[414], x[413]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[421], x[419], x[420], x[418], x[417], x[416], x[415], x[414], x[413]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[268], x[266], x[264], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[430], x[427], x[428], x[429], x[426], x[425], x[424], x[423], x[422], x[268], x[261], x[260], x[259], x[258], x[257]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[427], x[430], x[428], x[426], x[425], x[424], x[423], x[422], x[266], x[261], x[260], x[259], x[258], x[257]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[430], x[428], x[429], x[427], x[426], x[425], x[424], x[423], x[422], x[264], x[261], x[260], x[259], x[258], x[257]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[431]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[439], x[436], x[437], x[438], x[435], x[434], x[433], x[432], x[431]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[436], x[439], x[437], x[435], x[434], x[433], x[432], x[431]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[439], x[437], x[438], x[436], x[435], x[434], x[433], x[432], x[431]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[431]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[281], x[279], x[277], x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[275], x[274], x[273], x[272], x[271], x[270]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[448], x[445], x[446], x[447], x[444], x[443], x[442], x[441], x[440], x[281], x[274], x[273], x[272], x[271], x[270]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[445], x[448], x[446], x[444], x[443], x[442], x[441], x[440], x[279], x[274], x[273], x[272], x[271], x[270]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[448], x[446], x[447], x[445], x[444], x[443], x[442], x[441], x[440], x[277], x[274], x[273], x[272], x[271], x[270]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[275], x[274], x[273], x[272], x[271], x[270]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[457], x[456], x[455], x[454], x[453], x[452], x[451], x[450], x[449]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[457], x[454], x[455], x[456], x[453], x[452], x[451], x[450], x[449]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[454], x[457], x[455], x[453], x[452], x[451], x[450], x[449]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[457], x[455], x[456], x[454], x[453], x[452], x[451], x[450], x[449]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[457], x[456], x[455], x[454], x[453], x[452], x[451], x[450], x[449]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[294], x[292], x[290], x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[288], x[287], x[286], x[285], x[284], x[283]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[466], x[463], x[464], x[465], x[462], x[461], x[460], x[459], x[458], x[294], x[287], x[286], x[285], x[284], x[283]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[463], x[466], x[464], x[462], x[461], x[460], x[459], x[458], x[292], x[287], x[286], x[285], x[284], x[283]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[466], x[464], x[465], x[463], x[462], x[461], x[460], x[459], x[458], x[290], x[287], x[286], x[285], x[284], x[283]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[288], x[287], x[286], x[285], x[284], x[283]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[467]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[475], x[472], x[473], x[474], x[471], x[470], x[469], x[468], x[467]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[472], x[475], x[473], x[471], x[470], x[469], x[468], x[467]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[475], x[473], x[474], x[472], x[471], x[470], x[469], x[468], x[467]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[467]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[20], x[19], x[18], x[307], x[17], x[16], x[15], x[305], x[14], x[13], x[12], x[303], x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[476], x[23], x[22], x[21], x[301], x[300], x[299], x[298], x[297], x[296]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[484], x[481], x[482], x[483], x[480], x[479], x[478], x[477], x[476], x[20], x[19], x[18], x[307], x[300], x[299], x[298], x[297], x[296]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[481], x[484], x[482], x[480], x[479], x[478], x[477], x[476], x[17], x[16], x[15], x[305], x[300], x[299], x[298], x[297], x[296]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[484], x[482], x[483], x[481], x[480], x[479], x[478], x[477], x[476], x[14], x[13], x[12], x[303], x[300], x[299], x[298], x[297], x[296]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[476], x[23], x[22], x[21], x[301], x[300], x[299], x[298], x[297], x[296]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[229], x[227], x[225], x[493], x[492], x[491], x[490], x[489], x[488], x[487], x[486], x[485], x[223], x[222], x[221], x[220], x[219], x[218]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[493], x[490], x[491], x[492], x[489], x[488], x[487], x[486], x[485], x[229], x[222], x[221], x[220], x[219], x[218]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[490], x[493], x[491], x[489], x[488], x[487], x[486], x[485], x[227], x[222], x[221], x[220], x[219], x[218]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[493], x[491], x[492], x[490], x[489], x[488], x[487], x[486], x[485], x[225], x[222], x[221], x[220], x[219], x[218]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[493], x[492], x[491], x[490], x[489], x[488], x[487], x[486], x[485], x[223], x[222], x[221], x[220], x[219], x[218]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[242], x[240], x[238], x[502], x[501], x[500], x[499], x[498], x[497], x[496], x[495], x[494], x[236], x[235], x[234], x[233], x[232], x[231]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[502], x[499], x[500], x[501], x[498], x[497], x[496], x[495], x[494], x[242], x[235], x[234], x[233], x[232], x[231]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[499], x[502], x[500], x[498], x[497], x[496], x[495], x[494], x[240], x[235], x[234], x[233], x[232], x[231]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[502], x[500], x[501], x[499], x[498], x[497], x[496], x[495], x[494], x[238], x[235], x[234], x[233], x[232], x[231]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[502], x[501], x[500], x[499], x[498], x[497], x[496], x[495], x[494], x[236], x[235], x[234], x[233], x[232], x[231]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[255], x[253], x[11], x[10], x[9], x[251], x[511], x[510], x[509], x[508], x[507], x[506], x[505], x[504], x[503], x[8], x[7], x[6], x[249], x[248], x[247], x[246], x[245], x[244]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[511], x[508], x[509], x[510], x[507], x[506], x[505], x[504], x[503], x[255], x[248], x[247], x[246], x[245], x[244]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[508], x[511], x[509], x[507], x[506], x[505], x[504], x[503], x[253], x[248], x[247], x[246], x[245], x[244]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[511], x[509], x[510], x[508], x[507], x[506], x[505], x[504], x[503], x[11], x[10], x[9], x[251], x[248], x[247], x[246], x[245], x[244]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[511], x[510], x[509], x[508], x[507], x[506], x[505], x[504], x[503], x[8], x[7], x[6], x[249], x[248], x[247], x[246], x[245], x[244]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[216], x[214], x[212], x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[210], x[209], x[208], x[207], x[206], x[205]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[520], x[517], x[518], x[519], x[516], x[515], x[514], x[513], x[512], x[216], x[209], x[208], x[207], x[206], x[205]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[517], x[520], x[518], x[516], x[515], x[514], x[513], x[512], x[214], x[209], x[208], x[207], x[206], x[205]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[520], x[518], x[519], x[517], x[516], x[515], x[514], x[513], x[512], x[212], x[209], x[208], x[207], x[206], x[205]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[210], x[209], x[208], x[207], x[206], x[205]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[268], x[266], x[264], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[430], x[427], x[428], x[429], x[426], x[425], x[424], x[423], x[422], x[268], x[261], x[260], x[259], x[258], x[257]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[427], x[430], x[428], x[426], x[425], x[424], x[423], x[422], x[266], x[261], x[260], x[259], x[258], x[257]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[430], x[428], x[429], x[427], x[426], x[425], x[424], x[423], x[422], x[264], x[261], x[260], x[259], x[258], x[257]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[281], x[279], x[277], x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[275], x[274], x[273], x[272], x[271], x[270]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[448], x[445], x[446], x[447], x[444], x[443], x[442], x[441], x[440], x[281], x[274], x[273], x[272], x[271], x[270]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[445], x[448], x[446], x[444], x[443], x[442], x[441], x[440], x[279], x[274], x[273], x[272], x[271], x[270]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[448], x[446], x[447], x[445], x[444], x[443], x[442], x[441], x[440], x[277], x[274], x[273], x[272], x[271], x[270]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[448], x[447], x[446], x[445], x[444], x[443], x[442], x[441], x[440], x[275], x[274], x[273], x[272], x[271], x[270]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[294], x[292], x[290], x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[288], x[287], x[286], x[285], x[284], x[283]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[466], x[463], x[464], x[465], x[462], x[461], x[460], x[459], x[458], x[294], x[287], x[286], x[285], x[284], x[283]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[463], x[466], x[464], x[462], x[461], x[460], x[459], x[458], x[292], x[287], x[286], x[285], x[284], x[283]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[466], x[464], x[465], x[463], x[462], x[461], x[460], x[459], x[458], x[290], x[287], x[286], x[285], x[284], x[283]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[288], x[287], x[286], x[285], x[284], x[283]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[20], x[19], x[18], x[307], x[17], x[16], x[15], x[305], x[14], x[13], x[12], x[303], x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[476], x[23], x[22], x[21], x[301], x[300], x[299], x[298], x[297], x[296]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[484], x[481], x[482], x[483], x[480], x[479], x[478], x[477], x[476], x[20], x[19], x[18], x[307], x[300], x[299], x[298], x[297], x[296]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[481], x[484], x[482], x[480], x[479], x[478], x[477], x[476], x[17], x[16], x[15], x[305], x[300], x[299], x[298], x[297], x[296]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[484], x[482], x[483], x[481], x[480], x[479], x[478], x[477], x[476], x[14], x[13], x[12], x[303], x[300], x[299], x[298], x[297], x[296]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[476], x[23], x[22], x[21], x[301], x[300], x[299], x[298], x[297], x[296]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[529], x[528], x[527], x[526], x[525], x[524], x[523], x[522], x[521]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[529], x[526], x[527], x[528], x[525], x[524], x[523], x[522], x[521]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[526], x[529], x[527], x[525], x[524], x[523], x[522], x[521]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[529], x[527], x[528], x[526], x[525], x[524], x[523], x[522], x[521]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[529], x[528], x[527], x[526], x[525], x[524], x[523], x[522], x[521]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[538], x[537], x[536], x[535], x[534], x[533], x[532], x[531], x[530]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[538], x[535], x[536], x[537], x[534], x[533], x[532], x[531], x[530]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[535], x[538], x[536], x[534], x[533], x[532], x[531], x[530]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[538], x[536], x[537], x[535], x[534], x[533], x[532], x[531], x[530]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[538], x[537], x[536], x[535], x[534], x[533], x[532], x[531], x[530]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[547], x[544], x[545], x[546], x[543], x[542], x[541], x[540], x[539]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[544], x[547], x[545], x[543], x[542], x[541], x[540], x[539]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[547], x[545], x[546], x[544], x[543], x[542], x[541], x[540], x[539]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[547], x[546], x[545], x[544], x[543], x[542], x[541], x[540], x[539]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[556], x[555], x[554], x[553], x[552], x[551], x[550], x[549], x[548]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[556], x[553], x[554], x[555], x[552], x[551], x[550], x[549], x[548]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[553], x[556], x[554], x[552], x[551], x[550], x[549], x[548]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[556], x[554], x[555], x[553], x[552], x[551], x[550], x[549], x[548]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[556], x[555], x[554], x[553], x[552], x[551], x[550], x[549], x[548]}), .y(y[299]));
endmodule

