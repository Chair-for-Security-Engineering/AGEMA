module Reg1(x, y);
 input [74:0] x;
 output [73:0] y;

  register_stage #(.WIDTH(74)) inst_0(.clk(x[71]), .D({x[72],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[73],x[74],x[0],x[11],x[22],x[33],x[44],x[55],x[60],x[61],x[62],x[63],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[56],x[57],x[58],x[59]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73]}));
endmodule

module Reg2(x, y);
 input [148:0] x;
 output [147:0] y;

  register_stage #(.WIDTH(148)) inst_0(.clk(x[142]), .D({x[143],x[144],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[145],x[146],x[147],x[148],x[0],x[1],x[22],x[23],x[44],x[45],x[66],x[67],x[88],x[89],x[110],x[111],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [221:0] x;
 output [147:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[79], x[78]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[80], x[78]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[82], x[81]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[83], x[81]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[85], x[84]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[86], x[84]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[88], x[87]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[89], x[87]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[91], x[90]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[92], x[90]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[94], x[93]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[95], x[93]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[97], x[96]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[98], x[96]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[100], x[99]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[101], x[99]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[103], x[102]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[104], x[102]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[106], x[105]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[107], x[105]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[109], x[108]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[110], x[108]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[112], x[111]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[113], x[111]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[115], x[114]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[116], x[114]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[118], x[117]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[119], x[117]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[121], x[120]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[122], x[120]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[124], x[123]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[125], x[123]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[127], x[126]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[128], x[126]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[130], x[129]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[131], x[129]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[133], x[132]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[134], x[132]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[136], x[135]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[139], x[138]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[140], x[138]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[142], x[141]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[143], x[141]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[145], x[144]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[146], x[144]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[148], x[147]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[149], x[147]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[151], x[150]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[152], x[150]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[154], x[153]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[155], x[153]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[157], x[156]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[158], x[156]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[160], x[159]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[161], x[159]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[163], x[162]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[164], x[162]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[166], x[165]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[167], x[165]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[169], x[168]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[170], x[168]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[172], x[171]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[173], x[171]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[175], x[174]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[176], x[174]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[178], x[177]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[179], x[177]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[181], x[180]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[182], x[180]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[184], x[183]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[185], x[183]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[187], x[186]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[188], x[186]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[190], x[189]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[191], x[189]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[193], x[192]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[194], x[192]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[196], x[195]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[199], x[198]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[200], x[198]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[202], x[201]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[203], x[201]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[205], x[204]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[206], x[204]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[208], x[207]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[209], x[207]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[211], x[210]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[212], x[210]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[214], x[213]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[215], x[213]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[217], x[216]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[218], x[216]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[220], x[219]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[221], x[219]}), .y(y[147]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [21:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~x[0] & t[12];
  assign t[10] = ~x[0] & t[17];
  assign t[11] = ~x[0] & t[18];
  assign t[12] = t[19] ^ x[3];
  assign t[13] = t[20] ^ x[6];
  assign t[14] = t[21] ^ x[9];
  assign t[15] = t[22] ^ x[12];
  assign t[16] = t[23] ^ x[15];
  assign t[17] = t[24] ^ x[18];
  assign t[18] = t[25] ^ x[21];
  assign t[19] = (x[1] & x[2]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[20] = (x[4] & x[5]);
  assign t[21] = (x[7] & x[8]);
  assign t[22] = (x[10] & x[11]);
  assign t[23] = (x[13] & x[14]);
  assign t[24] = (x[16] & x[17]);
  assign t[25] = (x[19] & x[20]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[7]);
  assign t[4] = ~(~x[0] & ~t[13]);
  assign t[5] = ~x[0] & t[14];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~x[0] & t[15];
  assign t[9] = ~(~x[0] & ~t[16]);
  assign y = t[0] & t[1];
endmodule

module R1ind66(x, y);
 input [3:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = t[2] ^ x[3];
  assign t[2] = (x[1] & x[2]);
  assign y = ~(t[0]);
endmodule

module R1ind67(x, y);
 input [6:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = ~t[2];
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = t[5] ^ x[3];
  assign t[4] = t[6] ^ x[6];
  assign t[5] = (x[1] & x[2]);
  assign t[6] = (x[4] & x[5]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind68(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~x[0] & t[2];
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = t[4] ^ x[3];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[1] & x[2]);
  assign t[5] = (x[4] & x[5]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind73(x, y);
 input [3:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[3];
  assign t[1] = (x[1] & x[2]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind74(x, y);
 input [6:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = ~(~x[0] & ~t[2]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = t[4] ^ x[3];
  assign t[3] = t[5] ^ x[6];
  assign t[4] = (x[1] & x[2]);
  assign t[5] = (x[4] & x[5]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [18:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[12];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = t[21] ^ x[18];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[10] & x[11]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & x[14]);
  assign t[21] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[13] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] | t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind76(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind77(x, y);
 input [18:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[12];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = t[21] ^ x[18];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[10] & x[11]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & x[14]);
  assign t[21] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind78(x, y);
 input [18:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[12];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = t[22] ^ x[18];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[10] & x[11]);
  assign t[21] = (x[13] & x[14]);
  assign t[22] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind79(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind80(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind81(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind82(x, y);
 input [18:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[12];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = t[22] ^ x[18];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[10] & x[11]);
  assign t[21] = (x[13] & x[14]);
  assign t[22] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind83(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind84(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind85(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind86(x, y);
 input [18:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[12];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = t[22] ^ x[18];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[10] & x[11]);
  assign t[21] = (x[13] & x[14]);
  assign t[22] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind87(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind88(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind89(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind90(x, y);
 input [18:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[12];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = t[22] ^ x[18];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[10] & x[11]);
  assign t[21] = (x[13] & x[14]);
  assign t[22] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind91(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind92(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind93(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind94(x, y);
 input [18:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[12];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = t[22] ^ x[18];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[10] & x[11]);
  assign t[21] = (x[13] & x[14]);
  assign t[22] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind95(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind96(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind97(x, y);
 input [18:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[12];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = t[21] ^ x[18];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[10] & x[11]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & x[14]);
  assign t[21] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind98(x, y);
 input [18:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15]);
  assign t[11] = t[16] ^ x[6];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[12];
  assign t[14] = t[19] ^ x[15];
  assign t[15] = t[20] ^ x[18];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[11];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = t[9] | t[12];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[10] | t[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind99(x, y);
 input [18:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[12];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = t[21] ^ x[18];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[10] & x[11]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & x[14]);
  assign t[21] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[13] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] | t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind100(x, y);
 input [15:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~t[2];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[9];
  assign t[12] = t[16] ^ x[12];
  assign t[13] = t[17] ^ x[15];
  assign t[14] = (x[4] & x[5]);
  assign t[15] = (x[7] & x[8]);
  assign t[16] = (x[10] & x[11]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[10];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[11] & t[7]);
  assign t[6] = ~(t[12] & t[8]);
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[13] & t[9]);
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind101(x, y);
 input [18:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[14]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[17] ^ x[6];
  assign t[13] = t[18] ^ x[9];
  assign t[14] = t[19] ^ x[12];
  assign t[15] = t[20] ^ x[15];
  assign t[16] = t[21] ^ x[18];
  assign t[17] = (x[4] & x[5]);
  assign t[18] = (x[7] & x[8]);
  assign t[19] = (x[10] & x[11]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[13] & x[14]);
  assign t[21] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[12];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9] & t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind102(x, y);
 input [18:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15]);
  assign t[11] = t[16] ^ x[6];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[12];
  assign t[14] = t[19] ^ x[15];
  assign t[15] = t[20] ^ x[18];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~x[2] & t[11];
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = t[9] | t[12];
  assign t[7] = ~(t[13]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[10] | t[7]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind103(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] | t[13]);
  assign t[12] = ~(t[18]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[14] | t[11]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind104(x, y);
 input [15:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[15] & t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = t[19] ^ x[15];
  assign t[16] = (x[4] & x[5]);
  assign t[17] = (x[7] & x[8]);
  assign t[18] = (x[10] & x[11]);
  assign t[19] = (x[13] & x[14]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[12] & t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind105(x, y);
 input [18:0] x;
 output y;

 wire [23:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[17] & t[16]);
  assign t[13] = ~(t[18]);
  assign t[14] = t[19] ^ x[6];
  assign t[15] = t[20] ^ x[9];
  assign t[16] = t[21] ^ x[12];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = t[23] ^ x[18];
  assign t[19] = (x[4] & x[5]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = ~(t[11] & t[14]);
  assign t[8] = ~x[2] & t[15];
  assign t[9] = ~(t[16]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind106(x, y);
 input [18:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[12] | t[9]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[18] ^ x[6];
  assign t[14] = t[19] ^ x[9];
  assign t[15] = t[20] ^ x[12];
  assign t[16] = t[21] ^ x[15];
  assign t[17] = t[22] ^ x[18];
  assign t[18] = (x[4] & x[5]);
  assign t[19] = (x[7] & x[8]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = (x[10] & x[11]);
  assign t[21] = (x[13] & x[14]);
  assign t[22] = (x[16] & x[17]);
  assign t[2] = x[2] ? x[3] : t[4];
  assign t[3] = ~(t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] & t[10]);
  assign t[7] = t[11] | t[13];
  assign t[8] = ~x[2] & t[14];
  assign t[9] = ~(t[15]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind107(x, y);
 input [31:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[26] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[27] | t[20]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[16];
  assign t[29] = t[38] ^ x[19];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[25];
  assign t[32] = t[41] ^ x[28];
  assign t[33] = t[42] ^ x[31];
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[8] & x[9]);
  assign t[36] = (x[11] & x[12]);
  assign t[37] = (x[14] & x[15]);
  assign t[38] = (x[17] & x[18]);
  assign t[39] = (x[20] & x[21]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[23] & x[24]);
  assign t[41] = (x[26] & x[27]);
  assign t[42] = (x[29] & x[30]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind108(x, y);
 input [25:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[21] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[24] & t[17]);
  assign t[15] = ~(t[25]);
  assign t[16] = ~(t[25] & t[18]);
  assign t[17] = ~(t[20]);
  assign t[18] = ~(t[22]);
  assign t[19] = t[26] ^ x[5];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = t[27] ^ x[10];
  assign t[21] = t[28] ^ x[13];
  assign t[22] = t[29] ^ x[16];
  assign t[23] = t[30] ^ x[19];
  assign t[24] = t[31] ^ x[22];
  assign t[25] = t[32] ^ x[25];
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[8] & x[9]);
  assign t[28] = (x[11] & x[12]);
  assign t[29] = (x[14] & x[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[17] & x[18]);
  assign t[31] = (x[20] & x[21]);
  assign t[32] = (x[23] & x[24]);
  assign t[3] = ~x[2] & t[19];
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[6] : t[7];
  assign t[6] = x[2] ? x[7] : t[8];
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[20] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind109(x, y);
 input [31:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[26]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[29] & t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[31] & t[30]);
  assign t[24] = ~(t[33]);
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[16];
  assign t[29] = t[38] ^ x[19];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[25];
  assign t[32] = t[41] ^ x[28];
  assign t[33] = t[42] ^ x[31];
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[8] & x[9]);
  assign t[36] = (x[11] & x[12]);
  assign t[37] = (x[14] & x[15]);
  assign t[38] = (x[17] & x[18]);
  assign t[39] = (x[20] & x[21]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[23] & x[24]);
  assign t[41] = (x[26] & x[27]);
  assign t[42] = (x[29] & x[30]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind110(x, y);
 input [31:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = t[17] | t[24];
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = t[20] | t[25];
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[21] | t[15]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[29]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[22] | t[18]);
  assign t[21] = ~(t[30]);
  assign t[22] = ~(t[31]);
  assign t[23] = t[32] ^ x[7];
  assign t[24] = t[33] ^ x[10];
  assign t[25] = t[34] ^ x[13];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[22];
  assign t[29] = t[38] ^ x[25];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[28];
  assign t[31] = t[40] ^ x[31];
  assign t[32] = (x[5] & x[6]);
  assign t[33] = (x[8] & x[9]);
  assign t[34] = (x[11] & x[12]);
  assign t[35] = (x[14] & x[15]);
  assign t[36] = (x[17] & x[18]);
  assign t[37] = (x[20] & x[21]);
  assign t[38] = (x[23] & x[24]);
  assign t[39] = (x[26] & x[27]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[29] & x[30]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[23];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind111(x, y);
 input [31:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[24] | t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[25] | t[18]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[27]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[30]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = t[32] ^ x[5];
  assign t[24] = t[33] ^ x[10];
  assign t[25] = t[34] ^ x[13];
  assign t[26] = t[35] ^ x[16];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[22];
  assign t[29] = t[38] ^ x[25];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[28];
  assign t[31] = t[40] ^ x[31];
  assign t[32] = (x[3] & x[4]);
  assign t[33] = (x[8] & x[9]);
  assign t[34] = (x[11] & x[12]);
  assign t[35] = (x[14] & x[15]);
  assign t[36] = (x[17] & x[18]);
  assign t[37] = (x[20] & x[21]);
  assign t[38] = (x[23] & x[24]);
  assign t[39] = (x[26] & x[27]);
  assign t[3] = ~x[2] & t[23];
  assign t[40] = (x[29] & x[30]);
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[6] : t[7];
  assign t[6] = x[2] ? x[7] : t[8];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13] | t[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind112(x, y);
 input [25:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25] & t[18]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[26] & t[19]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[27] & t[20]);
  assign t[19] = ~(t[22]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[24]);
  assign t[21] = t[28] ^ x[7];
  assign t[22] = t[29] ^ x[10];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[16];
  assign t[25] = t[32] ^ x[19];
  assign t[26] = t[33] ^ x[22];
  assign t[27] = t[34] ^ x[25];
  assign t[28] = (x[5] & x[6]);
  assign t[29] = (x[8] & x[9]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[11] & x[12]);
  assign t[31] = (x[14] & x[15]);
  assign t[32] = (x[17] & x[18]);
  assign t[33] = (x[20] & x[21]);
  assign t[34] = (x[23] & x[24]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[21];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind113(x, y);
 input [31:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[26]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[29] & t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[31] & t[30]);
  assign t[24] = ~(t[33]);
  assign t[25] = t[34] ^ x[7];
  assign t[26] = t[35] ^ x[10];
  assign t[27] = t[36] ^ x[13];
  assign t[28] = t[37] ^ x[16];
  assign t[29] = t[38] ^ x[19];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[25];
  assign t[32] = t[41] ^ x[28];
  assign t[33] = t[42] ^ x[31];
  assign t[34] = (x[5] & x[6]);
  assign t[35] = (x[8] & x[9]);
  assign t[36] = (x[11] & x[12]);
  assign t[37] = (x[14] & x[15]);
  assign t[38] = (x[17] & x[18]);
  assign t[39] = (x[20] & x[21]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[23] & x[24]);
  assign t[41] = (x[26] & x[27]);
  assign t[42] = (x[29] & x[30]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~x[2] & t[25];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind114(x, y);
 input [31:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~t[2];
  assign t[10] = t[15] | t[22];
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = t[18] | t[23];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[19] | t[13]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[20] | t[16]);
  assign t[19] = ~(t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[29]);
  assign t[21] = t[30] ^ x[5];
  assign t[22] = t[31] ^ x[10];
  assign t[23] = t[32] ^ x[13];
  assign t[24] = t[33] ^ x[16];
  assign t[25] = t[34] ^ x[19];
  assign t[26] = t[35] ^ x[22];
  assign t[27] = t[36] ^ x[25];
  assign t[28] = t[37] ^ x[28];
  assign t[29] = t[38] ^ x[31];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (x[3] & x[4]);
  assign t[31] = (x[8] & x[9]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[3] = ~x[2] & t[21];
  assign t[4] = ~t[6];
  assign t[5] = x[2] ? x[6] : t[7];
  assign t[6] = x[2] ? x[7] : t[8];
  assign t[7] = ~(t[9] & t[10]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind115(x, y);
 input [34:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[28] | t[19]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[30] | t[22]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[19];
  assign t[32] = t[42] ^ x[22];
  assign t[33] = t[43] ^ x[25];
  assign t[34] = t[44] ^ x[28];
  assign t[35] = t[45] ^ x[31];
  assign t[36] = t[46] ^ x[34];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[43] = (x[23] & x[24]);
  assign t[44] = (x[26] & x[27]);
  assign t[45] = (x[29] & x[30]);
  assign t[46] = (x[32] & x[33]);
  assign t[4] = ~(~x[2] & ~t[27]);
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind116(x, y);
 input [28:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[24] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[27] & t[19]);
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[29] & t[21]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[30] & t[22]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[27]);
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[10];
  assign t[25] = t[33] ^ x[13];
  assign t[26] = t[34] ^ x[16];
  assign t[27] = t[35] ^ x[19];
  assign t[28] = t[36] ^ x[22];
  assign t[29] = t[37] ^ x[25];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[38] ^ x[28];
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[8] & x[9]);
  assign t[33] = (x[11] & x[12]);
  assign t[34] = (x[14] & x[15]);
  assign t[35] = (x[17] & x[18]);
  assign t[36] = (x[20] & x[21]);
  assign t[37] = (x[23] & x[24]);
  assign t[38] = (x[26] & x[27]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[4] = ~x[2] & t[23];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind117(x, y);
 input [34:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[28]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[30]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[32] & t[31]);
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[34] & t[33]);
  assign t[26] = ~(t[36]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[19];
  assign t[32] = t[42] ^ x[22];
  assign t[33] = t[43] ^ x[25];
  assign t[34] = t[44] ^ x[28];
  assign t[35] = t[45] ^ x[31];
  assign t[36] = t[46] ^ x[34];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[43] = (x[23] & x[24]);
  assign t[44] = (x[26] & x[27]);
  assign t[45] = (x[29] & x[30]);
  assign t[46] = (x[32] & x[33]);
  assign t[4] = ~x[2] & t[27];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind118(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = t[18] | t[24];
  assign t[13] = ~x[2] & t[25];
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = t[21] | t[26];
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[22] | t[16]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[23] | t[19]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[32]);
  assign t[24] = t[33] ^ x[7];
  assign t[25] = t[34] ^ x[10];
  assign t[26] = t[35] ^ x[13];
  assign t[27] = t[36] ^ x[16];
  assign t[28] = t[37] ^ x[19];
  assign t[29] = t[38] ^ x[22];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[39] ^ x[25];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[5] & x[6]);
  assign t[34] = (x[8] & x[9]);
  assign t[35] = (x[11] & x[12]);
  assign t[36] = (x[14] & x[15]);
  assign t[37] = (x[17] & x[18]);
  assign t[38] = (x[20] & x[21]);
  assign t[39] = (x[23] & x[24]);
  assign t[3] = t[6] ? x[1] : x[0];
  assign t[40] = (x[26] & x[27]);
  assign t[41] = (x[29] & x[30]);
  assign t[4] = ~t[7];
  assign t[5] = x[2] ? x[3] : t[8];
  assign t[6] = ~(t[9]);
  assign t[7] = x[2] ? x[4] : t[10];
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind119(x, y);
 input [34:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[28] | t[19]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[30] | t[22]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[35]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[19];
  assign t[32] = t[42] ^ x[22];
  assign t[33] = t[43] ^ x[25];
  assign t[34] = t[44] ^ x[28];
  assign t[35] = t[45] ^ x[31];
  assign t[36] = t[46] ^ x[34];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[43] = (x[23] & x[24]);
  assign t[44] = (x[26] & x[27]);
  assign t[45] = (x[29] & x[30]);
  assign t[46] = (x[32] & x[33]);
  assign t[4] = ~(~x[2] & ~t[27]);
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind120(x, y);
 input [28:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[24] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[27] & t[19]);
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[29] & t[21]);
  assign t[19] = ~(t[30]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[30] & t[22]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[27]);
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[10];
  assign t[25] = t[33] ^ x[13];
  assign t[26] = t[34] ^ x[16];
  assign t[27] = t[35] ^ x[19];
  assign t[28] = t[36] ^ x[22];
  assign t[29] = t[37] ^ x[25];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[38] ^ x[28];
  assign t[31] = (x[3] & x[4]);
  assign t[32] = (x[8] & x[9]);
  assign t[33] = (x[11] & x[12]);
  assign t[34] = (x[14] & x[15]);
  assign t[35] = (x[17] & x[18]);
  assign t[36] = (x[20] & x[21]);
  assign t[37] = (x[23] & x[24]);
  assign t[38] = (x[26] & x[27]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[4] = ~x[2] & t[23];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind121(x, y);
 input [34:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[28]);
  assign t[14] = ~x[2] & t[29];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[22] & t[30]);
  assign t[17] = ~(t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[23] & t[24]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[32] & t[31]);
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[34] & t[33]);
  assign t[26] = ~(t[36]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[10];
  assign t[29] = t[39] ^ x[13];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[16];
  assign t[31] = t[41] ^ x[19];
  assign t[32] = t[42] ^ x[22];
  assign t[33] = t[43] ^ x[25];
  assign t[34] = t[44] ^ x[28];
  assign t[35] = t[45] ^ x[31];
  assign t[36] = t[46] ^ x[34];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[8] & x[9]);
  assign t[39] = (x[11] & x[12]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[14] & x[15]);
  assign t[41] = (x[17] & x[18]);
  assign t[42] = (x[20] & x[21]);
  assign t[43] = (x[23] & x[24]);
  assign t[44] = (x[26] & x[27]);
  assign t[45] = (x[29] & x[30]);
  assign t[46] = (x[32] & x[33]);
  assign t[4] = ~x[2] & t[27];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind122(x, y);
 input [34:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[2];
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[26];
  assign t[14] = ~x[2] & t[27];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = t[22] | t[28];
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[23] | t[17]);
  assign t[1] = ~(t[3] ^ t[4]);
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[24] | t[20]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[34]);
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[10];
  assign t[27] = t[37] ^ x[13];
  assign t[28] = t[38] ^ x[16];
  assign t[29] = t[39] ^ x[19];
  assign t[2] = ~(t[5] ^ t[6]);
  assign t[30] = t[40] ^ x[22];
  assign t[31] = t[41] ^ x[25];
  assign t[32] = t[42] ^ x[28];
  assign t[33] = t[43] ^ x[31];
  assign t[34] = t[44] ^ x[34];
  assign t[35] = (x[3] & x[4]);
  assign t[36] = (x[8] & x[9]);
  assign t[37] = (x[11] & x[12]);
  assign t[38] = (x[14] & x[15]);
  assign t[39] = (x[17] & x[18]);
  assign t[3] = t[7] ? x[1] : x[0];
  assign t[40] = (x[20] & x[21]);
  assign t[41] = (x[23] & x[24]);
  assign t[42] = (x[26] & x[27]);
  assign t[43] = (x[29] & x[30]);
  assign t[44] = (x[32] & x[33]);
  assign t[4] = ~x[2] & t[25];
  assign t[5] = ~t[8];
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind123(x, y);
 input [44:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[20];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[23];
  assign t[41] = t[54] ^ x[26];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[32];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = t[58] ^ x[38];
  assign t[46] = t[59] ^ x[41];
  assign t[47] = t[60] ^ x[44];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[18] & x[19]);
  assign t[53] = (x[21] & x[22]);
  assign t[54] = (x[24] & x[25]);
  assign t[55] = (x[27] & x[28]);
  assign t[56] = (x[30] & x[31]);
  assign t[57] = (x[33] & x[34]);
  assign t[58] = (x[36] & x[37]);
  assign t[59] = (x[39] & x[40]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[42] & x[43]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind124(x, y);
 input [35:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = t[47] ^ x[32];
  assign t[38] = t[48] ^ x[35];
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[12] & x[13]);
  assign t[42] = (x[15] & x[16]);
  assign t[43] = (x[18] & x[19]);
  assign t[44] = (x[21] & x[22]);
  assign t[45] = (x[24] & x[25]);
  assign t[46] = (x[27] & x[28]);
  assign t[47] = (x[30] & x[31]);
  assign t[48] = (x[33] & x[34]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind125(x, y);
 input [44:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = ~(t[22] & t[36]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[37]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] & t[34]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[44] & t[43]);
  assign t[34] = ~(t[47]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[20];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[23];
  assign t[41] = t[54] ^ x[26];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[32];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = t[58] ^ x[38];
  assign t[46] = t[59] ^ x[41];
  assign t[47] = t[60] ^ x[44];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[18] & x[19]);
  assign t[53] = (x[21] & x[22]);
  assign t[54] = (x[24] & x[25]);
  assign t[55] = (x[27] & x[28]);
  assign t[56] = (x[30] & x[31]);
  assign t[57] = (x[33] & x[34]);
  assign t[58] = (x[36] & x[37]);
  assign t[59] = (x[39] & x[40]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[42] & x[43]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind126(x, y);
 input [44:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[8];
  assign t[33] = t[46] ^ x[11];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[20];
  assign t[37] = t[50] ^ x[23];
  assign t[38] = t[51] ^ x[26];
  assign t[39] = t[52] ^ x[29];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[32];
  assign t[41] = t[54] ^ x[35];
  assign t[42] = t[55] ^ x[38];
  assign t[43] = t[56] ^ x[41];
  assign t[44] = t[57] ^ x[44];
  assign t[45] = (x[6] & x[7]);
  assign t[46] = (x[9] & x[10]);
  assign t[47] = (x[12] & x[13]);
  assign t[48] = (x[15] & x[16]);
  assign t[49] = (x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[21] & x[22]);
  assign t[51] = (x[24] & x[25]);
  assign t[52] = (x[27] & x[28]);
  assign t[53] = (x[30] & x[31]);
  assign t[54] = (x[33] & x[34]);
  assign t[55] = (x[36] & x[37]);
  assign t[56] = (x[39] & x[40]);
  assign t[57] = (x[42] & x[43]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind127(x, y);
 input [44:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[20];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[23];
  assign t[41] = t[54] ^ x[26];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[32];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = t[58] ^ x[38];
  assign t[46] = t[59] ^ x[41];
  assign t[47] = t[60] ^ x[44];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[18] & x[19]);
  assign t[53] = (x[21] & x[22]);
  assign t[54] = (x[24] & x[25]);
  assign t[55] = (x[27] & x[28]);
  assign t[56] = (x[30] & x[31]);
  assign t[57] = (x[33] & x[34]);
  assign t[58] = (x[36] & x[37]);
  assign t[59] = (x[39] & x[40]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[42] & x[43]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind128(x, y);
 input [35:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[28] & t[18]);
  assign t[13] = ~(t[29] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[34] & t[24]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[35]);
  assign t[21] = ~(t[35] & t[25]);
  assign t[22] = ~(t[36]);
  assign t[23] = ~(t[36] & t[26]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[30]);
  assign t[26] = ~(t[32]);
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[11];
  assign t[29] = t[39] ^ x[14];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[17];
  assign t[31] = t[41] ^ x[20];
  assign t[32] = t[42] ^ x[23];
  assign t[33] = t[43] ^ x[26];
  assign t[34] = t[44] ^ x[29];
  assign t[35] = t[45] ^ x[32];
  assign t[36] = t[46] ^ x[35];
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[9] & x[10]);
  assign t[39] = (x[12] & x[13]);
  assign t[3] = ~x[2] & t[27];
  assign t[40] = (x[15] & x[16]);
  assign t[41] = (x[18] & x[19]);
  assign t[42] = (x[21] & x[22]);
  assign t[43] = (x[24] & x[25]);
  assign t[44] = (x[27] & x[28]);
  assign t[45] = (x[30] & x[31]);
  assign t[46] = (x[33] & x[34]);
  assign t[4] = t[6];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind129(x, y);
 input [44:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = ~(t[20] & t[34]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = ~(t[23] & t[35]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26] & t[36]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] & t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] & t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[38] & t[37]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[45]);
  assign t[33] = t[46] ^ x[5];
  assign t[34] = t[47] ^ x[11];
  assign t[35] = t[48] ^ x[14];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[20];
  assign t[38] = t[51] ^ x[23];
  assign t[39] = t[52] ^ x[26];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[29];
  assign t[41] = t[54] ^ x[32];
  assign t[42] = t[55] ^ x[35];
  assign t[43] = t[56] ^ x[38];
  assign t[44] = t[57] ^ x[41];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = (x[3] & x[4]);
  assign t[47] = (x[9] & x[10]);
  assign t[48] = (x[12] & x[13]);
  assign t[49] = (x[15] & x[16]);
  assign t[4] = t[6];
  assign t[50] = (x[18] & x[19]);
  assign t[51] = (x[21] & x[22]);
  assign t[52] = (x[24] & x[25]);
  assign t[53] = (x[27] & x[28]);
  assign t[54] = (x[30] & x[31]);
  assign t[55] = (x[33] & x[34]);
  assign t[56] = (x[36] & x[37]);
  assign t[57] = (x[39] & x[40]);
  assign t[58] = (x[42] & x[43]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind130(x, y);
 input [44:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[8];
  assign t[33] = t[46] ^ x[11];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[20];
  assign t[37] = t[50] ^ x[23];
  assign t[38] = t[51] ^ x[26];
  assign t[39] = t[52] ^ x[29];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[32];
  assign t[41] = t[54] ^ x[35];
  assign t[42] = t[55] ^ x[38];
  assign t[43] = t[56] ^ x[41];
  assign t[44] = t[57] ^ x[44];
  assign t[45] = (x[6] & x[7]);
  assign t[46] = (x[9] & x[10]);
  assign t[47] = (x[12] & x[13]);
  assign t[48] = (x[15] & x[16]);
  assign t[49] = (x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[21] & x[22]);
  assign t[51] = (x[24] & x[25]);
  assign t[52] = (x[27] & x[28]);
  assign t[53] = (x[30] & x[31]);
  assign t[54] = (x[33] & x[34]);
  assign t[55] = (x[36] & x[37]);
  assign t[56] = (x[39] & x[40]);
  assign t[57] = (x[42] & x[43]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind131(x, y);
 input [44:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[18] | t[19]);
  assign t[13] = ~(t[34] | t[20]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[15] = ~(t[35] | t[23]);
  assign t[16] = ~(t[24] | t[25]);
  assign t[17] = ~(t[36] | t[26]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] | t[32]);
  assign t[27] = ~(t[43]);
  assign t[28] = ~(t[37] | t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = t[46] ^ x[5];
  assign t[34] = t[47] ^ x[11];
  assign t[35] = t[48] ^ x[14];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[20];
  assign t[38] = t[51] ^ x[23];
  assign t[39] = t[52] ^ x[26];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[29];
  assign t[41] = t[54] ^ x[32];
  assign t[42] = t[55] ^ x[35];
  assign t[43] = t[56] ^ x[38];
  assign t[44] = t[57] ^ x[41];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = (x[3] & x[4]);
  assign t[47] = (x[9] & x[10]);
  assign t[48] = (x[12] & x[13]);
  assign t[49] = (x[15] & x[16]);
  assign t[4] = t[6];
  assign t[50] = (x[18] & x[19]);
  assign t[51] = (x[21] & x[22]);
  assign t[52] = (x[24] & x[25]);
  assign t[53] = (x[27] & x[28]);
  assign t[54] = (x[30] & x[31]);
  assign t[55] = (x[33] & x[34]);
  assign t[56] = (x[36] & x[37]);
  assign t[57] = (x[39] & x[40]);
  assign t[58] = (x[42] & x[43]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind132(x, y);
 input [35:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = t[47] ^ x[32];
  assign t[38] = t[48] ^ x[35];
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[12] & x[13]);
  assign t[42] = (x[15] & x[16]);
  assign t[43] = (x[18] & x[19]);
  assign t[44] = (x[21] & x[22]);
  assign t[45] = (x[24] & x[25]);
  assign t[46] = (x[27] & x[28]);
  assign t[47] = (x[30] & x[31]);
  assign t[48] = (x[33] & x[34]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind133(x, y);
 input [44:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = ~(t[22] & t[36]);
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = ~(t[25] & t[37]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] & t[34]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[44] & t[43]);
  assign t[34] = ~(t[47]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[20];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[23];
  assign t[41] = t[54] ^ x[26];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[32];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = t[58] ^ x[38];
  assign t[46] = t[59] ^ x[41];
  assign t[47] = t[60] ^ x[44];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[18] & x[19]);
  assign t[53] = (x[21] & x[22]);
  assign t[54] = (x[24] & x[25]);
  assign t[55] = (x[27] & x[28]);
  assign t[56] = (x[30] & x[31]);
  assign t[57] = (x[33] & x[34]);
  assign t[58] = (x[36] & x[37]);
  assign t[59] = (x[39] & x[40]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[42] & x[43]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind134(x, y);
 input [44:0] x;
 output y;

 wire [55:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = t[20] | t[31];
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = t[23] | t[32];
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = t[26] | t[33];
  assign t[18] = ~(t[34]);
  assign t[19] = ~(t[35]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] | t[18]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[28] | t[21]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[29] | t[24]);
  assign t[27] = ~(t[40]);
  assign t[28] = ~(t[41]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ x[5];
  assign t[31] = t[44] ^ x[11];
  assign t[32] = t[45] ^ x[14];
  assign t[33] = t[46] ^ x[17];
  assign t[34] = t[47] ^ x[20];
  assign t[35] = t[48] ^ x[23];
  assign t[36] = t[49] ^ x[26];
  assign t[37] = t[50] ^ x[29];
  assign t[38] = t[51] ^ x[32];
  assign t[39] = t[52] ^ x[35];
  assign t[3] = ~x[2] & t[30];
  assign t[40] = t[53] ^ x[38];
  assign t[41] = t[54] ^ x[41];
  assign t[42] = t[55] ^ x[44];
  assign t[43] = (x[3] & x[4]);
  assign t[44] = (x[9] & x[10]);
  assign t[45] = (x[12] & x[13]);
  assign t[46] = (x[15] & x[16]);
  assign t[47] = (x[18] & x[19]);
  assign t[48] = (x[21] & x[22]);
  assign t[49] = (x[24] & x[25]);
  assign t[4] = t[6];
  assign t[50] = (x[27] & x[28]);
  assign t[51] = (x[30] & x[31]);
  assign t[52] = (x[33] & x[34]);
  assign t[53] = (x[36] & x[37]);
  assign t[54] = (x[39] & x[40]);
  assign t[55] = (x[42] & x[43]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind135(x, y);
 input [44:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[35];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[36] | t[22]);
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = ~(t[37] | t[25]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[19] = ~(t[38] | t[28]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[29] | t[30]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[39] | t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[41] | t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[43] | t[44]);
  assign t[35] = t[48] ^ x[8];
  assign t[36] = t[49] ^ x[11];
  assign t[37] = t[50] ^ x[14];
  assign t[38] = t[51] ^ x[17];
  assign t[39] = t[52] ^ x[20];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[23];
  assign t[41] = t[54] ^ x[26];
  assign t[42] = t[55] ^ x[29];
  assign t[43] = t[56] ^ x[32];
  assign t[44] = t[57] ^ x[35];
  assign t[45] = t[58] ^ x[38];
  assign t[46] = t[59] ^ x[41];
  assign t[47] = t[60] ^ x[44];
  assign t[48] = (x[6] & x[7]);
  assign t[49] = (x[9] & x[10]);
  assign t[4] = t[7];
  assign t[50] = (x[12] & x[13]);
  assign t[51] = (x[15] & x[16]);
  assign t[52] = (x[18] & x[19]);
  assign t[53] = (x[21] & x[22]);
  assign t[54] = (x[24] & x[25]);
  assign t[55] = (x[27] & x[28]);
  assign t[56] = (x[30] & x[31]);
  assign t[57] = (x[33] & x[34]);
  assign t[58] = (x[36] & x[37]);
  assign t[59] = (x[39] & x[40]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = (x[42] & x[43]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind136(x, y);
 input [35:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[29];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[36] & t[26]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[37] & t[27]);
  assign t[24] = ~(t[38]);
  assign t[25] = ~(t[38] & t[28]);
  assign t[26] = ~(t[30]);
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[34]);
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = t[47] ^ x[32];
  assign t[38] = t[48] ^ x[35];
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[12] & x[13]);
  assign t[42] = (x[15] & x[16]);
  assign t[43] = (x[18] & x[19]);
  assign t[44] = (x[21] & x[22]);
  assign t[45] = (x[24] & x[25]);
  assign t[46] = (x[27] & x[28]);
  assign t[47] = (x[30] & x[31]);
  assign t[48] = (x[33] & x[34]);
  assign t[4] = t[7];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind137(x, y);
 input [44:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[18] & t[19]);
  assign t[13] = ~(t[20] & t[34]);
  assign t[14] = ~(t[21] & t[22]);
  assign t[15] = ~(t[23] & t[35]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(t[26] & t[36]);
  assign t[18] = ~(t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[27] & t[28]);
  assign t[21] = ~(t[39]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[29] & t[30]);
  assign t[24] = ~(t[41]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[38] & t[37]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[40] & t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[44]);
  assign t[31] = ~(t[42] & t[41]);
  assign t[32] = ~(t[45]);
  assign t[33] = t[46] ^ x[5];
  assign t[34] = t[47] ^ x[11];
  assign t[35] = t[48] ^ x[14];
  assign t[36] = t[49] ^ x[17];
  assign t[37] = t[50] ^ x[20];
  assign t[38] = t[51] ^ x[23];
  assign t[39] = t[52] ^ x[26];
  assign t[3] = ~x[2] & t[33];
  assign t[40] = t[53] ^ x[29];
  assign t[41] = t[54] ^ x[32];
  assign t[42] = t[55] ^ x[35];
  assign t[43] = t[56] ^ x[38];
  assign t[44] = t[57] ^ x[41];
  assign t[45] = t[58] ^ x[44];
  assign t[46] = (x[3] & x[4]);
  assign t[47] = (x[9] & x[10]);
  assign t[48] = (x[12] & x[13]);
  assign t[49] = (x[15] & x[16]);
  assign t[4] = t[6];
  assign t[50] = (x[18] & x[19]);
  assign t[51] = (x[21] & x[22]);
  assign t[52] = (x[24] & x[25]);
  assign t[53] = (x[27] & x[28]);
  assign t[54] = (x[30] & x[31]);
  assign t[55] = (x[33] & x[34]);
  assign t[56] = (x[36] & x[37]);
  assign t[57] = (x[39] & x[40]);
  assign t[58] = (x[42] & x[43]);
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[6] = x[2] ? x[6] : t[9];
  assign t[7] = x[2] ? x[7] : t[10];
  assign t[8] = x[2] ? x[8] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1ind138(x, y);
 input [44:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~t[2];
  assign t[10] = ~x[2] & t[32];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[21]);
  assign t[15] = t[22] | t[33];
  assign t[16] = ~(t[23] & t[24]);
  assign t[17] = t[25] | t[34];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[35];
  assign t[1] = t[3] ? x[1] : x[0];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[29] | t[20]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[30] | t[23]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[31] | t[26]);
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = t[45] ^ x[8];
  assign t[33] = t[46] ^ x[11];
  assign t[34] = t[47] ^ x[14];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[20];
  assign t[37] = t[50] ^ x[23];
  assign t[38] = t[51] ^ x[26];
  assign t[39] = t[52] ^ x[29];
  assign t[3] = ~(t[6]);
  assign t[40] = t[53] ^ x[32];
  assign t[41] = t[54] ^ x[35];
  assign t[42] = t[55] ^ x[38];
  assign t[43] = t[56] ^ x[41];
  assign t[44] = t[57] ^ x[44];
  assign t[45] = (x[6] & x[7]);
  assign t[46] = (x[9] & x[10]);
  assign t[47] = (x[12] & x[13]);
  assign t[48] = (x[15] & x[16]);
  assign t[49] = (x[18] & x[19]);
  assign t[4] = t[7];
  assign t[50] = (x[21] & x[22]);
  assign t[51] = (x[24] & x[25]);
  assign t[52] = (x[27] & x[28]);
  assign t[53] = (x[30] & x[31]);
  assign t[54] = (x[33] & x[34]);
  assign t[55] = (x[36] & x[37]);
  assign t[56] = (x[39] & x[40]);
  assign t[57] = (x[42] & x[43]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = x[2] ? x[3] : t[11];
  assign t[8] = x[2] ? x[4] : t[12];
  assign t[9] = x[2] ? x[5] : t[13];
  assign y = ~(t[0] ^ t[1]);
endmodule

module R1_ind(x, y);
 input [414:0] x;
 output [138:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[8], x[7], x[6]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[11], x[10], x[9]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[14], x[13], x[12]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[17], x[16], x[15]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[20], x[19], x[18]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[23], x[22], x[21]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[26], x[25], x[24]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[29], x[28], x[27]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[35], x[34], x[33]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[38], x[37], x[36]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[41], x[40], x[39]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[44], x[43], x[42]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[47], x[46], x[45]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[50], x[49], x[48]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[53], x[52], x[51]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[56], x[55], x[54]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[59], x[58], x[57]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[61], x[60]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[68], x[67], x[66]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[71], x[70], x[69]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[74], x[73], x[72]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[77], x[76], x[75]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[80], x[79], x[78]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[82], x[81]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[86], x[85], x[84]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[89], x[88], x[87]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[92], x[91], x[90]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[95], x[94], x[93]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[98], x[97], x[96]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[101], x[100], x[99]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[103], x[102]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[107], x[106], x[105]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[110], x[109], x[108]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[113], x[112], x[111]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[116], x[115], x[114]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[119], x[118], x[117]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[122], x[121], x[120]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[128], x[127], x[126]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[131], x[130], x[129]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[134], x[133], x[132]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[137], x[136], x[135]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[140], x[139], x[138]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[143], x[142], x[141]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[146], x[145], x[144]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[149], x[148], x[147]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[152], x[151], x[150]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[155], x[154], x[153]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[158], x[157], x[156]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[161], x[160], x[159]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[164], x[163], x[162]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[167], x[166], x[165]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[170], x[169], x[168]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[173], x[172], x[171]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[176], x[175], x[174]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[179], x[178], x[177]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[182], x[181], x[180]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[185], x[184], x[183]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[188], x[187], x[186]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[191], x[190], x[189]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[194], x[193], x[192]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[219], x[218], x[217], x[195]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[219], x[218], x[217], x[222], x[221], x[220], x[195]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[207], x[206], x[205], x[195]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[204], x[203], x[202], x[195]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[201], x[200], x[199], x[207], x[206], x[205], x[195]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[213], x[212], x[211], x[195]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[216], x[215], x[214], x[195]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[198], x[197], x[196], x[195]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[213], x[212], x[211], x[210], x[209], x[208], x[195]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[185], x[184], x[183], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[219], x[218], x[217], x[225], x[195], x[224], x[223]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[194], x[193], x[192], x[219], x[218], x[217], x[185], x[184], x[183], x[191], x[190], x[189], x[228], x[195], x[227], x[226]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[191], x[190], x[189], x[185], x[184], x[183], x[194], x[193], x[192], x[188], x[187], x[186], x[219], x[218], x[217], x[231], x[195], x[230], x[229]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[191], x[190], x[189], x[185], x[184], x[183], x[194], x[193], x[192], x[219], x[218], x[217], x[188], x[187], x[186], x[234], x[195], x[233], x[232]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[149], x[148], x[147], x[158], x[157], x[156], x[155], x[154], x[153], x[219], x[218], x[217], x[152], x[151], x[150], x[237], x[195], x[236], x[235]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[158], x[157], x[156], x[219], x[218], x[217], x[149], x[148], x[147], x[155], x[154], x[153], x[240], x[195], x[239], x[238]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[155], x[154], x[153], x[149], x[148], x[147], x[158], x[157], x[156], x[219], x[218], x[217], x[152], x[151], x[150], x[243], x[195], x[242], x[241]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[155], x[154], x[153], x[149], x[148], x[147], x[158], x[157], x[156], x[219], x[218], x[217], x[152], x[151], x[150], x[246], x[195], x[245], x[244]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[161], x[160], x[159], x[170], x[169], x[168], x[167], x[166], x[165], x[219], x[218], x[217], x[164], x[163], x[162], x[249], x[195], x[248], x[247]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[170], x[169], x[168], x[219], x[218], x[217], x[161], x[160], x[159], x[167], x[166], x[165], x[252], x[195], x[251], x[250]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[167], x[166], x[165], x[161], x[160], x[159], x[170], x[169], x[168], x[219], x[218], x[217], x[164], x[163], x[162], x[255], x[195], x[254], x[253]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[167], x[166], x[165], x[161], x[160], x[159], x[170], x[169], x[168], x[219], x[218], x[217], x[164], x[163], x[162], x[258], x[195], x[257], x[256]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[173], x[172], x[171], x[182], x[181], x[180], x[179], x[178], x[177], x[219], x[218], x[217], x[176], x[175], x[174], x[261], x[195], x[260], x[259]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[182], x[181], x[180], x[219], x[218], x[217], x[173], x[172], x[171], x[179], x[178], x[177], x[264], x[195], x[263], x[262]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[179], x[178], x[177], x[173], x[172], x[171], x[182], x[181], x[180], x[219], x[218], x[217], x[176], x[175], x[174], x[267], x[195], x[266], x[265]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[179], x[178], x[177], x[173], x[172], x[171], x[182], x[181], x[180], x[219], x[218], x[217], x[176], x[175], x[174], x[270], x[195], x[269], x[268]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[101], x[100], x[99], x[110], x[109], x[108], x[107], x[106], x[105], x[219], x[218], x[217], x[104], x[103], x[102], x[273], x[195], x[272], x[271]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[110], x[109], x[108], x[219], x[218], x[217], x[101], x[100], x[99], x[107], x[106], x[105], x[276], x[195], x[275], x[274]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[107], x[106], x[105], x[101], x[100], x[99], x[110], x[109], x[108], x[219], x[218], x[217], x[104], x[103], x[102], x[279], x[195], x[278], x[277]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[107], x[106], x[105], x[101], x[100], x[99], x[110], x[109], x[108], x[219], x[218], x[217], x[104], x[103], x[102], x[282], x[195], x[281], x[280]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[137], x[136], x[135], x[146], x[145], x[144], x[143], x[142], x[141], x[219], x[218], x[217], x[140], x[139], x[138], x[285], x[195], x[284], x[283]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[146], x[145], x[144], x[219], x[218], x[217], x[137], x[136], x[135], x[143], x[142], x[141], x[288], x[195], x[287], x[286]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[143], x[142], x[141], x[137], x[136], x[135], x[146], x[145], x[144], x[140], x[139], x[138], x[219], x[218], x[217], x[291], x[195], x[290], x[289]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[143], x[142], x[141], x[137], x[136], x[135], x[146], x[145], x[144], x[140], x[139], x[138], x[219], x[218], x[217], x[294], x[195], x[293], x[292]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[125], x[124], x[123], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[219], x[218], x[217], x[297], x[195], x[296], x[295]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[134], x[133], x[132], x[125], x[124], x[123], x[131], x[130], x[129], x[219], x[218], x[217], x[300], x[195], x[299], x[298]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[131], x[130], x[129], x[125], x[124], x[123], x[134], x[133], x[132], x[128], x[127], x[126], x[219], x[218], x[217], x[303], x[195], x[302], x[301]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[131], x[130], x[129], x[125], x[124], x[123], x[134], x[133], x[132], x[128], x[127], x[126], x[219], x[218], x[217], x[306], x[195], x[305], x[304]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[113], x[112], x[111], x[122], x[121], x[120], x[119], x[118], x[117], x[219], x[218], x[217], x[116], x[115], x[114], x[309], x[195], x[308], x[307]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[122], x[121], x[120], x[219], x[218], x[217], x[113], x[112], x[111], x[119], x[118], x[117], x[312], x[195], x[311], x[310]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[119], x[118], x[117], x[113], x[112], x[111], x[122], x[121], x[120], x[219], x[218], x[217], x[116], x[115], x[114], x[315], x[195], x[314], x[313]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[119], x[118], x[117], x[113], x[112], x[111], x[122], x[121], x[120], x[219], x[218], x[217], x[116], x[115], x[114], x[318], x[195], x[317], x[316]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[53], x[52], x[51], x[185], x[184], x[183], x[62], x[61], x[60], x[59], x[58], x[57], x[194], x[193], x[192], x[191], x[190], x[189], x[56], x[55], x[54], x[188], x[187], x[186], x[219], x[218], x[217], x[321], x[225], x[195], x[320], x[319]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[62], x[61], x[60], x[194], x[193], x[192], x[53], x[52], x[51], x[59], x[58], x[57], x[185], x[184], x[183], x[191], x[190], x[189], x[324], x[228], x[219], x[218], x[217], x[195], x[323], x[322]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[59], x[58], x[57], x[191], x[190], x[189], x[53], x[52], x[51], x[62], x[61], x[60], x[185], x[184], x[183], x[194], x[193], x[192], x[56], x[55], x[54], x[188], x[187], x[186], x[219], x[218], x[217], x[327], x[231], x[195], x[326], x[325]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[59], x[58], x[57], x[191], x[190], x[189], x[53], x[52], x[51], x[62], x[61], x[60], x[185], x[184], x[183], x[194], x[193], x[192], x[56], x[55], x[54], x[188], x[187], x[186], x[219], x[218], x[217], x[330], x[234], x[195], x[329], x[328]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[89], x[88], x[87], x[149], x[148], x[147], x[98], x[97], x[96], x[95], x[94], x[93], x[158], x[157], x[156], x[155], x[154], x[153], x[92], x[91], x[90], x[152], x[151], x[150], x[333], x[237], x[219], x[218], x[217], x[195], x[332], x[331]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[98], x[97], x[96], x[158], x[157], x[156], x[89], x[88], x[87], x[95], x[94], x[93], x[149], x[148], x[147], x[155], x[154], x[153], x[219], x[218], x[217], x[336], x[240], x[195], x[335], x[334]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[95], x[94], x[93], x[155], x[154], x[153], x[89], x[88], x[87], x[98], x[97], x[96], x[149], x[148], x[147], x[158], x[157], x[156], x[92], x[91], x[90], x[152], x[151], x[150], x[219], x[218], x[217], x[339], x[243], x[195], x[338], x[337]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[95], x[94], x[93], x[155], x[154], x[153], x[89], x[88], x[87], x[98], x[97], x[96], x[149], x[148], x[147], x[158], x[157], x[156], x[92], x[91], x[90], x[152], x[151], x[150], x[342], x[246], x[219], x[218], x[217], x[195], x[341], x[340]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[77], x[76], x[75], x[161], x[160], x[159], x[86], x[85], x[84], x[83], x[82], x[81], x[170], x[169], x[168], x[167], x[166], x[165], x[80], x[79], x[78], x[219], x[218], x[217], x[164], x[163], x[162], x[345], x[249], x[201], x[200], x[199], x[195], x[344], x[343]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[86], x[85], x[84], x[170], x[169], x[168], x[77], x[76], x[75], x[83], x[82], x[81], x[219], x[218], x[217], x[161], x[160], x[159], x[167], x[166], x[165], x[348], x[252], x[207], x[206], x[205], x[195], x[347], x[346]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[83], x[82], x[81], x[167], x[166], x[165], x[77], x[76], x[75], x[86], x[85], x[84], x[161], x[160], x[159], x[170], x[169], x[168], x[80], x[79], x[78], x[219], x[218], x[217], x[164], x[163], x[162], x[351], x[255], x[204], x[203], x[202], x[195], x[350], x[349]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[83], x[82], x[81], x[167], x[166], x[165], x[77], x[76], x[75], x[86], x[85], x[84], x[161], x[160], x[159], x[170], x[169], x[168], x[80], x[79], x[78], x[219], x[218], x[217], x[164], x[163], x[162], x[354], x[258], x[195], x[353], x[352]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[65], x[64], x[63], x[173], x[172], x[171], x[74], x[73], x[72], x[71], x[70], x[69], x[182], x[181], x[180], x[179], x[178], x[177], x[68], x[67], x[66], x[219], x[218], x[217], x[176], x[175], x[174], x[357], x[261], x[210], x[209], x[208], x[195], x[356], x[355]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[74], x[73], x[72], x[182], x[181], x[180], x[65], x[64], x[63], x[71], x[70], x[69], x[219], x[218], x[217], x[173], x[172], x[171], x[179], x[178], x[177], x[360], x[264], x[213], x[212], x[211], x[195], x[359], x[358]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[71], x[70], x[69], x[179], x[178], x[177], x[65], x[64], x[63], x[74], x[73], x[72], x[173], x[172], x[171], x[182], x[181], x[180], x[68], x[67], x[66], x[219], x[218], x[217], x[176], x[175], x[174], x[363], x[267], x[216], x[215], x[214], x[195], x[362], x[361]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[71], x[70], x[69], x[179], x[178], x[177], x[65], x[64], x[63], x[74], x[73], x[72], x[173], x[172], x[171], x[182], x[181], x[180], x[68], x[67], x[66], x[219], x[218], x[217], x[176], x[175], x[174], x[366], x[270], x[198], x[197], x[196], x[195], x[365], x[364]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[185], x[184], x[183], x[101], x[100], x[99], x[17], x[16], x[15], x[194], x[193], x[192], x[191], x[190], x[189], x[110], x[109], x[108], x[107], x[106], x[105], x[26], x[25], x[24], x[23], x[22], x[21], x[188], x[187], x[186], x[104], x[103], x[102], x[20], x[19], x[18], x[219], x[218], x[217], x[225], x[273], x[369], x[195], x[368], x[367]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[194], x[193], x[192], x[110], x[109], x[108], x[26], x[25], x[24], x[185], x[184], x[183], x[191], x[190], x[189], x[101], x[100], x[99], x[107], x[106], x[105], x[17], x[16], x[15], x[23], x[22], x[21], x[219], x[218], x[217], x[228], x[276], x[372], x[195], x[371], x[370]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[191], x[190], x[189], x[107], x[106], x[105], x[23], x[22], x[21], x[185], x[184], x[183], x[194], x[193], x[192], x[101], x[100], x[99], x[110], x[109], x[108], x[17], x[16], x[15], x[26], x[25], x[24], x[188], x[187], x[186], x[104], x[103], x[102], x[20], x[19], x[18], x[219], x[218], x[217], x[231], x[279], x[375], x[195], x[374], x[373]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[191], x[190], x[189], x[107], x[106], x[105], x[23], x[22], x[21], x[185], x[184], x[183], x[194], x[193], x[192], x[101], x[100], x[99], x[110], x[109], x[108], x[17], x[16], x[15], x[26], x[25], x[24], x[188], x[187], x[186], x[104], x[103], x[102], x[20], x[19], x[18], x[219], x[218], x[217], x[234], x[282], x[378], x[195], x[377], x[376]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[149], x[148], x[147], x[137], x[136], x[135], x[29], x[28], x[27], x[158], x[157], x[156], x[155], x[154], x[153], x[146], x[145], x[144], x[143], x[142], x[141], x[38], x[37], x[36], x[35], x[34], x[33], x[152], x[151], x[150], x[140], x[139], x[138], x[32], x[31], x[30], x[219], x[218], x[217], x[237], x[285], x[381], x[195], x[380], x[379]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[158], x[157], x[156], x[146], x[145], x[144], x[38], x[37], x[36], x[149], x[148], x[147], x[155], x[154], x[153], x[137], x[136], x[135], x[143], x[142], x[141], x[29], x[28], x[27], x[35], x[34], x[33], x[240], x[288], x[384], x[219], x[218], x[217], x[195], x[383], x[382]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[155], x[154], x[153], x[143], x[142], x[141], x[35], x[34], x[33], x[149], x[148], x[147], x[158], x[157], x[156], x[137], x[136], x[135], x[146], x[145], x[144], x[29], x[28], x[27], x[38], x[37], x[36], x[152], x[151], x[150], x[140], x[139], x[138], x[32], x[31], x[30], x[243], x[291], x[387], x[219], x[218], x[217], x[195], x[386], x[385]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[155], x[154], x[153], x[143], x[142], x[141], x[35], x[34], x[33], x[149], x[148], x[147], x[158], x[157], x[156], x[137], x[136], x[135], x[146], x[145], x[144], x[29], x[28], x[27], x[38], x[37], x[36], x[152], x[151], x[150], x[140], x[139], x[138], x[32], x[31], x[30], x[219], x[218], x[217], x[246], x[294], x[390], x[195], x[389], x[388]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[161], x[160], x[159], x[125], x[124], x[123], x[41], x[40], x[39], x[170], x[169], x[168], x[167], x[166], x[165], x[134], x[133], x[132], x[131], x[130], x[129], x[50], x[49], x[48], x[47], x[46], x[45], x[164], x[163], x[162], x[128], x[127], x[126], x[44], x[43], x[42], x[249], x[297], x[393], x[219], x[218], x[217], x[195], x[392], x[391]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[170], x[169], x[168], x[134], x[133], x[132], x[50], x[49], x[48], x[161], x[160], x[159], x[167], x[166], x[165], x[125], x[124], x[123], x[131], x[130], x[129], x[41], x[40], x[39], x[47], x[46], x[45], x[219], x[218], x[217], x[252], x[300], x[396], x[195], x[395], x[394]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[167], x[166], x[165], x[131], x[130], x[129], x[47], x[46], x[45], x[161], x[160], x[159], x[170], x[169], x[168], x[125], x[124], x[123], x[134], x[133], x[132], x[41], x[40], x[39], x[50], x[49], x[48], x[164], x[163], x[162], x[128], x[127], x[126], x[44], x[43], x[42], x[219], x[218], x[217], x[255], x[303], x[399], x[195], x[398], x[397]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[167], x[166], x[165], x[131], x[130], x[129], x[47], x[46], x[45], x[161], x[160], x[159], x[170], x[169], x[168], x[125], x[124], x[123], x[134], x[133], x[132], x[41], x[40], x[39], x[50], x[49], x[48], x[164], x[163], x[162], x[128], x[127], x[126], x[44], x[43], x[42], x[258], x[306], x[402], x[219], x[218], x[217], x[195], x[401], x[400]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[173], x[172], x[171], x[113], x[112], x[111], x[5], x[4], x[3], x[182], x[181], x[180], x[179], x[178], x[177], x[122], x[121], x[120], x[119], x[118], x[117], x[14], x[13], x[12], x[11], x[10], x[9], x[176], x[175], x[174], x[116], x[115], x[114], x[8], x[7], x[6], x[219], x[218], x[217], x[261], x[309], x[405], x[195], x[404], x[403]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[182], x[181], x[180], x[122], x[121], x[120], x[14], x[13], x[12], x[173], x[172], x[171], x[179], x[178], x[177], x[113], x[112], x[111], x[119], x[118], x[117], x[5], x[4], x[3], x[11], x[10], x[9], x[219], x[218], x[217], x[264], x[312], x[408], x[195], x[407], x[406]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[179], x[178], x[177], x[119], x[118], x[117], x[11], x[10], x[9], x[173], x[172], x[171], x[182], x[181], x[180], x[113], x[112], x[111], x[122], x[121], x[120], x[5], x[4], x[3], x[14], x[13], x[12], x[176], x[175], x[174], x[116], x[115], x[114], x[8], x[7], x[6], x[267], x[315], x[411], x[219], x[218], x[217], x[195], x[410], x[409]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[179], x[178], x[177], x[119], x[118], x[117], x[11], x[10], x[9], x[173], x[172], x[171], x[182], x[181], x[180], x[113], x[112], x[111], x[122], x[121], x[120], x[5], x[4], x[3], x[14], x[13], x[12], x[176], x[175], x[174], x[116], x[115], x[114], x[8], x[7], x[6], x[219], x[218], x[217], x[270], x[318], x[414], x[195], x[413], x[412]}), .y(y[138]));
endmodule

module R2ind0(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (t[2] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[1];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [21:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[11] = ~x[0] & t[18];
  assign t[12] = ~x[0] & t[19];
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[27] ^ x[3];
  assign t[21] = t[28] ^ x[6];
  assign t[22] = t[29] ^ x[9];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[18];
  assign t[26] = t[33] ^ x[21];
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[40] & ~t[41]);
  assign t[31] = (t[42] & ~t[43]);
  assign t[32] = (t[44] & ~t[45]);
  assign t[33] = (t[46] & ~t[47]);
  assign t[34] = t[48] ^ x[3];
  assign t[35] = t[49] ^ x[2];
  assign t[36] = t[50] ^ x[6];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[9];
  assign t[39] = t[53] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[11];
  assign t[42] = t[56] ^ x[15];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[17];
  assign t[46] = t[60] ^ x[21];
  assign t[47] = t[61] ^ x[20];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = (x[4]);
  assign t[51] = (x[4]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[10]);
  assign t[55] = (x[10]);
  assign t[56] = (x[13]);
  assign t[57] = (x[13]);
  assign t[58] = (x[16]);
  assign t[59] = (x[16]);
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = (x[19]);
  assign t[61] = (x[19]);
  assign t[6] = ~x[0] & t[15];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0]);
endmodule

module R2ind3(x, y);
 input [21:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(~x[0] & ~t[17]);
  assign t[11] = ~x[0] & t[18];
  assign t[12] = ~x[0] & t[19];
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = (t[26]);
  assign t[1] = ~x[0] & t[13];
  assign t[20] = t[27] ^ x[3];
  assign t[21] = t[28] ^ x[6];
  assign t[22] = t[29] ^ x[9];
  assign t[23] = t[30] ^ x[12];
  assign t[24] = t[31] ^ x[15];
  assign t[25] = t[32] ^ x[18];
  assign t[26] = t[33] ^ x[21];
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[40] & ~t[41]);
  assign t[31] = (t[42] & ~t[43]);
  assign t[32] = (t[44] & ~t[45]);
  assign t[33] = (t[46] & ~t[47]);
  assign t[34] = t[48] ^ x[3];
  assign t[35] = t[49] ^ x[2];
  assign t[36] = t[50] ^ x[6];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[9];
  assign t[39] = t[53] ^ x[8];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[11];
  assign t[42] = t[56] ^ x[15];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[17];
  assign t[46] = t[60] ^ x[21];
  assign t[47] = t[61] ^ x[20];
  assign t[48] = (x[1]);
  assign t[49] = (x[1]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[50] = (x[4]);
  assign t[51] = (x[4]);
  assign t[52] = (x[7]);
  assign t[53] = (x[7]);
  assign t[54] = (x[10]);
  assign t[55] = (x[10]);
  assign t[56] = (x[13]);
  assign t[57] = (x[13]);
  assign t[58] = (x[16]);
  assign t[59] = (x[16]);
  assign t[5] = ~(~x[0] & ~t[14]);
  assign t[60] = (x[19]);
  assign t[61] = (x[19]);
  assign t[6] = ~x[0] & t[15];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~x[0] & t[16];
  assign y = (t[0]);
endmodule

module R2ind4(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind5(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind6(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~x[0] & t[3];
  assign t[2] = ~(~x[0] & ~t[4]);
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [3:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[3];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[3];
  assign t[5] = t[7] ^ x[2];
  assign t[6] = (x[1]);
  assign t[7] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = ~x[0] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [6:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[5];
  assign t[13] = (x[1]);
  assign t[14] = (x[1]);
  assign t[15] = (x[4]);
  assign t[16] = (x[4]);
  assign t[1] = ~(~x[0] & ~t[3]);
  assign t[2] = ~x[0] & t[4];
  assign t[3] = (t[5]);
  assign t[4] = (t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[6];
  assign t[7] = (t[9] & ~t[10]);
  assign t[8] = (t[11] & ~t[12]);
  assign t[9] = t[13] ^ x[3];
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~x[0] & t[2];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [3:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = ~x[0] & t[2];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[3];
  assign t[4] = (t[5] & ~t[6]);
  assign t[5] = t[7] ^ x[3];
  assign t[6] = t[8] ^ x[2];
  assign t[7] = (x[1]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [6:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[2];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[5];
  assign t[14] = (x[1]);
  assign t[15] = (x[1]);
  assign t[16] = (x[4]);
  assign t[17] = (x[4]);
  assign t[1] = ~t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = ~x[0] & t[5];
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[6];
  assign t[8] = (t[10] & ~t[11]);
  assign t[9] = (t[12] & ~t[13]);
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [6:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[2];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[5];
  assign t[14] = (x[1]);
  assign t[15] = (x[1]);
  assign t[16] = (x[4]);
  assign t[17] = (x[4]);
  assign t[1] = ~t[3];
  assign t[2] = ~x[0] & t[4];
  assign t[3] = ~x[0] & t[5];
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[3];
  assign t[7] = t[9] ^ x[6];
  assign t[8] = (t[10] & ~t[11]);
  assign t[9] = (t[12] & ~t[13]);
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind26(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind27(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind28(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind29(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind31(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind36(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind41(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind46(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind51(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind56(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind61(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind66(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [18:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[8]);
  assign t[11] = ~(t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[15];
  assign t[21] = t[26] ^ x[18];
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = (t[33] & ~t[34]);
  assign t[26] = (t[35] & ~t[36]);
  assign t[27] = t[37] ^ x[6];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[15];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[18];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = (x[4]);
  assign t[38] = (x[4]);
  assign t[39] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[10]);
  assign t[42] = (x[10]);
  assign t[43] = (x[13]);
  assign t[44] = (x[13]);
  assign t[45] = (x[16]);
  assign t[46] = (x[16]);
  assign t[4] = ~x[2] & t[12];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = t[10] | t[13];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [18:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[8]);
  assign t[11] = ~(t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[15];
  assign t[21] = t[26] ^ x[18];
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = (t[33] & ~t[34]);
  assign t[26] = (t[35] & ~t[36]);
  assign t[27] = t[37] ^ x[6];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[15];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[18];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = (x[4]);
  assign t[38] = (x[4]);
  assign t[39] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[10]);
  assign t[42] = (x[10]);
  assign t[43] = (x[13]);
  assign t[44] = (x[13]);
  assign t[45] = (x[16]);
  assign t[46] = (x[16]);
  assign t[4] = ~x[2] & t[12];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = t[10] | t[13];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind71(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[12]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [15:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = t[22] ^ x[15];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = ~t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[15];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[14];
  assign t[31] = (x[4]);
  assign t[32] = (x[4]);
  assign t[33] = (x[7]);
  assign t[34] = (x[7]);
  assign t[35] = (x[10]);
  assign t[36] = (x[10]);
  assign t[37] = (x[13]);
  assign t[38] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~x[2] & t[11];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[12] & t[8]);
  assign t[7] = ~(t[13] & t[9]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[14] & t[10]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [15:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[12]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = t[22] ^ x[15];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = ~t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[15];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[14];
  assign t[31] = (x[4]);
  assign t[32] = (x[4]);
  assign t[33] = (x[7]);
  assign t[34] = (x[7]);
  assign t[35] = (x[10]);
  assign t[36] = (x[10]);
  assign t[37] = (x[13]);
  assign t[38] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[4] = ~x[2] & t[11];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[12] & t[8]);
  assign t[7] = ~(t[13] & t[9]);
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[14] & t[10]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[16] & t[15]);
  assign t[12] = ~(t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = t[23] ^ x[6];
  assign t[19] = t[24] ^ x[9];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[12];
  assign t[21] = t[26] ^ x[15];
  assign t[22] = t[27] ^ x[18];
  assign t[23] = (t[28] & ~t[29]);
  assign t[24] = (t[30] & ~t[31]);
  assign t[25] = (t[32] & ~t[33]);
  assign t[26] = (t[34] & ~t[35]);
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = t[38] ^ x[6];
  assign t[29] = t[39] ^ x[5];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[9];
  assign t[31] = t[41] ^ x[8];
  assign t[32] = t[42] ^ x[12];
  assign t[33] = t[43] ^ x[11];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[14];
  assign t[36] = t[46] ^ x[18];
  assign t[37] = t[47] ^ x[17];
  assign t[38] = (x[4]);
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[7]);
  assign t[42] = (x[10]);
  assign t[43] = (x[10]);
  assign t[44] = (x[13]);
  assign t[45] = (x[13]);
  assign t[46] = (x[16]);
  assign t[47] = (x[16]);
  assign t[4] = ~x[2] & t[13];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10] & t[14]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16]);
  assign y = (t[0]);
endmodule

module R2ind76(x, y);
 input [18:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[8]);
  assign t[11] = ~(t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[15];
  assign t[21] = t[26] ^ x[18];
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = (t[33] & ~t[34]);
  assign t[26] = (t[35] & ~t[36]);
  assign t[27] = t[37] ^ x[6];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[15];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[18];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = (x[4]);
  assign t[38] = (x[4]);
  assign t[39] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[10]);
  assign t[42] = (x[10]);
  assign t[43] = (x[13]);
  assign t[44] = (x[13]);
  assign t[45] = (x[16]);
  assign t[46] = (x[16]);
  assign t[4] = ~x[2] & t[12];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = t[10] | t[13];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [18:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[11] | t[8]);
  assign t[11] = ~(t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = t[22] ^ x[6];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[15];
  assign t[21] = t[26] ^ x[18];
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = (t[33] & ~t[34]);
  assign t[26] = (t[35] & ~t[36]);
  assign t[27] = t[37] ^ x[6];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[9];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[15];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[18];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = (x[4]);
  assign t[38] = (x[4]);
  assign t[39] = (x[7]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[7]);
  assign t[41] = (x[10]);
  assign t[42] = (x[10]);
  assign t[43] = (x[13]);
  assign t[44] = (x[13]);
  assign t[45] = (x[16]);
  assign t[46] = (x[16]);
  assign t[4] = ~x[2] & t[12];
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = t[10] | t[13];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[19]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[15] | t[12]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind81(x, y);
 input [15:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[16] & t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = (t[19]);
  assign t[16] = (t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[9];
  assign t[19] = t[23] ^ x[12];
  assign t[1] = ~t[3];
  assign t[20] = t[24] ^ x[15];
  assign t[21] = (t[25] & ~t[26]);
  assign t[22] = (t[27] & ~t[28]);
  assign t[23] = (t[29] & ~t[30]);
  assign t[24] = (t[31] & ~t[32]);
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[8];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[38] ^ x[11];
  assign t[31] = t[39] ^ x[15];
  assign t[32] = t[40] ^ x[14];
  assign t[33] = (x[4]);
  assign t[34] = (x[4]);
  assign t[35] = (x[7]);
  assign t[36] = (x[7]);
  assign t[37] = (x[10]);
  assign t[38] = (x[10]);
  assign t[39] = (x[13]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[13]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[13] & t[10]);
  assign t[8] = ~(t[14] & t[11]);
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [18:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[18] & t[17]);
  assign t[14] = ~(t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = (t[24]);
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[6];
  assign t[21] = t[26] ^ x[9];
  assign t[22] = t[27] ^ x[12];
  assign t[23] = t[28] ^ x[15];
  assign t[24] = t[29] ^ x[18];
  assign t[25] = (t[30] & ~t[31]);
  assign t[26] = (t[32] & ~t[33]);
  assign t[27] = (t[34] & ~t[35]);
  assign t[28] = (t[36] & ~t[37]);
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[6];
  assign t[31] = t[41] ^ x[5];
  assign t[32] = t[42] ^ x[9];
  assign t[33] = t[43] ^ x[8];
  assign t[34] = t[44] ^ x[12];
  assign t[35] = t[45] ^ x[11];
  assign t[36] = t[46] ^ x[15];
  assign t[37] = t[47] ^ x[14];
  assign t[38] = t[48] ^ x[18];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[4]);
  assign t[42] = (x[7]);
  assign t[43] = (x[7]);
  assign t[44] = (x[10]);
  assign t[45] = (x[10]);
  assign t[46] = (x[13]);
  assign t[47] = (x[13]);
  assign t[48] = (x[16]);
  assign t[49] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[15]);
  assign t[9] = ~x[2] & t[16];
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [18:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16]);
  assign t[11] = ~(t[17]);
  assign t[12] = ~(t[13] | t[10]);
  assign t[13] = ~(t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = (t[21]);
  assign t[17] = (t[22]);
  assign t[18] = (t[23]);
  assign t[19] = t[24] ^ x[6];
  assign t[1] = ~t[3];
  assign t[20] = t[25] ^ x[9];
  assign t[21] = t[26] ^ x[12];
  assign t[22] = t[27] ^ x[15];
  assign t[23] = t[28] ^ x[18];
  assign t[24] = (t[29] & ~t[30]);
  assign t[25] = (t[31] & ~t[32]);
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = t[39] ^ x[6];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[40] ^ x[5];
  assign t[31] = t[41] ^ x[9];
  assign t[32] = t[42] ^ x[8];
  assign t[33] = t[43] ^ x[12];
  assign t[34] = t[44] ^ x[11];
  assign t[35] = t[45] ^ x[15];
  assign t[36] = t[46] ^ x[14];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = t[48] ^ x[17];
  assign t[39] = (x[4]);
  assign t[3] = x[2] ? x[3] : t[5];
  assign t[40] = (x[4]);
  assign t[41] = (x[7]);
  assign t[42] = (x[7]);
  assign t[43] = (x[10]);
  assign t[44] = (x[10]);
  assign t[45] = (x[13]);
  assign t[46] = (x[13]);
  assign t[47] = (x[16]);
  assign t[48] = (x[16]);
  assign t[4] = ~(t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = t[12] | t[14];
  assign t[9] = ~x[2] & t[15];
  assign y = (t[0]);
endmodule

module R2ind86(x, y);
 input [31:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[27] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[28] | t[21]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[31];
  assign t[44] = (t[53] & ~t[54]);
  assign t[45] = (t[55] & ~t[56]);
  assign t[46] = (t[57] & ~t[58]);
  assign t[47] = (t[59] & ~t[60]);
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = t[71] ^ x[7];
  assign t[54] = t[72] ^ x[6];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[13];
  assign t[58] = t[76] ^ x[12];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[22];
  assign t[64] = t[82] ^ x[21];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[24];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[27];
  assign t[69] = t[87] ^ x[31];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = (x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8]);
  assign t[74] = (x[8]);
  assign t[75] = (x[11]);
  assign t[76] = (x[11]);
  assign t[77] = (x[14]);
  assign t[78] = (x[14]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17]);
  assign t[81] = (x[20]);
  assign t[82] = (x[20]);
  assign t[83] = (x[23]);
  assign t[84] = (x[23]);
  assign t[85] = (x[26]);
  assign t[86] = (x[26]);
  assign t[87] = (x[29]);
  assign t[88] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [31:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[27] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[28] | t[21]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[31];
  assign t[44] = (t[53] & ~t[54]);
  assign t[45] = (t[55] & ~t[56]);
  assign t[46] = (t[57] & ~t[58]);
  assign t[47] = (t[59] & ~t[60]);
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = t[71] ^ x[7];
  assign t[54] = t[72] ^ x[6];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[13];
  assign t[58] = t[76] ^ x[12];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[22];
  assign t[64] = t[82] ^ x[21];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[24];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[27];
  assign t[69] = t[87] ^ x[31];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = (x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8]);
  assign t[74] = (x[8]);
  assign t[75] = (x[11]);
  assign t[76] = (x[11]);
  assign t[77] = (x[14]);
  assign t[78] = (x[14]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17]);
  assign t[81] = (x[20]);
  assign t[82] = (x[20]);
  assign t[83] = (x[23]);
  assign t[84] = (x[23]);
  assign t[85] = (x[26]);
  assign t[86] = (x[26]);
  assign t[87] = (x[29]);
  assign t[88] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[25] & t[18]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[26] & t[19]);
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[23]);
  assign t[1] = ~t[3];
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = (t[33]);
  assign t[27] = t[34] ^ x[5];
  assign t[28] = t[35] ^ x[10];
  assign t[29] = t[36] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[16];
  assign t[31] = t[38] ^ x[19];
  assign t[32] = t[39] ^ x[22];
  assign t[33] = t[40] ^ x[25];
  assign t[34] = (t[41] & ~t[42]);
  assign t[35] = (t[43] & ~t[44]);
  assign t[36] = (t[45] & ~t[46]);
  assign t[37] = (t[47] & ~t[48]);
  assign t[38] = (t[49] & ~t[50]);
  assign t[39] = (t[51] & ~t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53] & ~t[54]);
  assign t[41] = t[55] ^ x[5];
  assign t[42] = t[56] ^ x[4];
  assign t[43] = t[57] ^ x[10];
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[13];
  assign t[46] = t[60] ^ x[12];
  assign t[47] = t[61] ^ x[16];
  assign t[48] = t[62] ^ x[15];
  assign t[49] = t[63] ^ x[19];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[22];
  assign t[52] = t[66] ^ x[21];
  assign t[53] = t[67] ^ x[25];
  assign t[54] = t[68] ^ x[24];
  assign t[55] = (x[3]);
  assign t[56] = (x[3]);
  assign t[57] = (x[8]);
  assign t[58] = (x[8]);
  assign t[59] = (x[11]);
  assign t[5] = ~t[7];
  assign t[60] = (x[11]);
  assign t[61] = (x[14]);
  assign t[62] = (x[14]);
  assign t[63] = (x[17]);
  assign t[64] = (x[17]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[23]);
  assign t[68] = (x[23]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21] & t[14]);
  assign t[11] = ~(t[22] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[25] & t[18]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[26] & t[19]);
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[23]);
  assign t[1] = ~t[3];
  assign t[20] = (t[27]);
  assign t[21] = (t[28]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = (t[33]);
  assign t[27] = t[34] ^ x[5];
  assign t[28] = t[35] ^ x[10];
  assign t[29] = t[36] ^ x[13];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[16];
  assign t[31] = t[38] ^ x[19];
  assign t[32] = t[39] ^ x[22];
  assign t[33] = t[40] ^ x[25];
  assign t[34] = (t[41] & ~t[42]);
  assign t[35] = (t[43] & ~t[44]);
  assign t[36] = (t[45] & ~t[46]);
  assign t[37] = (t[47] & ~t[48]);
  assign t[38] = (t[49] & ~t[50]);
  assign t[39] = (t[51] & ~t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53] & ~t[54]);
  assign t[41] = t[55] ^ x[5];
  assign t[42] = t[56] ^ x[4];
  assign t[43] = t[57] ^ x[10];
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[13];
  assign t[46] = t[60] ^ x[12];
  assign t[47] = t[61] ^ x[16];
  assign t[48] = t[62] ^ x[15];
  assign t[49] = t[63] ^ x[19];
  assign t[4] = ~x[2] & t[20];
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[22];
  assign t[52] = t[66] ^ x[21];
  assign t[53] = t[67] ^ x[25];
  assign t[54] = t[68] ^ x[24];
  assign t[55] = (x[3]);
  assign t[56] = (x[3]);
  assign t[57] = (x[8]);
  assign t[58] = (x[8]);
  assign t[59] = (x[11]);
  assign t[5] = ~t[7];
  assign t[60] = (x[11]);
  assign t[61] = (x[14]);
  assign t[62] = (x[14]);
  assign t[63] = (x[17]);
  assign t[64] = (x[17]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[23]);
  assign t[68] = (x[23]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [31:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[27]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[32] & t[31]);
  assign t[25] = ~(t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[31];
  assign t[44] = (t[53] & ~t[54]);
  assign t[45] = (t[55] & ~t[56]);
  assign t[46] = (t[57] & ~t[58]);
  assign t[47] = (t[59] & ~t[60]);
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = t[71] ^ x[7];
  assign t[54] = t[72] ^ x[6];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[13];
  assign t[58] = t[76] ^ x[12];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[22];
  assign t[64] = t[82] ^ x[21];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[24];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[27];
  assign t[69] = t[87] ^ x[31];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = (x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8]);
  assign t[74] = (x[8]);
  assign t[75] = (x[11]);
  assign t[76] = (x[11]);
  assign t[77] = (x[14]);
  assign t[78] = (x[14]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17]);
  assign t[81] = (x[20]);
  assign t[82] = (x[20]);
  assign t[83] = (x[23]);
  assign t[84] = (x[23]);
  assign t[85] = (x[26]);
  assign t[86] = (x[26]);
  assign t[87] = (x[29]);
  assign t[88] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind91(x, y);
 input [31:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[27]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[32] & t[31]);
  assign t[25] = ~(t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[31];
  assign t[44] = (t[53] & ~t[54]);
  assign t[45] = (t[55] & ~t[56]);
  assign t[46] = (t[57] & ~t[58]);
  assign t[47] = (t[59] & ~t[60]);
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = t[71] ^ x[7];
  assign t[54] = t[72] ^ x[6];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[13];
  assign t[58] = t[76] ^ x[12];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[22];
  assign t[64] = t[82] ^ x[21];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[24];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[27];
  assign t[69] = t[87] ^ x[31];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = (x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8]);
  assign t[74] = (x[8]);
  assign t[75] = (x[11]);
  assign t[76] = (x[11]);
  assign t[77] = (x[14]);
  assign t[78] = (x[14]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17]);
  assign t[81] = (x[20]);
  assign t[82] = (x[20]);
  assign t[83] = (x[23]);
  assign t[84] = (x[23]);
  assign t[85] = (x[26]);
  assign t[86] = (x[26]);
  assign t[87] = (x[29]);
  assign t[88] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[24];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = t[18] | t[25];
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = t[21] | t[26];
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[22] | t[16]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[23] | t[19]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = t[42] ^ x[7];
  assign t[34] = t[43] ^ x[10];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[22];
  assign t[39] = t[48] ^ x[25];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[28];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = (t[51] & ~t[52]);
  assign t[43] = (t[53] & ~t[54]);
  assign t[44] = (t[55] & ~t[56]);
  assign t[45] = (t[57] & ~t[58]);
  assign t[46] = (t[59] & ~t[60]);
  assign t[47] = (t[61] & ~t[62]);
  assign t[48] = (t[63] & ~t[64]);
  assign t[49] = (t[65] & ~t[66]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[67] & ~t[68]);
  assign t[51] = t[69] ^ x[7];
  assign t[52] = t[70] ^ x[6];
  assign t[53] = t[71] ^ x[10];
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[13];
  assign t[56] = t[74] ^ x[12];
  assign t[57] = t[75] ^ x[16];
  assign t[58] = t[76] ^ x[15];
  assign t[59] = t[77] ^ x[19];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[22];
  assign t[62] = t[80] ^ x[21];
  assign t[63] = t[81] ^ x[25];
  assign t[64] = t[82] ^ x[24];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[31];
  assign t[68] = t[86] ^ x[30];
  assign t[69] = (x[5]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[5]);
  assign t[71] = (x[8]);
  assign t[72] = (x[8]);
  assign t[73] = (x[11]);
  assign t[74] = (x[11]);
  assign t[75] = (x[14]);
  assign t[76] = (x[14]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[20]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[20]);
  assign t[81] = (x[23]);
  assign t[82] = (x[23]);
  assign t[83] = (x[26]);
  assign t[84] = (x[26]);
  assign t[85] = (x[29]);
  assign t[86] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[24];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = t[18] | t[25];
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = t[21] | t[26];
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[22] | t[16]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[23] | t[19]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = t[42] ^ x[7];
  assign t[34] = t[43] ^ x[10];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[22];
  assign t[39] = t[48] ^ x[25];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[28];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = (t[51] & ~t[52]);
  assign t[43] = (t[53] & ~t[54]);
  assign t[44] = (t[55] & ~t[56]);
  assign t[45] = (t[57] & ~t[58]);
  assign t[46] = (t[59] & ~t[60]);
  assign t[47] = (t[61] & ~t[62]);
  assign t[48] = (t[63] & ~t[64]);
  assign t[49] = (t[65] & ~t[66]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[67] & ~t[68]);
  assign t[51] = t[69] ^ x[7];
  assign t[52] = t[70] ^ x[6];
  assign t[53] = t[71] ^ x[10];
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[13];
  assign t[56] = t[74] ^ x[12];
  assign t[57] = t[75] ^ x[16];
  assign t[58] = t[76] ^ x[15];
  assign t[59] = t[77] ^ x[19];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[22];
  assign t[62] = t[80] ^ x[21];
  assign t[63] = t[81] ^ x[25];
  assign t[64] = t[82] ^ x[24];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[31];
  assign t[68] = t[86] ^ x[30];
  assign t[69] = (x[5]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[5]);
  assign t[71] = (x[8]);
  assign t[72] = (x[8]);
  assign t[73] = (x[11]);
  assign t[74] = (x[11]);
  assign t[75] = (x[14]);
  assign t[76] = (x[14]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[20]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[20]);
  assign t[81] = (x[23]);
  assign t[82] = (x[23]);
  assign t[83] = (x[26]);
  assign t[84] = (x[26]);
  assign t[85] = (x[29]);
  assign t[86] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[25] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[26] | t[19]);
  assign t[14] = ~(t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[27] | t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = t[42] ^ x[5];
  assign t[34] = t[43] ^ x[10];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[22];
  assign t[39] = t[48] ^ x[25];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[28];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = (t[51] & ~t[52]);
  assign t[43] = (t[53] & ~t[54]);
  assign t[44] = (t[55] & ~t[56]);
  assign t[45] = (t[57] & ~t[58]);
  assign t[46] = (t[59] & ~t[60]);
  assign t[47] = (t[61] & ~t[62]);
  assign t[48] = (t[63] & ~t[64]);
  assign t[49] = (t[65] & ~t[66]);
  assign t[4] = ~x[2] & t[24];
  assign t[50] = (t[67] & ~t[68]);
  assign t[51] = t[69] ^ x[5];
  assign t[52] = t[70] ^ x[4];
  assign t[53] = t[71] ^ x[10];
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[13];
  assign t[56] = t[74] ^ x[12];
  assign t[57] = t[75] ^ x[16];
  assign t[58] = t[76] ^ x[15];
  assign t[59] = t[77] ^ x[19];
  assign t[5] = ~t[7];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[22];
  assign t[62] = t[80] ^ x[21];
  assign t[63] = t[81] ^ x[25];
  assign t[64] = t[82] ^ x[24];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[31];
  assign t[68] = t[86] ^ x[30];
  assign t[69] = (x[3]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (x[3]);
  assign t[71] = (x[8]);
  assign t[72] = (x[8]);
  assign t[73] = (x[11]);
  assign t[74] = (x[11]);
  assign t[75] = (x[14]);
  assign t[76] = (x[14]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[20]);
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[80] = (x[20]);
  assign t[81] = (x[23]);
  assign t[82] = (x[23]);
  assign t[83] = (x[26]);
  assign t[84] = (x[26]);
  assign t[85] = (x[29]);
  assign t[86] = (x[29]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [31:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[25] | t[16]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[26] | t[19]);
  assign t[14] = ~(t[27]);
  assign t[15] = ~(t[28]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[29]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[27] | t[28]);
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = t[42] ^ x[5];
  assign t[34] = t[43] ^ x[10];
  assign t[35] = t[44] ^ x[13];
  assign t[36] = t[45] ^ x[16];
  assign t[37] = t[46] ^ x[19];
  assign t[38] = t[47] ^ x[22];
  assign t[39] = t[48] ^ x[25];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[28];
  assign t[41] = t[50] ^ x[31];
  assign t[42] = (t[51] & ~t[52]);
  assign t[43] = (t[53] & ~t[54]);
  assign t[44] = (t[55] & ~t[56]);
  assign t[45] = (t[57] & ~t[58]);
  assign t[46] = (t[59] & ~t[60]);
  assign t[47] = (t[61] & ~t[62]);
  assign t[48] = (t[63] & ~t[64]);
  assign t[49] = (t[65] & ~t[66]);
  assign t[4] = ~x[2] & t[24];
  assign t[50] = (t[67] & ~t[68]);
  assign t[51] = t[69] ^ x[5];
  assign t[52] = t[70] ^ x[4];
  assign t[53] = t[71] ^ x[10];
  assign t[54] = t[72] ^ x[9];
  assign t[55] = t[73] ^ x[13];
  assign t[56] = t[74] ^ x[12];
  assign t[57] = t[75] ^ x[16];
  assign t[58] = t[76] ^ x[15];
  assign t[59] = t[77] ^ x[19];
  assign t[5] = ~t[7];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[22];
  assign t[62] = t[80] ^ x[21];
  assign t[63] = t[81] ^ x[25];
  assign t[64] = t[82] ^ x[24];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[31];
  assign t[68] = t[86] ^ x[30];
  assign t[69] = (x[3]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (x[3]);
  assign t[71] = (x[8]);
  assign t[72] = (x[8]);
  assign t[73] = (x[11]);
  assign t[74] = (x[11]);
  assign t[75] = (x[14]);
  assign t[76] = (x[14]);
  assign t[77] = (x[17]);
  assign t[78] = (x[17]);
  assign t[79] = (x[20]);
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[80] = (x[20]);
  assign t[81] = (x[23]);
  assign t[82] = (x[23]);
  assign t[83] = (x[26]);
  assign t[84] = (x[26]);
  assign t[85] = (x[29]);
  assign t[86] = (x[29]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind96(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[22];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25] & t[18]);
  assign t[15] = ~(t[26] & t[19]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[27] & t[20]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[28] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[25]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = (t[33]);
  assign t[27] = (t[34]);
  assign t[28] = (t[35]);
  assign t[29] = t[36] ^ x[7];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[10];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[16];
  assign t[33] = t[40] ^ x[19];
  assign t[34] = t[41] ^ x[22];
  assign t[35] = t[42] ^ x[25];
  assign t[36] = (t[43] & ~t[44]);
  assign t[37] = (t[45] & ~t[46]);
  assign t[38] = (t[47] & ~t[48]);
  assign t[39] = (t[49] & ~t[50]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[51] & ~t[52]);
  assign t[41] = (t[53] & ~t[54]);
  assign t[42] = (t[55] & ~t[56]);
  assign t[43] = t[57] ^ x[7];
  assign t[44] = t[58] ^ x[6];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[9];
  assign t[47] = t[61] ^ x[13];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[16];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[15];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[25];
  assign t[56] = t[70] ^ x[24];
  assign t[57] = (x[5]);
  assign t[58] = (x[5]);
  assign t[59] = (x[8]);
  assign t[5] = ~t[8];
  assign t[60] = (x[8]);
  assign t[61] = (x[11]);
  assign t[62] = (x[11]);
  assign t[63] = (x[14]);
  assign t[64] = (x[14]);
  assign t[65] = (x[17]);
  assign t[66] = (x[17]);
  assign t[67] = (x[20]);
  assign t[68] = (x[20]);
  assign t[69] = (x[23]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[23]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [25:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[22];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[23] & t[16]);
  assign t[13] = ~(t[24] & t[17]);
  assign t[14] = ~(t[25] & t[18]);
  assign t[15] = ~(t[26] & t[19]);
  assign t[16] = ~(t[27]);
  assign t[17] = ~(t[27] & t[20]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[28] & t[21]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[25]);
  assign t[22] = (t[29]);
  assign t[23] = (t[30]);
  assign t[24] = (t[31]);
  assign t[25] = (t[32]);
  assign t[26] = (t[33]);
  assign t[27] = (t[34]);
  assign t[28] = (t[35]);
  assign t[29] = t[36] ^ x[7];
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = t[37] ^ x[10];
  assign t[31] = t[38] ^ x[13];
  assign t[32] = t[39] ^ x[16];
  assign t[33] = t[40] ^ x[19];
  assign t[34] = t[41] ^ x[22];
  assign t[35] = t[42] ^ x[25];
  assign t[36] = (t[43] & ~t[44]);
  assign t[37] = (t[45] & ~t[46]);
  assign t[38] = (t[47] & ~t[48]);
  assign t[39] = (t[49] & ~t[50]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[51] & ~t[52]);
  assign t[41] = (t[53] & ~t[54]);
  assign t[42] = (t[55] & ~t[56]);
  assign t[43] = t[57] ^ x[7];
  assign t[44] = t[58] ^ x[6];
  assign t[45] = t[59] ^ x[10];
  assign t[46] = t[60] ^ x[9];
  assign t[47] = t[61] ^ x[13];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[16];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[15];
  assign t[51] = t[65] ^ x[19];
  assign t[52] = t[66] ^ x[18];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[25];
  assign t[56] = t[70] ^ x[24];
  assign t[57] = (x[5]);
  assign t[58] = (x[5]);
  assign t[59] = (x[8]);
  assign t[5] = ~t[8];
  assign t[60] = (x[8]);
  assign t[61] = (x[11]);
  assign t[62] = (x[11]);
  assign t[63] = (x[14]);
  assign t[64] = (x[14]);
  assign t[65] = (x[17]);
  assign t[66] = (x[17]);
  assign t[67] = (x[20]);
  assign t[68] = (x[20]);
  assign t[69] = (x[23]);
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[23]);
  assign t[7] = ~(t[10]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [31:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[27]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[32] & t[31]);
  assign t[25] = ~(t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[31];
  assign t[44] = (t[53] & ~t[54]);
  assign t[45] = (t[55] & ~t[56]);
  assign t[46] = (t[57] & ~t[58]);
  assign t[47] = (t[59] & ~t[60]);
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = t[71] ^ x[7];
  assign t[54] = t[72] ^ x[6];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[13];
  assign t[58] = t[76] ^ x[12];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[22];
  assign t[64] = t[82] ^ x[21];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[24];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[27];
  assign t[69] = t[87] ^ x[31];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = (x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8]);
  assign t[74] = (x[8]);
  assign t[75] = (x[11]);
  assign t[76] = (x[11]);
  assign t[77] = (x[14]);
  assign t[78] = (x[14]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17]);
  assign t[81] = (x[20]);
  assign t[82] = (x[20]);
  assign t[83] = (x[23]);
  assign t[84] = (x[23]);
  assign t[85] = (x[26]);
  assign t[86] = (x[26]);
  assign t[87] = (x[29]);
  assign t[88] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [31:0] x;
 output y;

 wire [88:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~x[2] & t[26];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[27]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[28]);
  assign t[16] = ~(t[29]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[31]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[32]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = ~(t[33]);
  assign t[24] = ~(t[32] & t[31]);
  assign t[25] = ~(t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = (t[43]);
  assign t[35] = t[44] ^ x[7];
  assign t[36] = t[45] ^ x[10];
  assign t[37] = t[46] ^ x[13];
  assign t[38] = t[47] ^ x[16];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[22];
  assign t[41] = t[50] ^ x[25];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[31];
  assign t[44] = (t[53] & ~t[54]);
  assign t[45] = (t[55] & ~t[56]);
  assign t[46] = (t[57] & ~t[58]);
  assign t[47] = (t[59] & ~t[60]);
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = t[71] ^ x[7];
  assign t[54] = t[72] ^ x[6];
  assign t[55] = t[73] ^ x[10];
  assign t[56] = t[74] ^ x[9];
  assign t[57] = t[75] ^ x[13];
  assign t[58] = t[76] ^ x[12];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[22];
  assign t[64] = t[82] ^ x[21];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[24];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[27];
  assign t[69] = t[87] ^ x[31];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = (x[5]);
  assign t[72] = (x[5]);
  assign t[73] = (x[8]);
  assign t[74] = (x[8]);
  assign t[75] = (x[11]);
  assign t[76] = (x[11]);
  assign t[77] = (x[14]);
  assign t[78] = (x[14]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[17]);
  assign t[81] = (x[20]);
  assign t[82] = (x[20]);
  assign t[83] = (x[23]);
  assign t[84] = (x[23]);
  assign t[85] = (x[26]);
  assign t[86] = (x[26]);
  assign t[87] = (x[29]);
  assign t[88] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [31:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = t[16] | t[23];
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[24];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[20] | t[14]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[21] | t[17]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29]);
  assign t[21] = ~(t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = t[40] ^ x[5];
  assign t[32] = t[41] ^ x[10];
  assign t[33] = t[42] ^ x[13];
  assign t[34] = t[43] ^ x[16];
  assign t[35] = t[44] ^ x[19];
  assign t[36] = t[45] ^ x[22];
  assign t[37] = t[46] ^ x[25];
  assign t[38] = t[47] ^ x[28];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[52]);
  assign t[42] = (t[53] & ~t[54]);
  assign t[43] = (t[55] & ~t[56]);
  assign t[44] = (t[57] & ~t[58]);
  assign t[45] = (t[59] & ~t[60]);
  assign t[46] = (t[61] & ~t[62]);
  assign t[47] = (t[63] & ~t[64]);
  assign t[48] = (t[65] & ~t[66]);
  assign t[49] = t[67] ^ x[5];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[68] ^ x[4];
  assign t[51] = t[69] ^ x[10];
  assign t[52] = t[70] ^ x[9];
  assign t[53] = t[71] ^ x[13];
  assign t[54] = t[72] ^ x[12];
  assign t[55] = t[73] ^ x[16];
  assign t[56] = t[74] ^ x[15];
  assign t[57] = t[75] ^ x[19];
  assign t[58] = t[76] ^ x[18];
  assign t[59] = t[77] ^ x[22];
  assign t[5] = ~t[7];
  assign t[60] = t[78] ^ x[21];
  assign t[61] = t[79] ^ x[25];
  assign t[62] = t[80] ^ x[24];
  assign t[63] = t[81] ^ x[28];
  assign t[64] = t[82] ^ x[27];
  assign t[65] = t[83] ^ x[31];
  assign t[66] = t[84] ^ x[30];
  assign t[67] = (x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[8]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (x[8]);
  assign t[71] = (x[11]);
  assign t[72] = (x[11]);
  assign t[73] = (x[14]);
  assign t[74] = (x[14]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[20]);
  assign t[78] = (x[20]);
  assign t[79] = (x[23]);
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[80] = (x[23]);
  assign t[81] = (x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29]);
  assign t[84] = (x[29]);
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind101(x, y);
 input [31:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14] & t[15]);
  assign t[11] = t[16] | t[23];
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[24];
  assign t[14] = ~(t[25]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[20] | t[14]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[28]);
  assign t[19] = ~(t[21] | t[17]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29]);
  assign t[21] = ~(t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[39]);
  assign t[31] = t[40] ^ x[5];
  assign t[32] = t[41] ^ x[10];
  assign t[33] = t[42] ^ x[13];
  assign t[34] = t[43] ^ x[16];
  assign t[35] = t[44] ^ x[19];
  assign t[36] = t[45] ^ x[22];
  assign t[37] = t[46] ^ x[25];
  assign t[38] = t[47] ^ x[28];
  assign t[39] = t[48] ^ x[31];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[49] & ~t[50]);
  assign t[41] = (t[51] & ~t[52]);
  assign t[42] = (t[53] & ~t[54]);
  assign t[43] = (t[55] & ~t[56]);
  assign t[44] = (t[57] & ~t[58]);
  assign t[45] = (t[59] & ~t[60]);
  assign t[46] = (t[61] & ~t[62]);
  assign t[47] = (t[63] & ~t[64]);
  assign t[48] = (t[65] & ~t[66]);
  assign t[49] = t[67] ^ x[5];
  assign t[4] = ~x[2] & t[22];
  assign t[50] = t[68] ^ x[4];
  assign t[51] = t[69] ^ x[10];
  assign t[52] = t[70] ^ x[9];
  assign t[53] = t[71] ^ x[13];
  assign t[54] = t[72] ^ x[12];
  assign t[55] = t[73] ^ x[16];
  assign t[56] = t[74] ^ x[15];
  assign t[57] = t[75] ^ x[19];
  assign t[58] = t[76] ^ x[18];
  assign t[59] = t[77] ^ x[22];
  assign t[5] = ~t[7];
  assign t[60] = t[78] ^ x[21];
  assign t[61] = t[79] ^ x[25];
  assign t[62] = t[80] ^ x[24];
  assign t[63] = t[81] ^ x[28];
  assign t[64] = t[82] ^ x[27];
  assign t[65] = t[83] ^ x[31];
  assign t[66] = t[84] ^ x[30];
  assign t[67] = (x[3]);
  assign t[68] = (x[3]);
  assign t[69] = (x[8]);
  assign t[6] = x[2] ? x[6] : t[8];
  assign t[70] = (x[8]);
  assign t[71] = (x[11]);
  assign t[72] = (x[11]);
  assign t[73] = (x[14]);
  assign t[74] = (x[14]);
  assign t[75] = (x[17]);
  assign t[76] = (x[17]);
  assign t[77] = (x[20]);
  assign t[78] = (x[20]);
  assign t[79] = (x[23]);
  assign t[7] = x[2] ? x[7] : t[9];
  assign t[80] = (x[23]);
  assign t[81] = (x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29]);
  assign t[84] = (x[29]);
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[29] | t[20]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[31] | t[23]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~(~x[2] & ~t[28]);
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[29] | t[20]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[31] | t[23]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~(~x[2] & ~t[28]);
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [28:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~(t[26] & t[19]);
  assign t[15] = ~x[2] & t[27];
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29] & t[21]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[31] & t[23]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[28]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = t[47] ^ x[28];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = (t[48] & ~t[49]);
  assign t[41] = (t[50] & ~t[51]);
  assign t[42] = (t[52] & ~t[53]);
  assign t[43] = (t[54] & ~t[55]);
  assign t[44] = (t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[59]);
  assign t[46] = (t[60] & ~t[61]);
  assign t[47] = (t[62] & ~t[63]);
  assign t[48] = t[64] ^ x[5];
  assign t[49] = t[65] ^ x[4];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = t[66] ^ x[10];
  assign t[51] = t[67] ^ x[9];
  assign t[52] = t[68] ^ x[13];
  assign t[53] = t[69] ^ x[12];
  assign t[54] = t[70] ^ x[16];
  assign t[55] = t[71] ^ x[15];
  assign t[56] = t[72] ^ x[19];
  assign t[57] = t[73] ^ x[18];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[21];
  assign t[5] = ~x[2] & t[24];
  assign t[60] = t[76] ^ x[25];
  assign t[61] = t[77] ^ x[24];
  assign t[62] = t[78] ^ x[28];
  assign t[63] = t[79] ^ x[27];
  assign t[64] = (x[3]);
  assign t[65] = (x[3]);
  assign t[66] = (x[8]);
  assign t[67] = (x[8]);
  assign t[68] = (x[11]);
  assign t[69] = (x[11]);
  assign t[6] = ~t[9];
  assign t[70] = (x[14]);
  assign t[71] = (x[14]);
  assign t[72] = (x[17]);
  assign t[73] = (x[17]);
  assign t[74] = (x[20]);
  assign t[75] = (x[20]);
  assign t[76] = (x[23]);
  assign t[77] = (x[23]);
  assign t[78] = (x[26]);
  assign t[79] = (x[26]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [28:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~(t[26] & t[19]);
  assign t[15] = ~x[2] & t[27];
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29] & t[21]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[31] & t[23]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[28]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = t[47] ^ x[28];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = (t[48] & ~t[49]);
  assign t[41] = (t[50] & ~t[51]);
  assign t[42] = (t[52] & ~t[53]);
  assign t[43] = (t[54] & ~t[55]);
  assign t[44] = (t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[59]);
  assign t[46] = (t[60] & ~t[61]);
  assign t[47] = (t[62] & ~t[63]);
  assign t[48] = t[64] ^ x[5];
  assign t[49] = t[65] ^ x[4];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = t[66] ^ x[10];
  assign t[51] = t[67] ^ x[9];
  assign t[52] = t[68] ^ x[13];
  assign t[53] = t[69] ^ x[12];
  assign t[54] = t[70] ^ x[16];
  assign t[55] = t[71] ^ x[15];
  assign t[56] = t[72] ^ x[19];
  assign t[57] = t[73] ^ x[18];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[21];
  assign t[5] = ~x[2] & t[24];
  assign t[60] = t[76] ^ x[25];
  assign t[61] = t[77] ^ x[24];
  assign t[62] = t[78] ^ x[28];
  assign t[63] = t[79] ^ x[27];
  assign t[64] = (x[3]);
  assign t[65] = (x[3]);
  assign t[66] = (x[8]);
  assign t[67] = (x[8]);
  assign t[68] = (x[11]);
  assign t[69] = (x[11]);
  assign t[6] = ~t[9];
  assign t[70] = (x[14]);
  assign t[71] = (x[14]);
  assign t[72] = (x[17]);
  assign t[73] = (x[17]);
  assign t[74] = (x[20]);
  assign t[75] = (x[20]);
  assign t[76] = (x[23]);
  assign t[77] = (x[23]);
  assign t[78] = (x[26]);
  assign t[79] = (x[26]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind106(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[29]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[33] & t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] & t[34]);
  assign t[27] = ~(t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~x[2] & t[28];
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[29]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[33] & t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] & t[34]);
  assign t[27] = ~(t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~x[2] & t[28];
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [31:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[25];
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = t[22] | t[27];
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[23] | t[17]);
  assign t[1] = t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[24] | t[20]);
  assign t[23] = ~(t[32]);
  assign t[24] = ~(t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[10];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[16];
  assign t[38] = t[47] ^ x[19];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[25];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[31];
  assign t[43] = (t[52] & ~t[53]);
  assign t[44] = (t[54] & ~t[55]);
  assign t[45] = (t[56] & ~t[57]);
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = t[7] ? x[1] : x[0];
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = t[70] ^ x[7];
  assign t[53] = t[71] ^ x[6];
  assign t[54] = t[72] ^ x[10];
  assign t[55] = t[73] ^ x[9];
  assign t[56] = t[74] ^ x[13];
  assign t[57] = t[75] ^ x[12];
  assign t[58] = t[76] ^ x[16];
  assign t[59] = t[77] ^ x[15];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[19];
  assign t[61] = t[79] ^ x[18];
  assign t[62] = t[80] ^ x[22];
  assign t[63] = t[81] ^ x[21];
  assign t[64] = t[82] ^ x[25];
  assign t[65] = t[83] ^ x[24];
  assign t[66] = t[84] ^ x[28];
  assign t[67] = t[85] ^ x[27];
  assign t[68] = t[86] ^ x[31];
  assign t[69] = t[87] ^ x[30];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[5]);
  assign t[71] = (x[5]);
  assign t[72] = (x[8]);
  assign t[73] = (x[8]);
  assign t[74] = (x[11]);
  assign t[75] = (x[11]);
  assign t[76] = (x[14]);
  assign t[77] = (x[14]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[20]);
  assign t[81] = (x[20]);
  assign t[82] = (x[23]);
  assign t[83] = (x[23]);
  assign t[84] = (x[26]);
  assign t[85] = (x[26]);
  assign t[86] = (x[29]);
  assign t[87] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [31:0] x;
 output y;

 wire [87:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = t[19] | t[25];
  assign t[14] = ~x[2] & t[26];
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = t[22] | t[27];
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[29]);
  assign t[19] = ~(t[23] | t[17]);
  assign t[1] = t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31]);
  assign t[22] = ~(t[24] | t[20]);
  assign t[23] = ~(t[32]);
  assign t[24] = ~(t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = (t[37]);
  assign t[29] = (t[38]);
  assign t[2] = ~t[4];
  assign t[30] = (t[39]);
  assign t[31] = (t[40]);
  assign t[32] = (t[41]);
  assign t[33] = (t[42]);
  assign t[34] = t[43] ^ x[7];
  assign t[35] = t[44] ^ x[10];
  assign t[36] = t[45] ^ x[13];
  assign t[37] = t[46] ^ x[16];
  assign t[38] = t[47] ^ x[19];
  assign t[39] = t[48] ^ x[22];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[49] ^ x[25];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[31];
  assign t[43] = (t[52] & ~t[53]);
  assign t[44] = (t[54] & ~t[55]);
  assign t[45] = (t[56] & ~t[57]);
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = t[7] ? x[1] : x[0];
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = t[70] ^ x[7];
  assign t[53] = t[71] ^ x[6];
  assign t[54] = t[72] ^ x[10];
  assign t[55] = t[73] ^ x[9];
  assign t[56] = t[74] ^ x[13];
  assign t[57] = t[75] ^ x[12];
  assign t[58] = t[76] ^ x[16];
  assign t[59] = t[77] ^ x[15];
  assign t[5] = ~t[8];
  assign t[60] = t[78] ^ x[19];
  assign t[61] = t[79] ^ x[18];
  assign t[62] = t[80] ^ x[22];
  assign t[63] = t[81] ^ x[21];
  assign t[64] = t[82] ^ x[25];
  assign t[65] = t[83] ^ x[24];
  assign t[66] = t[84] ^ x[28];
  assign t[67] = t[85] ^ x[27];
  assign t[68] = t[86] ^ x[31];
  assign t[69] = t[87] ^ x[30];
  assign t[6] = x[2] ? x[3] : t[9];
  assign t[70] = (x[5]);
  assign t[71] = (x[5]);
  assign t[72] = (x[8]);
  assign t[73] = (x[8]);
  assign t[74] = (x[11]);
  assign t[75] = (x[11]);
  assign t[76] = (x[14]);
  assign t[77] = (x[14]);
  assign t[78] = (x[17]);
  assign t[79] = (x[17]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[20]);
  assign t[81] = (x[20]);
  assign t[82] = (x[23]);
  assign t[83] = (x[23]);
  assign t[84] = (x[26]);
  assign t[85] = (x[26]);
  assign t[86] = (x[29]);
  assign t[87] = (x[29]);
  assign t[8] = x[2] ? x[4] : t[11];
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[29] | t[20]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[31] | t[23]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~(~x[2] & ~t[28]);
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind111(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = ~(t[29] | t[20]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] | t[22]);
  assign t[17] = ~(t[31] | t[23]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[37]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~(~x[2] & ~t[28]);
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [28:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~(t[26] & t[19]);
  assign t[15] = ~x[2] & t[27];
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29] & t[21]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[31] & t[23]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[28]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = t[47] ^ x[28];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = (t[48] & ~t[49]);
  assign t[41] = (t[50] & ~t[51]);
  assign t[42] = (t[52] & ~t[53]);
  assign t[43] = (t[54] & ~t[55]);
  assign t[44] = (t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[59]);
  assign t[46] = (t[60] & ~t[61]);
  assign t[47] = (t[62] & ~t[63]);
  assign t[48] = t[64] ^ x[5];
  assign t[49] = t[65] ^ x[4];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = t[66] ^ x[10];
  assign t[51] = t[67] ^ x[9];
  assign t[52] = t[68] ^ x[13];
  assign t[53] = t[69] ^ x[12];
  assign t[54] = t[70] ^ x[16];
  assign t[55] = t[71] ^ x[15];
  assign t[56] = t[72] ^ x[19];
  assign t[57] = t[73] ^ x[18];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[21];
  assign t[5] = ~x[2] & t[24];
  assign t[60] = t[76] ^ x[25];
  assign t[61] = t[77] ^ x[24];
  assign t[62] = t[78] ^ x[28];
  assign t[63] = t[79] ^ x[27];
  assign t[64] = (x[3]);
  assign t[65] = (x[3]);
  assign t[66] = (x[8]);
  assign t[67] = (x[8]);
  assign t[68] = (x[11]);
  assign t[69] = (x[11]);
  assign t[6] = ~t[9];
  assign t[70] = (x[14]);
  assign t[71] = (x[14]);
  assign t[72] = (x[17]);
  assign t[73] = (x[17]);
  assign t[74] = (x[20]);
  assign t[75] = (x[20]);
  assign t[76] = (x[23]);
  assign t[77] = (x[23]);
  assign t[78] = (x[26]);
  assign t[79] = (x[26]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [28:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[25] & t[18]);
  assign t[14] = ~(t[26] & t[19]);
  assign t[15] = ~x[2] & t[27];
  assign t[16] = ~(t[28] & t[20]);
  assign t[17] = ~(t[29] & t[21]);
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = t[3];
  assign t[20] = ~(t[31]);
  assign t[21] = ~(t[31] & t[23]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[28]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[5];
  assign t[33] = t[41] ^ x[10];
  assign t[34] = t[42] ^ x[13];
  assign t[35] = t[43] ^ x[16];
  assign t[36] = t[44] ^ x[19];
  assign t[37] = t[45] ^ x[22];
  assign t[38] = t[46] ^ x[25];
  assign t[39] = t[47] ^ x[28];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = (t[48] & ~t[49]);
  assign t[41] = (t[50] & ~t[51]);
  assign t[42] = (t[52] & ~t[53]);
  assign t[43] = (t[54] & ~t[55]);
  assign t[44] = (t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[59]);
  assign t[46] = (t[60] & ~t[61]);
  assign t[47] = (t[62] & ~t[63]);
  assign t[48] = t[64] ^ x[5];
  assign t[49] = t[65] ^ x[4];
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = t[66] ^ x[10];
  assign t[51] = t[67] ^ x[9];
  assign t[52] = t[68] ^ x[13];
  assign t[53] = t[69] ^ x[12];
  assign t[54] = t[70] ^ x[16];
  assign t[55] = t[71] ^ x[15];
  assign t[56] = t[72] ^ x[19];
  assign t[57] = t[73] ^ x[18];
  assign t[58] = t[74] ^ x[22];
  assign t[59] = t[75] ^ x[21];
  assign t[5] = ~x[2] & t[24];
  assign t[60] = t[76] ^ x[25];
  assign t[61] = t[77] ^ x[24];
  assign t[62] = t[78] ^ x[28];
  assign t[63] = t[79] ^ x[27];
  assign t[64] = (x[3]);
  assign t[65] = (x[3]);
  assign t[66] = (x[8]);
  assign t[67] = (x[8]);
  assign t[68] = (x[11]);
  assign t[69] = (x[11]);
  assign t[6] = ~t[9];
  assign t[70] = (x[14]);
  assign t[71] = (x[14]);
  assign t[72] = (x[17]);
  assign t[73] = (x[17]);
  assign t[74] = (x[20]);
  assign t[75] = (x[20]);
  assign t[76] = (x[23]);
  assign t[77] = (x[23]);
  assign t[78] = (x[26]);
  assign t[79] = (x[26]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[29]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[33] & t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] & t[34]);
  assign t[27] = ~(t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~x[2] & t[28];
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [34:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[20] & t[29]);
  assign t[15] = ~x[2] & t[30];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[23] & t[31]);
  assign t[18] = ~(t[32]);
  assign t[19] = ~(t[33]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] & t[25]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[26] & t[27]);
  assign t[24] = ~(t[33] & t[32]);
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[35] & t[34]);
  assign t[27] = ~(t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[10];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[13];
  assign t[41] = t[51] ^ x[16];
  assign t[42] = t[52] ^ x[19];
  assign t[43] = t[53] ^ x[22];
  assign t[44] = t[54] ^ x[25];
  assign t[45] = t[55] ^ x[28];
  assign t[46] = t[56] ^ x[31];
  assign t[47] = t[57] ^ x[34];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = ~x[2] & t[28];
  assign t[60] = t[80] ^ x[10];
  assign t[61] = t[81] ^ x[9];
  assign t[62] = t[82] ^ x[13];
  assign t[63] = t[83] ^ x[12];
  assign t[64] = t[84] ^ x[16];
  assign t[65] = t[85] ^ x[15];
  assign t[66] = t[86] ^ x[19];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[22];
  assign t[69] = t[89] ^ x[21];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[25];
  assign t[71] = t[91] ^ x[24];
  assign t[72] = t[92] ^ x[28];
  assign t[73] = t[93] ^ x[27];
  assign t[74] = t[94] ^ x[31];
  assign t[75] = t[95] ^ x[30];
  assign t[76] = t[96] ^ x[34];
  assign t[77] = t[97] ^ x[33];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[8]);
  assign t[81] = (x[8]);
  assign t[82] = (x[11]);
  assign t[83] = (x[11]);
  assign t[84] = (x[14]);
  assign t[85] = (x[14]);
  assign t[86] = (x[17]);
  assign t[87] = (x[17]);
  assign t[88] = (x[20]);
  assign t[89] = (x[20]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[23]);
  assign t[91] = (x[23]);
  assign t[92] = (x[26]);
  assign t[93] = (x[26]);
  assign t[94] = (x[29]);
  assign t[95] = (x[29]);
  assign t[96] = (x[32]);
  assign t[97] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind116(x, y);
 input [34:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = t[20] | t[27];
  assign t[15] = ~x[2] & t[28];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = t[23] | t[29];
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[18]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[25] | t[21]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = t[46] ^ x[5];
  assign t[37] = t[47] ^ x[10];
  assign t[38] = t[48] ^ x[13];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[19];
  assign t[41] = t[51] ^ x[22];
  assign t[42] = t[52] ^ x[25];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[31];
  assign t[45] = t[55] ^ x[34];
  assign t[46] = (t[56] & ~t[57]);
  assign t[47] = (t[58] & ~t[59]);
  assign t[48] = (t[60] & ~t[61]);
  assign t[49] = (t[62] & ~t[63]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = t[76] ^ x[5];
  assign t[57] = t[77] ^ x[4];
  assign t[58] = t[78] ^ x[10];
  assign t[59] = t[79] ^ x[9];
  assign t[5] = ~x[2] & t[26];
  assign t[60] = t[80] ^ x[13];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[16];
  assign t[63] = t[83] ^ x[15];
  assign t[64] = t[84] ^ x[19];
  assign t[65] = t[85] ^ x[18];
  assign t[66] = t[86] ^ x[22];
  assign t[67] = t[87] ^ x[21];
  assign t[68] = t[88] ^ x[25];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[28];
  assign t[71] = t[91] ^ x[27];
  assign t[72] = t[92] ^ x[31];
  assign t[73] = t[93] ^ x[30];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[33];
  assign t[76] = (x[3]);
  assign t[77] = (x[3]);
  assign t[78] = (x[8]);
  assign t[79] = (x[8]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[11]);
  assign t[81] = (x[11]);
  assign t[82] = (x[14]);
  assign t[83] = (x[14]);
  assign t[84] = (x[17]);
  assign t[85] = (x[17]);
  assign t[86] = (x[20]);
  assign t[87] = (x[20]);
  assign t[88] = (x[23]);
  assign t[89] = (x[23]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[26]);
  assign t[91] = (x[26]);
  assign t[92] = (x[29]);
  assign t[93] = (x[29]);
  assign t[94] = (x[32]);
  assign t[95] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [34:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = t[20] | t[27];
  assign t[15] = ~x[2] & t[28];
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = t[23] | t[29];
  assign t[18] = ~(t[30]);
  assign t[19] = ~(t[31]);
  assign t[1] = t[3];
  assign t[20] = ~(t[24] | t[18]);
  assign t[21] = ~(t[32]);
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[25] | t[21]);
  assign t[24] = ~(t[34]);
  assign t[25] = ~(t[35]);
  assign t[26] = (t[36]);
  assign t[27] = (t[37]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = t[46] ^ x[5];
  assign t[37] = t[47] ^ x[10];
  assign t[38] = t[48] ^ x[13];
  assign t[39] = t[49] ^ x[16];
  assign t[3] = ~(t[6] ^ t[7]);
  assign t[40] = t[50] ^ x[19];
  assign t[41] = t[51] ^ x[22];
  assign t[42] = t[52] ^ x[25];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[31];
  assign t[45] = t[55] ^ x[34];
  assign t[46] = (t[56] & ~t[57]);
  assign t[47] = (t[58] & ~t[59]);
  assign t[48] = (t[60] & ~t[61]);
  assign t[49] = (t[62] & ~t[63]);
  assign t[4] = t[8] ? x[1] : x[0];
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = t[76] ^ x[5];
  assign t[57] = t[77] ^ x[4];
  assign t[58] = t[78] ^ x[10];
  assign t[59] = t[79] ^ x[9];
  assign t[5] = ~x[2] & t[26];
  assign t[60] = t[80] ^ x[13];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[16];
  assign t[63] = t[83] ^ x[15];
  assign t[64] = t[84] ^ x[19];
  assign t[65] = t[85] ^ x[18];
  assign t[66] = t[86] ^ x[22];
  assign t[67] = t[87] ^ x[21];
  assign t[68] = t[88] ^ x[25];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~t[9];
  assign t[70] = t[90] ^ x[28];
  assign t[71] = t[91] ^ x[27];
  assign t[72] = t[92] ^ x[31];
  assign t[73] = t[93] ^ x[30];
  assign t[74] = t[94] ^ x[34];
  assign t[75] = t[95] ^ x[33];
  assign t[76] = (x[3]);
  assign t[77] = (x[3]);
  assign t[78] = (x[8]);
  assign t[79] = (x[8]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[11]);
  assign t[81] = (x[11]);
  assign t[82] = (x[14]);
  assign t[83] = (x[14]);
  assign t[84] = (x[17]);
  assign t[85] = (x[17]);
  assign t[86] = (x[20]);
  assign t[87] = (x[20]);
  assign t[88] = (x[23]);
  assign t[89] = (x[23]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[26]);
  assign t[91] = (x[26]);
  assign t[92] = (x[29]);
  assign t[93] = (x[29]);
  assign t[94] = (x[32]);
  assign t[95] = (x[32]);
  assign t[9] = x[2] ? x[7] : t[12];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[11];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[17];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[23];
  assign t[46] = t[56] ^ x[26];
  assign t[47] = t[57] ^ x[29];
  assign t[48] = t[58] ^ x[32];
  assign t[49] = t[59] ^ x[35];
  assign t[4] = ~(t[7]);
  assign t[50] = (t[60] & ~t[61]);
  assign t[51] = (t[62] & ~t[63]);
  assign t[52] = (t[64] & ~t[65]);
  assign t[53] = (t[66] & ~t[67]);
  assign t[54] = (t[68] & ~t[69]);
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[11];
  assign t[63] = t[83] ^ x[10];
  assign t[64] = t[84] ^ x[14];
  assign t[65] = t[85] ^ x[13];
  assign t[66] = t[86] ^ x[17];
  assign t[67] = t[87] ^ x[16];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[23];
  assign t[71] = t[91] ^ x[22];
  assign t[72] = t[92] ^ x[26];
  assign t[73] = t[93] ^ x[25];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[28];
  assign t[76] = t[96] ^ x[32];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[35];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = ~(t[11]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind121(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[11];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[17];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[23];
  assign t[46] = t[56] ^ x[26];
  assign t[47] = t[57] ^ x[29];
  assign t[48] = t[58] ^ x[32];
  assign t[49] = t[59] ^ x[35];
  assign t[4] = ~(t[7]);
  assign t[50] = (t[60] & ~t[61]);
  assign t[51] = (t[62] & ~t[63]);
  assign t[52] = (t[64] & ~t[65]);
  assign t[53] = (t[66] & ~t[67]);
  assign t[54] = (t[68] & ~t[69]);
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[11];
  assign t[63] = t[83] ^ x[10];
  assign t[64] = t[84] ^ x[14];
  assign t[65] = t[85] ^ x[13];
  assign t[66] = t[86] ^ x[17];
  assign t[67] = t[87] ^ x[16];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[23];
  assign t[71] = t[91] ^ x[22];
  assign t[72] = t[92] ^ x[26];
  assign t[73] = t[93] ^ x[25];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[28];
  assign t[76] = t[96] ^ x[32];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[35];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = ~(t[11]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[38]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[45] & t[44]);
  assign t[35] = ~(t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[38]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[45] & t[44]);
  assign t[35] = ~(t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [44:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[9]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[15]);
  assign t[105] = (x[15]);
  assign t[106] = (x[18]);
  assign t[107] = (x[18]);
  assign t[108] = (x[21]);
  assign t[109] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[24]);
  assign t[111] = (x[24]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[30]);
  assign t[115] = (x[30]);
  assign t[116] = (x[33]);
  assign t[117] = (x[33]);
  assign t[118] = (x[36]);
  assign t[119] = (x[36]);
  assign t[11] = ~x[2] & t[33];
  assign t[120] = (x[39]);
  assign t[121] = (x[39]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[17];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[20];
  assign t[51] = t[64] ^ x[23];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[32];
  assign t[55] = t[68] ^ x[35];
  assign t[56] = t[69] ^ x[38];
  assign t[57] = t[70] ^ x[41];
  assign t[58] = t[71] ^ x[44];
  assign t[59] = (t[72] & ~t[73]);
  assign t[5] = t[8];
  assign t[60] = (t[74] & ~t[75]);
  assign t[61] = (t[76] & ~t[77]);
  assign t[62] = (t[78] & ~t[79]);
  assign t[63] = (t[80] & ~t[81]);
  assign t[64] = (t[82] & ~t[83]);
  assign t[65] = (t[84] & ~t[85]);
  assign t[66] = (t[86] & ~t[87]);
  assign t[67] = (t[88] & ~t[89]);
  assign t[68] = (t[90] & ~t[91]);
  assign t[69] = (t[92] & ~t[93]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[94] & ~t[95]);
  assign t[71] = (t[96] & ~t[97]);
  assign t[72] = t[98] ^ x[8];
  assign t[73] = t[99] ^ x[7];
  assign t[74] = t[100] ^ x[11];
  assign t[75] = t[101] ^ x[10];
  assign t[76] = t[102] ^ x[14];
  assign t[77] = t[103] ^ x[13];
  assign t[78] = t[104] ^ x[17];
  assign t[79] = t[105] ^ x[16];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[20];
  assign t[81] = t[107] ^ x[19];
  assign t[82] = t[108] ^ x[23];
  assign t[83] = t[109] ^ x[22];
  assign t[84] = t[110] ^ x[26];
  assign t[85] = t[111] ^ x[25];
  assign t[86] = t[112] ^ x[29];
  assign t[87] = t[113] ^ x[28];
  assign t[88] = t[114] ^ x[32];
  assign t[89] = t[115] ^ x[31];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[35];
  assign t[91] = t[117] ^ x[34];
  assign t[92] = t[118] ^ x[38];
  assign t[93] = t[119] ^ x[37];
  assign t[94] = t[120] ^ x[41];
  assign t[95] = t[121] ^ x[40];
  assign t[96] = t[122] ^ x[44];
  assign t[97] = t[123] ^ x[43];
  assign t[98] = (x[6]);
  assign t[99] = (x[6]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [44:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[9]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[15]);
  assign t[105] = (x[15]);
  assign t[106] = (x[18]);
  assign t[107] = (x[18]);
  assign t[108] = (x[21]);
  assign t[109] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[24]);
  assign t[111] = (x[24]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[30]);
  assign t[115] = (x[30]);
  assign t[116] = (x[33]);
  assign t[117] = (x[33]);
  assign t[118] = (x[36]);
  assign t[119] = (x[36]);
  assign t[11] = ~x[2] & t[33];
  assign t[120] = (x[39]);
  assign t[121] = (x[39]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[17];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[20];
  assign t[51] = t[64] ^ x[23];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[32];
  assign t[55] = t[68] ^ x[35];
  assign t[56] = t[69] ^ x[38];
  assign t[57] = t[70] ^ x[41];
  assign t[58] = t[71] ^ x[44];
  assign t[59] = (t[72] & ~t[73]);
  assign t[5] = t[8];
  assign t[60] = (t[74] & ~t[75]);
  assign t[61] = (t[76] & ~t[77]);
  assign t[62] = (t[78] & ~t[79]);
  assign t[63] = (t[80] & ~t[81]);
  assign t[64] = (t[82] & ~t[83]);
  assign t[65] = (t[84] & ~t[85]);
  assign t[66] = (t[86] & ~t[87]);
  assign t[67] = (t[88] & ~t[89]);
  assign t[68] = (t[90] & ~t[91]);
  assign t[69] = (t[92] & ~t[93]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[94] & ~t[95]);
  assign t[71] = (t[96] & ~t[97]);
  assign t[72] = t[98] ^ x[8];
  assign t[73] = t[99] ^ x[7];
  assign t[74] = t[100] ^ x[11];
  assign t[75] = t[101] ^ x[10];
  assign t[76] = t[102] ^ x[14];
  assign t[77] = t[103] ^ x[13];
  assign t[78] = t[104] ^ x[17];
  assign t[79] = t[105] ^ x[16];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[20];
  assign t[81] = t[107] ^ x[19];
  assign t[82] = t[108] ^ x[23];
  assign t[83] = t[109] ^ x[22];
  assign t[84] = t[110] ^ x[26];
  assign t[85] = t[111] ^ x[25];
  assign t[86] = t[112] ^ x[29];
  assign t[87] = t[113] ^ x[28];
  assign t[88] = t[114] ^ x[32];
  assign t[89] = t[115] ^ x[31];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[35];
  assign t[91] = t[117] ^ x[34];
  assign t[92] = t[118] ^ x[38];
  assign t[93] = t[119] ^ x[37];
  assign t[94] = t[120] ^ x[41];
  assign t[95] = t[121] ^ x[40];
  assign t[96] = t[122] ^ x[44];
  assign t[97] = t[123] ^ x[43];
  assign t[98] = (x[6]);
  assign t[99] = (x[6]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind126(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [35:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[29] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[35] & t[25]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[36] & t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = ~(t[37] & t[27]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[31]);
  assign t[27] = ~(t[33]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[11];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[14];
  assign t[41] = t[51] ^ x[17];
  assign t[42] = t[52] ^ x[20];
  assign t[43] = t[53] ^ x[23];
  assign t[44] = t[54] ^ x[26];
  assign t[45] = t[55] ^ x[29];
  assign t[46] = t[56] ^ x[32];
  assign t[47] = t[57] ^ x[35];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = ~x[2] & t[28];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = t[7];
  assign t[60] = t[80] ^ x[11];
  assign t[61] = t[81] ^ x[10];
  assign t[62] = t[82] ^ x[14];
  assign t[63] = t[83] ^ x[13];
  assign t[64] = t[84] ^ x[17];
  assign t[65] = t[85] ^ x[16];
  assign t[66] = t[86] ^ x[20];
  assign t[67] = t[87] ^ x[19];
  assign t[68] = t[88] ^ x[23];
  assign t[69] = t[89] ^ x[22];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[26];
  assign t[71] = t[91] ^ x[25];
  assign t[72] = t[92] ^ x[29];
  assign t[73] = t[93] ^ x[28];
  assign t[74] = t[94] ^ x[32];
  assign t[75] = t[95] ^ x[31];
  assign t[76] = t[96] ^ x[35];
  assign t[77] = t[97] ^ x[34];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[9]);
  assign t[81] = (x[9]);
  assign t[82] = (x[12]);
  assign t[83] = (x[12]);
  assign t[84] = (x[15]);
  assign t[85] = (x[15]);
  assign t[86] = (x[18]);
  assign t[87] = (x[18]);
  assign t[88] = (x[21]);
  assign t[89] = (x[21]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = (x[24]);
  assign t[91] = (x[24]);
  assign t[92] = (x[27]);
  assign t[93] = (x[27]);
  assign t[94] = (x[30]);
  assign t[95] = (x[30]);
  assign t[96] = (x[33]);
  assign t[97] = (x[33]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [35:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[29] & t[19]);
  assign t[14] = ~(t[30] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[35] & t[25]);
  assign t[21] = ~(t[36]);
  assign t[22] = ~(t[36] & t[26]);
  assign t[23] = ~(t[37]);
  assign t[24] = ~(t[37] & t[27]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[31]);
  assign t[27] = ~(t[33]);
  assign t[28] = (t[38]);
  assign t[29] = (t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = t[48] ^ x[5];
  assign t[39] = t[49] ^ x[11];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[14];
  assign t[41] = t[51] ^ x[17];
  assign t[42] = t[52] ^ x[20];
  assign t[43] = t[53] ^ x[23];
  assign t[44] = t[54] ^ x[26];
  assign t[45] = t[55] ^ x[29];
  assign t[46] = t[56] ^ x[32];
  assign t[47] = t[57] ^ x[35];
  assign t[48] = (t[58] & ~t[59]);
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = ~x[2] & t[28];
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = t[78] ^ x[5];
  assign t[59] = t[79] ^ x[4];
  assign t[5] = t[7];
  assign t[60] = t[80] ^ x[11];
  assign t[61] = t[81] ^ x[10];
  assign t[62] = t[82] ^ x[14];
  assign t[63] = t[83] ^ x[13];
  assign t[64] = t[84] ^ x[17];
  assign t[65] = t[85] ^ x[16];
  assign t[66] = t[86] ^ x[20];
  assign t[67] = t[87] ^ x[19];
  assign t[68] = t[88] ^ x[23];
  assign t[69] = t[89] ^ x[22];
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[90] ^ x[26];
  assign t[71] = t[91] ^ x[25];
  assign t[72] = t[92] ^ x[29];
  assign t[73] = t[93] ^ x[28];
  assign t[74] = t[94] ^ x[32];
  assign t[75] = t[95] ^ x[31];
  assign t[76] = t[96] ^ x[35];
  assign t[77] = t[97] ^ x[34];
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = (x[9]);
  assign t[81] = (x[9]);
  assign t[82] = (x[12]);
  assign t[83] = (x[12]);
  assign t[84] = (x[15]);
  assign t[85] = (x[15]);
  assign t[86] = (x[18]);
  assign t[87] = (x[18]);
  assign t[88] = (x[21]);
  assign t[89] = (x[21]);
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = (x[24]);
  assign t[91] = (x[24]);
  assign t[92] = (x[27]);
  assign t[93] = (x[27]);
  assign t[94] = (x[30]);
  assign t[95] = (x[30]);
  assign t[96] = (x[33]);
  assign t[97] = (x[33]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [44:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = ~(t[21] & t[35]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[36]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[39] & t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[11];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[17];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[23];
  assign t[53] = t[66] ^ x[26];
  assign t[54] = t[67] ^ x[29];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = t[70] ^ x[38];
  assign t[58] = t[71] ^ x[41];
  assign t[59] = t[72] ^ x[44];
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]);
  assign t[61] = (t[75] & ~t[76]);
  assign t[62] = (t[77] & ~t[78]);
  assign t[63] = (t[79] & ~t[80]);
  assign t[64] = (t[81] & ~t[82]);
  assign t[65] = (t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[86]);
  assign t[67] = (t[87] & ~t[88]);
  assign t[68] = (t[89] & ~t[90]);
  assign t[69] = (t[91] & ~t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[93] & ~t[94]);
  assign t[71] = (t[95] & ~t[96]);
  assign t[72] = (t[97] & ~t[98]);
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[4];
  assign t[75] = t[101] ^ x[11];
  assign t[76] = t[102] ^ x[10];
  assign t[77] = t[103] ^ x[14];
  assign t[78] = t[104] ^ x[13];
  assign t[79] = t[105] ^ x[17];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[16];
  assign t[81] = t[107] ^ x[20];
  assign t[82] = t[108] ^ x[19];
  assign t[83] = t[109] ^ x[23];
  assign t[84] = t[110] ^ x[22];
  assign t[85] = t[111] ^ x[26];
  assign t[86] = t[112] ^ x[25];
  assign t[87] = t[113] ^ x[29];
  assign t[88] = t[114] ^ x[28];
  assign t[89] = t[115] ^ x[32];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[31];
  assign t[91] = t[117] ^ x[35];
  assign t[92] = t[118] ^ x[34];
  assign t[93] = t[119] ^ x[38];
  assign t[94] = t[120] ^ x[37];
  assign t[95] = t[121] ^ x[41];
  assign t[96] = t[122] ^ x[40];
  assign t[97] = t[123] ^ x[44];
  assign t[98] = t[124] ^ x[43];
  assign t[99] = (x[3]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind131(x, y);
 input [44:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = ~(t[21] & t[35]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[36]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[39] & t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[11];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[17];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[23];
  assign t[53] = t[66] ^ x[26];
  assign t[54] = t[67] ^ x[29];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = t[70] ^ x[38];
  assign t[58] = t[71] ^ x[41];
  assign t[59] = t[72] ^ x[44];
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]);
  assign t[61] = (t[75] & ~t[76]);
  assign t[62] = (t[77] & ~t[78]);
  assign t[63] = (t[79] & ~t[80]);
  assign t[64] = (t[81] & ~t[82]);
  assign t[65] = (t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[86]);
  assign t[67] = (t[87] & ~t[88]);
  assign t[68] = (t[89] & ~t[90]);
  assign t[69] = (t[91] & ~t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[93] & ~t[94]);
  assign t[71] = (t[95] & ~t[96]);
  assign t[72] = (t[97] & ~t[98]);
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[4];
  assign t[75] = t[101] ^ x[11];
  assign t[76] = t[102] ^ x[10];
  assign t[77] = t[103] ^ x[14];
  assign t[78] = t[104] ^ x[13];
  assign t[79] = t[105] ^ x[17];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[16];
  assign t[81] = t[107] ^ x[20];
  assign t[82] = t[108] ^ x[19];
  assign t[83] = t[109] ^ x[23];
  assign t[84] = t[110] ^ x[22];
  assign t[85] = t[111] ^ x[26];
  assign t[86] = t[112] ^ x[25];
  assign t[87] = t[113] ^ x[29];
  assign t[88] = t[114] ^ x[28];
  assign t[89] = t[115] ^ x[32];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[31];
  assign t[91] = t[117] ^ x[35];
  assign t[92] = t[118] ^ x[34];
  assign t[93] = t[119] ^ x[38];
  assign t[94] = t[120] ^ x[37];
  assign t[95] = t[121] ^ x[41];
  assign t[96] = t[122] ^ x[40];
  assign t[97] = t[123] ^ x[44];
  assign t[98] = t[124] ^ x[43];
  assign t[99] = (x[3]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [44:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[9]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[15]);
  assign t[105] = (x[15]);
  assign t[106] = (x[18]);
  assign t[107] = (x[18]);
  assign t[108] = (x[21]);
  assign t[109] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[24]);
  assign t[111] = (x[24]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[30]);
  assign t[115] = (x[30]);
  assign t[116] = (x[33]);
  assign t[117] = (x[33]);
  assign t[118] = (x[36]);
  assign t[119] = (x[36]);
  assign t[11] = ~x[2] & t[33];
  assign t[120] = (x[39]);
  assign t[121] = (x[39]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[17];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[20];
  assign t[51] = t[64] ^ x[23];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[32];
  assign t[55] = t[68] ^ x[35];
  assign t[56] = t[69] ^ x[38];
  assign t[57] = t[70] ^ x[41];
  assign t[58] = t[71] ^ x[44];
  assign t[59] = (t[72] & ~t[73]);
  assign t[5] = t[8];
  assign t[60] = (t[74] & ~t[75]);
  assign t[61] = (t[76] & ~t[77]);
  assign t[62] = (t[78] & ~t[79]);
  assign t[63] = (t[80] & ~t[81]);
  assign t[64] = (t[82] & ~t[83]);
  assign t[65] = (t[84] & ~t[85]);
  assign t[66] = (t[86] & ~t[87]);
  assign t[67] = (t[88] & ~t[89]);
  assign t[68] = (t[90] & ~t[91]);
  assign t[69] = (t[92] & ~t[93]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[94] & ~t[95]);
  assign t[71] = (t[96] & ~t[97]);
  assign t[72] = t[98] ^ x[8];
  assign t[73] = t[99] ^ x[7];
  assign t[74] = t[100] ^ x[11];
  assign t[75] = t[101] ^ x[10];
  assign t[76] = t[102] ^ x[14];
  assign t[77] = t[103] ^ x[13];
  assign t[78] = t[104] ^ x[17];
  assign t[79] = t[105] ^ x[16];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[20];
  assign t[81] = t[107] ^ x[19];
  assign t[82] = t[108] ^ x[23];
  assign t[83] = t[109] ^ x[22];
  assign t[84] = t[110] ^ x[26];
  assign t[85] = t[111] ^ x[25];
  assign t[86] = t[112] ^ x[29];
  assign t[87] = t[113] ^ x[28];
  assign t[88] = t[114] ^ x[32];
  assign t[89] = t[115] ^ x[31];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[35];
  assign t[91] = t[117] ^ x[34];
  assign t[92] = t[118] ^ x[38];
  assign t[93] = t[119] ^ x[37];
  assign t[94] = t[120] ^ x[41];
  assign t[95] = t[121] ^ x[40];
  assign t[96] = t[122] ^ x[44];
  assign t[97] = t[123] ^ x[43];
  assign t[98] = (x[6]);
  assign t[99] = (x[6]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [44:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[9]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[15]);
  assign t[105] = (x[15]);
  assign t[106] = (x[18]);
  assign t[107] = (x[18]);
  assign t[108] = (x[21]);
  assign t[109] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[24]);
  assign t[111] = (x[24]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[30]);
  assign t[115] = (x[30]);
  assign t[116] = (x[33]);
  assign t[117] = (x[33]);
  assign t[118] = (x[36]);
  assign t[119] = (x[36]);
  assign t[11] = ~x[2] & t[33];
  assign t[120] = (x[39]);
  assign t[121] = (x[39]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[17];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[20];
  assign t[51] = t[64] ^ x[23];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[32];
  assign t[55] = t[68] ^ x[35];
  assign t[56] = t[69] ^ x[38];
  assign t[57] = t[70] ^ x[41];
  assign t[58] = t[71] ^ x[44];
  assign t[59] = (t[72] & ~t[73]);
  assign t[5] = t[8];
  assign t[60] = (t[74] & ~t[75]);
  assign t[61] = (t[76] & ~t[77]);
  assign t[62] = (t[78] & ~t[79]);
  assign t[63] = (t[80] & ~t[81]);
  assign t[64] = (t[82] & ~t[83]);
  assign t[65] = (t[84] & ~t[85]);
  assign t[66] = (t[86] & ~t[87]);
  assign t[67] = (t[88] & ~t[89]);
  assign t[68] = (t[90] & ~t[91]);
  assign t[69] = (t[92] & ~t[93]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[94] & ~t[95]);
  assign t[71] = (t[96] & ~t[97]);
  assign t[72] = t[98] ^ x[8];
  assign t[73] = t[99] ^ x[7];
  assign t[74] = t[100] ^ x[11];
  assign t[75] = t[101] ^ x[10];
  assign t[76] = t[102] ^ x[14];
  assign t[77] = t[103] ^ x[13];
  assign t[78] = t[104] ^ x[17];
  assign t[79] = t[105] ^ x[16];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[20];
  assign t[81] = t[107] ^ x[19];
  assign t[82] = t[108] ^ x[23];
  assign t[83] = t[109] ^ x[22];
  assign t[84] = t[110] ^ x[26];
  assign t[85] = t[111] ^ x[25];
  assign t[86] = t[112] ^ x[29];
  assign t[87] = t[113] ^ x[28];
  assign t[88] = t[114] ^ x[32];
  assign t[89] = t[115] ^ x[31];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[35];
  assign t[91] = t[117] ^ x[34];
  assign t[92] = t[118] ^ x[38];
  assign t[93] = t[119] ^ x[37];
  assign t[94] = t[120] ^ x[41];
  assign t[95] = t[121] ^ x[40];
  assign t[96] = t[122] ^ x[44];
  assign t[97] = t[123] ^ x[43];
  assign t[98] = (x[6]);
  assign t[99] = (x[6]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [44:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[14] = ~(t[35] | t[21]);
  assign t[15] = ~(t[22] | t[23]);
  assign t[16] = ~(t[36] | t[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[18] = ~(t[37] | t[27]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[44]);
  assign t[29] = ~(t[38] | t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[11];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[17];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[23];
  assign t[53] = t[66] ^ x[26];
  assign t[54] = t[67] ^ x[29];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = t[70] ^ x[38];
  assign t[58] = t[71] ^ x[41];
  assign t[59] = t[72] ^ x[44];
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]);
  assign t[61] = (t[75] & ~t[76]);
  assign t[62] = (t[77] & ~t[78]);
  assign t[63] = (t[79] & ~t[80]);
  assign t[64] = (t[81] & ~t[82]);
  assign t[65] = (t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[86]);
  assign t[67] = (t[87] & ~t[88]);
  assign t[68] = (t[89] & ~t[90]);
  assign t[69] = (t[91] & ~t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[93] & ~t[94]);
  assign t[71] = (t[95] & ~t[96]);
  assign t[72] = (t[97] & ~t[98]);
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[4];
  assign t[75] = t[101] ^ x[11];
  assign t[76] = t[102] ^ x[10];
  assign t[77] = t[103] ^ x[14];
  assign t[78] = t[104] ^ x[13];
  assign t[79] = t[105] ^ x[17];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[16];
  assign t[81] = t[107] ^ x[20];
  assign t[82] = t[108] ^ x[19];
  assign t[83] = t[109] ^ x[23];
  assign t[84] = t[110] ^ x[22];
  assign t[85] = t[111] ^ x[26];
  assign t[86] = t[112] ^ x[25];
  assign t[87] = t[113] ^ x[29];
  assign t[88] = t[114] ^ x[28];
  assign t[89] = t[115] ^ x[32];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[31];
  assign t[91] = t[117] ^ x[35];
  assign t[92] = t[118] ^ x[34];
  assign t[93] = t[119] ^ x[38];
  assign t[94] = t[120] ^ x[37];
  assign t[95] = t[121] ^ x[41];
  assign t[96] = t[122] ^ x[40];
  assign t[97] = t[123] ^ x[44];
  assign t[98] = t[124] ^ x[43];
  assign t[99] = (x[3]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [44:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[13] | t[14]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[14] = ~(t[35] | t[21]);
  assign t[15] = ~(t[22] | t[23]);
  assign t[16] = ~(t[36] | t[24]);
  assign t[17] = ~(t[25] | t[26]);
  assign t[18] = ~(t[37] | t[27]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] | t[33]);
  assign t[28] = ~(t[44]);
  assign t[29] = ~(t[38] | t[39]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[46]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[11];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[17];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[23];
  assign t[53] = t[66] ^ x[26];
  assign t[54] = t[67] ^ x[29];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = t[70] ^ x[38];
  assign t[58] = t[71] ^ x[41];
  assign t[59] = t[72] ^ x[44];
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]);
  assign t[61] = (t[75] & ~t[76]);
  assign t[62] = (t[77] & ~t[78]);
  assign t[63] = (t[79] & ~t[80]);
  assign t[64] = (t[81] & ~t[82]);
  assign t[65] = (t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[86]);
  assign t[67] = (t[87] & ~t[88]);
  assign t[68] = (t[89] & ~t[90]);
  assign t[69] = (t[91] & ~t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[93] & ~t[94]);
  assign t[71] = (t[95] & ~t[96]);
  assign t[72] = (t[97] & ~t[98]);
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[4];
  assign t[75] = t[101] ^ x[11];
  assign t[76] = t[102] ^ x[10];
  assign t[77] = t[103] ^ x[14];
  assign t[78] = t[104] ^ x[13];
  assign t[79] = t[105] ^ x[17];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[16];
  assign t[81] = t[107] ^ x[20];
  assign t[82] = t[108] ^ x[19];
  assign t[83] = t[109] ^ x[23];
  assign t[84] = t[110] ^ x[22];
  assign t[85] = t[111] ^ x[26];
  assign t[86] = t[112] ^ x[25];
  assign t[87] = t[113] ^ x[29];
  assign t[88] = t[114] ^ x[28];
  assign t[89] = t[115] ^ x[32];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[31];
  assign t[91] = t[117] ^ x[35];
  assign t[92] = t[118] ^ x[34];
  assign t[93] = t[119] ^ x[38];
  assign t[94] = t[120] ^ x[37];
  assign t[95] = t[121] ^ x[41];
  assign t[96] = t[122] ^ x[40];
  assign t[97] = t[123] ^ x[44];
  assign t[98] = t[124] ^ x[43];
  assign t[99] = (x[3]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind136(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[11];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[17];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[23];
  assign t[46] = t[56] ^ x[26];
  assign t[47] = t[57] ^ x[29];
  assign t[48] = t[58] ^ x[32];
  assign t[49] = t[59] ^ x[35];
  assign t[4] = ~(t[7]);
  assign t[50] = (t[60] & ~t[61]);
  assign t[51] = (t[62] & ~t[63]);
  assign t[52] = (t[64] & ~t[65]);
  assign t[53] = (t[66] & ~t[67]);
  assign t[54] = (t[68] & ~t[69]);
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[11];
  assign t[63] = t[83] ^ x[10];
  assign t[64] = t[84] ^ x[14];
  assign t[65] = t[85] ^ x[13];
  assign t[66] = t[86] ^ x[17];
  assign t[67] = t[87] ^ x[16];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[23];
  assign t[71] = t[91] ^ x[22];
  assign t[72] = t[92] ^ x[26];
  assign t[73] = t[93] ^ x[25];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[28];
  assign t[76] = t[96] ^ x[32];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[35];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = ~(t[11]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[11];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[17];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[23];
  assign t[46] = t[56] ^ x[26];
  assign t[47] = t[57] ^ x[29];
  assign t[48] = t[58] ^ x[32];
  assign t[49] = t[59] ^ x[35];
  assign t[4] = ~(t[7]);
  assign t[50] = (t[60] & ~t[61]);
  assign t[51] = (t[62] & ~t[63]);
  assign t[52] = (t[64] & ~t[65]);
  assign t[53] = (t[66] & ~t[67]);
  assign t[54] = (t[68] & ~t[69]);
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[11];
  assign t[63] = t[83] ^ x[10];
  assign t[64] = t[84] ^ x[14];
  assign t[65] = t[85] ^ x[13];
  assign t[66] = t[86] ^ x[17];
  assign t[67] = t[87] ^ x[16];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[23];
  assign t[71] = t[91] ^ x[22];
  assign t[72] = t[92] ^ x[26];
  assign t[73] = t[93] ^ x[25];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[28];
  assign t[76] = t[96] ^ x[32];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[35];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = ~(t[11]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[38]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[45] & t[44]);
  assign t[35] = ~(t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[38]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[29] & t[39]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] & t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] & t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[47]);
  assign t[34] = ~(t[45] & t[44]);
  assign t[35] = ~(t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [44:0] x;
 output y;

 wire [121:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = t[21] | t[32];
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = t[24] | t[33];
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] | t[34];
  assign t[19] = ~(t[35]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[28] | t[19]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] | t[22]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[30] | t[25]);
  assign t[28] = ~(t[41]);
  assign t[29] = ~(t[42]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = t[57] ^ x[5];
  assign t[45] = t[58] ^ x[11];
  assign t[46] = t[59] ^ x[14];
  assign t[47] = t[60] ^ x[17];
  assign t[48] = t[61] ^ x[20];
  assign t[49] = t[62] ^ x[23];
  assign t[4] = ~x[2] & t[31];
  assign t[50] = t[63] ^ x[26];
  assign t[51] = t[64] ^ x[29];
  assign t[52] = t[65] ^ x[32];
  assign t[53] = t[66] ^ x[35];
  assign t[54] = t[67] ^ x[38];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[44];
  assign t[57] = (t[70] & ~t[71]);
  assign t[58] = (t[72] & ~t[73]);
  assign t[59] = (t[74] & ~t[75]);
  assign t[5] = t[7];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[96] ^ x[5];
  assign t[71] = t[97] ^ x[4];
  assign t[72] = t[98] ^ x[11];
  assign t[73] = t[99] ^ x[10];
  assign t[74] = t[100] ^ x[14];
  assign t[75] = t[101] ^ x[13];
  assign t[76] = t[102] ^ x[17];
  assign t[77] = t[103] ^ x[16];
  assign t[78] = t[104] ^ x[20];
  assign t[79] = t[105] ^ x[19];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[23];
  assign t[81] = t[107] ^ x[22];
  assign t[82] = t[108] ^ x[26];
  assign t[83] = t[109] ^ x[25];
  assign t[84] = t[110] ^ x[29];
  assign t[85] = t[111] ^ x[28];
  assign t[86] = t[112] ^ x[32];
  assign t[87] = t[113] ^ x[31];
  assign t[88] = t[114] ^ x[35];
  assign t[89] = t[115] ^ x[34];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[38];
  assign t[91] = t[117] ^ x[37];
  assign t[92] = t[118] ^ x[41];
  assign t[93] = t[119] ^ x[40];
  assign t[94] = t[120] ^ x[44];
  assign t[95] = t[121] ^ x[43];
  assign t[96] = (x[3]);
  assign t[97] = (x[3]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind141(x, y);
 input [44:0] x;
 output y;

 wire [121:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = (x[42]);
  assign t[121] = (x[42]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = t[21] | t[32];
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = t[24] | t[33];
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] | t[34];
  assign t[19] = ~(t[35]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[28] | t[19]);
  assign t[22] = ~(t[37]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[29] | t[22]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = ~(t[30] | t[25]);
  assign t[28] = ~(t[41]);
  assign t[29] = ~(t[42]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = t[57] ^ x[5];
  assign t[45] = t[58] ^ x[11];
  assign t[46] = t[59] ^ x[14];
  assign t[47] = t[60] ^ x[17];
  assign t[48] = t[61] ^ x[20];
  assign t[49] = t[62] ^ x[23];
  assign t[4] = ~x[2] & t[31];
  assign t[50] = t[63] ^ x[26];
  assign t[51] = t[64] ^ x[29];
  assign t[52] = t[65] ^ x[32];
  assign t[53] = t[66] ^ x[35];
  assign t[54] = t[67] ^ x[38];
  assign t[55] = t[68] ^ x[41];
  assign t[56] = t[69] ^ x[44];
  assign t[57] = (t[70] & ~t[71]);
  assign t[58] = (t[72] & ~t[73]);
  assign t[59] = (t[74] & ~t[75]);
  assign t[5] = t[7];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = t[96] ^ x[5];
  assign t[71] = t[97] ^ x[4];
  assign t[72] = t[98] ^ x[11];
  assign t[73] = t[99] ^ x[10];
  assign t[74] = t[100] ^ x[14];
  assign t[75] = t[101] ^ x[13];
  assign t[76] = t[102] ^ x[17];
  assign t[77] = t[103] ^ x[16];
  assign t[78] = t[104] ^ x[20];
  assign t[79] = t[105] ^ x[19];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[23];
  assign t[81] = t[107] ^ x[22];
  assign t[82] = t[108] ^ x[26];
  assign t[83] = t[109] ^ x[25];
  assign t[84] = t[110] ^ x[29];
  assign t[85] = t[111] ^ x[28];
  assign t[86] = t[112] ^ x[32];
  assign t[87] = t[113] ^ x[31];
  assign t[88] = t[114] ^ x[35];
  assign t[89] = t[115] ^ x[34];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[38];
  assign t[91] = t[117] ^ x[37];
  assign t[92] = t[118] ^ x[41];
  assign t[93] = t[119] ^ x[40];
  assign t[94] = t[120] ^ x[44];
  assign t[95] = t[121] ^ x[43];
  assign t[96] = (x[3]);
  assign t[97] = (x[3]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [44:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = t[126] ^ x[43];
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~x[2] & t[36];
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[125] = (x[42]);
  assign t[126] = (x[42]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[37] | t[23]);
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = ~(t[38] | t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39] | t[29]);
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[41]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[42]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[44]);
  assign t[28] = ~(t[45]);
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[46]);
  assign t[31] = ~(t[40] | t[41]);
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[42] | t[43]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[44] | t[45]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = (t[60]);
  assign t[48] = (t[61]);
  assign t[49] = t[62] ^ x[8];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[11];
  assign t[51] = t[64] ^ x[14];
  assign t[52] = t[65] ^ x[17];
  assign t[53] = t[66] ^ x[20];
  assign t[54] = t[67] ^ x[23];
  assign t[55] = t[68] ^ x[26];
  assign t[56] = t[69] ^ x[29];
  assign t[57] = t[70] ^ x[32];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[38];
  assign t[5] = t[8];
  assign t[60] = t[73] ^ x[41];
  assign t[61] = t[74] ^ x[44];
  assign t[62] = (t[75] & ~t[76]);
  assign t[63] = (t[77] & ~t[78]);
  assign t[64] = (t[79] & ~t[80]);
  assign t[65] = (t[81] & ~t[82]);
  assign t[66] = (t[83] & ~t[84]);
  assign t[67] = (t[85] & ~t[86]);
  assign t[68] = (t[87] & ~t[88]);
  assign t[69] = (t[89] & ~t[90]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[91] & ~t[92]);
  assign t[71] = (t[93] & ~t[94]);
  assign t[72] = (t[95] & ~t[96]);
  assign t[73] = (t[97] & ~t[98]);
  assign t[74] = (t[99] & ~t[100]);
  assign t[75] = t[101] ^ x[8];
  assign t[76] = t[102] ^ x[7];
  assign t[77] = t[103] ^ x[11];
  assign t[78] = t[104] ^ x[10];
  assign t[79] = t[105] ^ x[14];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[13];
  assign t[81] = t[107] ^ x[17];
  assign t[82] = t[108] ^ x[16];
  assign t[83] = t[109] ^ x[20];
  assign t[84] = t[110] ^ x[19];
  assign t[85] = t[111] ^ x[23];
  assign t[86] = t[112] ^ x[22];
  assign t[87] = t[113] ^ x[26];
  assign t[88] = t[114] ^ x[25];
  assign t[89] = t[115] ^ x[29];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[28];
  assign t[91] = t[117] ^ x[32];
  assign t[92] = t[118] ^ x[31];
  assign t[93] = t[119] ^ x[35];
  assign t[94] = t[120] ^ x[34];
  assign t[95] = t[121] ^ x[38];
  assign t[96] = t[122] ^ x[37];
  assign t[97] = t[123] ^ x[41];
  assign t[98] = t[124] ^ x[40];
  assign t[99] = t[125] ^ x[44];
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[11];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[17];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[23];
  assign t[46] = t[56] ^ x[26];
  assign t[47] = t[57] ^ x[29];
  assign t[48] = t[58] ^ x[32];
  assign t[49] = t[59] ^ x[35];
  assign t[4] = ~(t[7]);
  assign t[50] = (t[60] & ~t[61]);
  assign t[51] = (t[62] & ~t[63]);
  assign t[52] = (t[64] & ~t[65]);
  assign t[53] = (t[66] & ~t[67]);
  assign t[54] = (t[68] & ~t[69]);
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[11];
  assign t[63] = t[83] ^ x[10];
  assign t[64] = t[84] ^ x[14];
  assign t[65] = t[85] ^ x[13];
  assign t[66] = t[86] ^ x[17];
  assign t[67] = t[87] ^ x[16];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[23];
  assign t[71] = t[91] ^ x[22];
  assign t[72] = t[92] ^ x[26];
  assign t[73] = t[93] ^ x[25];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[28];
  assign t[76] = t[96] ^ x[32];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[35];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = ~(t[11]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[11] = ~x[2] & t[30];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[31] & t[21]);
  assign t[16] = ~(t[32] & t[22]);
  assign t[17] = ~(t[33] & t[23]);
  assign t[18] = ~(t[34] & t[24]);
  assign t[19] = ~(t[35] & t[25]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[36] & t[26]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[37] & t[27]);
  assign t[23] = ~(t[38]);
  assign t[24] = ~(t[38] & t[28]);
  assign t[25] = ~(t[39]);
  assign t[26] = ~(t[39] & t[29]);
  assign t[27] = ~(t[31]);
  assign t[28] = ~(t[33]);
  assign t[29] = ~(t[35]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = (t[40]);
  assign t[31] = (t[41]);
  assign t[32] = (t[42]);
  assign t[33] = (t[43]);
  assign t[34] = (t[44]);
  assign t[35] = (t[45]);
  assign t[36] = (t[46]);
  assign t[37] = (t[47]);
  assign t[38] = (t[48]);
  assign t[39] = (t[49]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ x[8];
  assign t[41] = t[51] ^ x[11];
  assign t[42] = t[52] ^ x[14];
  assign t[43] = t[53] ^ x[17];
  assign t[44] = t[54] ^ x[20];
  assign t[45] = t[55] ^ x[23];
  assign t[46] = t[56] ^ x[26];
  assign t[47] = t[57] ^ x[29];
  assign t[48] = t[58] ^ x[32];
  assign t[49] = t[59] ^ x[35];
  assign t[4] = ~(t[7]);
  assign t[50] = (t[60] & ~t[61]);
  assign t[51] = (t[62] & ~t[63]);
  assign t[52] = (t[64] & ~t[65]);
  assign t[53] = (t[66] & ~t[67]);
  assign t[54] = (t[68] & ~t[69]);
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[11];
  assign t[63] = t[83] ^ x[10];
  assign t[64] = t[84] ^ x[14];
  assign t[65] = t[85] ^ x[13];
  assign t[66] = t[86] ^ x[17];
  assign t[67] = t[87] ^ x[16];
  assign t[68] = t[88] ^ x[20];
  assign t[69] = t[89] ^ x[19];
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = t[90] ^ x[23];
  assign t[71] = t[91] ^ x[22];
  assign t[72] = t[92] ^ x[26];
  assign t[73] = t[93] ^ x[25];
  assign t[74] = t[94] ^ x[29];
  assign t[75] = t[95] ^ x[28];
  assign t[76] = t[96] ^ x[32];
  assign t[77] = t[97] ^ x[31];
  assign t[78] = t[98] ^ x[35];
  assign t[79] = t[99] ^ x[34];
  assign t[7] = ~(t[11]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind146(x, y);
 input [44:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = ~(t[21] & t[35]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[36]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[39] & t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[11];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[17];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[23];
  assign t[53] = t[66] ^ x[26];
  assign t[54] = t[67] ^ x[29];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = t[70] ^ x[38];
  assign t[58] = t[71] ^ x[41];
  assign t[59] = t[72] ^ x[44];
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]);
  assign t[61] = (t[75] & ~t[76]);
  assign t[62] = (t[77] & ~t[78]);
  assign t[63] = (t[79] & ~t[80]);
  assign t[64] = (t[81] & ~t[82]);
  assign t[65] = (t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[86]);
  assign t[67] = (t[87] & ~t[88]);
  assign t[68] = (t[89] & ~t[90]);
  assign t[69] = (t[91] & ~t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[93] & ~t[94]);
  assign t[71] = (t[95] & ~t[96]);
  assign t[72] = (t[97] & ~t[98]);
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[4];
  assign t[75] = t[101] ^ x[11];
  assign t[76] = t[102] ^ x[10];
  assign t[77] = t[103] ^ x[14];
  assign t[78] = t[104] ^ x[13];
  assign t[79] = t[105] ^ x[17];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[16];
  assign t[81] = t[107] ^ x[20];
  assign t[82] = t[108] ^ x[19];
  assign t[83] = t[109] ^ x[23];
  assign t[84] = t[110] ^ x[22];
  assign t[85] = t[111] ^ x[26];
  assign t[86] = t[112] ^ x[25];
  assign t[87] = t[113] ^ x[29];
  assign t[88] = t[114] ^ x[28];
  assign t[89] = t[115] ^ x[32];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[31];
  assign t[91] = t[117] ^ x[35];
  assign t[92] = t[118] ^ x[34];
  assign t[93] = t[119] ^ x[38];
  assign t[94] = t[120] ^ x[37];
  assign t[95] = t[121] ^ x[41];
  assign t[96] = t[122] ^ x[40];
  assign t[97] = t[123] ^ x[44];
  assign t[98] = t[124] ^ x[43];
  assign t[99] = (x[3]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [44:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[13] & t[14]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = ~(t[15] & t[16]);
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[123] = (x[42]);
  assign t[124] = (x[42]);
  assign t[12] = ~(t[17] & t[18]);
  assign t[13] = ~(t[19] & t[20]);
  assign t[14] = ~(t[21] & t[35]);
  assign t[15] = ~(t[22] & t[23]);
  assign t[16] = ~(t[24] & t[36]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[27] & t[37]);
  assign t[19] = ~(t[38]);
  assign t[1] = ~t[3];
  assign t[20] = ~(t[39]);
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[40]);
  assign t[23] = ~(t[41]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43]);
  assign t[27] = ~(t[32] & t[33]);
  assign t[28] = ~(t[39] & t[38]);
  assign t[29] = ~(t[44]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[41] & t[40]);
  assign t[31] = ~(t[45]);
  assign t[32] = ~(t[43] & t[42]);
  assign t[33] = ~(t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = (t[59]);
  assign t[47] = t[60] ^ x[5];
  assign t[48] = t[61] ^ x[11];
  assign t[49] = t[62] ^ x[14];
  assign t[4] = ~x[2] & t[34];
  assign t[50] = t[63] ^ x[17];
  assign t[51] = t[64] ^ x[20];
  assign t[52] = t[65] ^ x[23];
  assign t[53] = t[66] ^ x[26];
  assign t[54] = t[67] ^ x[29];
  assign t[55] = t[68] ^ x[32];
  assign t[56] = t[69] ^ x[35];
  assign t[57] = t[70] ^ x[38];
  assign t[58] = t[71] ^ x[41];
  assign t[59] = t[72] ^ x[44];
  assign t[5] = t[7];
  assign t[60] = (t[73] & ~t[74]);
  assign t[61] = (t[75] & ~t[76]);
  assign t[62] = (t[77] & ~t[78]);
  assign t[63] = (t[79] & ~t[80]);
  assign t[64] = (t[81] & ~t[82]);
  assign t[65] = (t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[86]);
  assign t[67] = (t[87] & ~t[88]);
  assign t[68] = (t[89] & ~t[90]);
  assign t[69] = (t[91] & ~t[92]);
  assign t[6] = ~(t[8] ^ t[9]);
  assign t[70] = (t[93] & ~t[94]);
  assign t[71] = (t[95] & ~t[96]);
  assign t[72] = (t[97] & ~t[98]);
  assign t[73] = t[99] ^ x[5];
  assign t[74] = t[100] ^ x[4];
  assign t[75] = t[101] ^ x[11];
  assign t[76] = t[102] ^ x[10];
  assign t[77] = t[103] ^ x[14];
  assign t[78] = t[104] ^ x[13];
  assign t[79] = t[105] ^ x[17];
  assign t[7] = x[2] ? x[6] : t[10];
  assign t[80] = t[106] ^ x[16];
  assign t[81] = t[107] ^ x[20];
  assign t[82] = t[108] ^ x[19];
  assign t[83] = t[109] ^ x[23];
  assign t[84] = t[110] ^ x[22];
  assign t[85] = t[111] ^ x[26];
  assign t[86] = t[112] ^ x[25];
  assign t[87] = t[113] ^ x[29];
  assign t[88] = t[114] ^ x[28];
  assign t[89] = t[115] ^ x[32];
  assign t[8] = x[2] ? x[7] : t[11];
  assign t[90] = t[116] ^ x[31];
  assign t[91] = t[117] ^ x[35];
  assign t[92] = t[118] ^ x[34];
  assign t[93] = t[119] ^ x[38];
  assign t[94] = t[120] ^ x[37];
  assign t[95] = t[121] ^ x[41];
  assign t[96] = t[122] ^ x[40];
  assign t[97] = t[123] ^ x[44];
  assign t[98] = t[124] ^ x[43];
  assign t[99] = (x[3]);
  assign t[9] = x[2] ? x[8] : t[12];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [44:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[9]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[15]);
  assign t[105] = (x[15]);
  assign t[106] = (x[18]);
  assign t[107] = (x[18]);
  assign t[108] = (x[21]);
  assign t[109] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[24]);
  assign t[111] = (x[24]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[30]);
  assign t[115] = (x[30]);
  assign t[116] = (x[33]);
  assign t[117] = (x[33]);
  assign t[118] = (x[36]);
  assign t[119] = (x[36]);
  assign t[11] = ~x[2] & t[33];
  assign t[120] = (x[39]);
  assign t[121] = (x[39]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[17];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[20];
  assign t[51] = t[64] ^ x[23];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[32];
  assign t[55] = t[68] ^ x[35];
  assign t[56] = t[69] ^ x[38];
  assign t[57] = t[70] ^ x[41];
  assign t[58] = t[71] ^ x[44];
  assign t[59] = (t[72] & ~t[73]);
  assign t[5] = t[8];
  assign t[60] = (t[74] & ~t[75]);
  assign t[61] = (t[76] & ~t[77]);
  assign t[62] = (t[78] & ~t[79]);
  assign t[63] = (t[80] & ~t[81]);
  assign t[64] = (t[82] & ~t[83]);
  assign t[65] = (t[84] & ~t[85]);
  assign t[66] = (t[86] & ~t[87]);
  assign t[67] = (t[88] & ~t[89]);
  assign t[68] = (t[90] & ~t[91]);
  assign t[69] = (t[92] & ~t[93]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[94] & ~t[95]);
  assign t[71] = (t[96] & ~t[97]);
  assign t[72] = t[98] ^ x[8];
  assign t[73] = t[99] ^ x[7];
  assign t[74] = t[100] ^ x[11];
  assign t[75] = t[101] ^ x[10];
  assign t[76] = t[102] ^ x[14];
  assign t[77] = t[103] ^ x[13];
  assign t[78] = t[104] ^ x[17];
  assign t[79] = t[105] ^ x[16];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[20];
  assign t[81] = t[107] ^ x[19];
  assign t[82] = t[108] ^ x[23];
  assign t[83] = t[109] ^ x[22];
  assign t[84] = t[110] ^ x[26];
  assign t[85] = t[111] ^ x[25];
  assign t[86] = t[112] ^ x[29];
  assign t[87] = t[113] ^ x[28];
  assign t[88] = t[114] ^ x[32];
  assign t[89] = t[115] ^ x[31];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[35];
  assign t[91] = t[117] ^ x[34];
  assign t[92] = t[118] ^ x[38];
  assign t[93] = t[119] ^ x[37];
  assign t[94] = t[120] ^ x[41];
  assign t[95] = t[121] ^ x[40];
  assign t[96] = t[122] ^ x[44];
  assign t[97] = t[123] ^ x[43];
  assign t[98] = (x[6]);
  assign t[99] = (x[6]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [44:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[100] = (x[9]);
  assign t[101] = (x[9]);
  assign t[102] = (x[12]);
  assign t[103] = (x[12]);
  assign t[104] = (x[15]);
  assign t[105] = (x[15]);
  assign t[106] = (x[18]);
  assign t[107] = (x[18]);
  assign t[108] = (x[21]);
  assign t[109] = (x[21]);
  assign t[10] = x[2] ? x[5] : t[14];
  assign t[110] = (x[24]);
  assign t[111] = (x[24]);
  assign t[112] = (x[27]);
  assign t[113] = (x[27]);
  assign t[114] = (x[30]);
  assign t[115] = (x[30]);
  assign t[116] = (x[33]);
  assign t[117] = (x[33]);
  assign t[118] = (x[36]);
  assign t[119] = (x[36]);
  assign t[11] = ~x[2] & t[33];
  assign t[120] = (x[39]);
  assign t[121] = (x[39]);
  assign t[122] = (x[42]);
  assign t[123] = (x[42]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = t[23] | t[34];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = t[26] | t[35];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~t[3];
  assign t[20] = t[29] | t[36];
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[38]);
  assign t[23] = ~(t[30] | t[21]);
  assign t[24] = ~(t[39]);
  assign t[25] = ~(t[40]);
  assign t[26] = ~(t[31] | t[24]);
  assign t[27] = ~(t[41]);
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[32] | t[27]);
  assign t[2] = t[4] ? x[1] : x[0];
  assign t[30] = ~(t[43]);
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = (t[50]);
  assign t[38] = (t[51]);
  assign t[39] = (t[52]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = (t[53]);
  assign t[41] = (t[54]);
  assign t[42] = (t[55]);
  assign t[43] = (t[56]);
  assign t[44] = (t[57]);
  assign t[45] = (t[58]);
  assign t[46] = t[59] ^ x[8];
  assign t[47] = t[60] ^ x[11];
  assign t[48] = t[61] ^ x[14];
  assign t[49] = t[62] ^ x[17];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ x[20];
  assign t[51] = t[64] ^ x[23];
  assign t[52] = t[65] ^ x[26];
  assign t[53] = t[66] ^ x[29];
  assign t[54] = t[67] ^ x[32];
  assign t[55] = t[68] ^ x[35];
  assign t[56] = t[69] ^ x[38];
  assign t[57] = t[70] ^ x[41];
  assign t[58] = t[71] ^ x[44];
  assign t[59] = (t[72] & ~t[73]);
  assign t[5] = t[8];
  assign t[60] = (t[74] & ~t[75]);
  assign t[61] = (t[76] & ~t[77]);
  assign t[62] = (t[78] & ~t[79]);
  assign t[63] = (t[80] & ~t[81]);
  assign t[64] = (t[82] & ~t[83]);
  assign t[65] = (t[84] & ~t[85]);
  assign t[66] = (t[86] & ~t[87]);
  assign t[67] = (t[88] & ~t[89]);
  assign t[68] = (t[90] & ~t[91]);
  assign t[69] = (t[92] & ~t[93]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[94] & ~t[95]);
  assign t[71] = (t[96] & ~t[97]);
  assign t[72] = t[98] ^ x[8];
  assign t[73] = t[99] ^ x[7];
  assign t[74] = t[100] ^ x[11];
  assign t[75] = t[101] ^ x[10];
  assign t[76] = t[102] ^ x[14];
  assign t[77] = t[103] ^ x[13];
  assign t[78] = t[104] ^ x[17];
  assign t[79] = t[105] ^ x[16];
  assign t[7] = ~(t[11]);
  assign t[80] = t[106] ^ x[20];
  assign t[81] = t[107] ^ x[19];
  assign t[82] = t[108] ^ x[23];
  assign t[83] = t[109] ^ x[22];
  assign t[84] = t[110] ^ x[26];
  assign t[85] = t[111] ^ x[25];
  assign t[86] = t[112] ^ x[29];
  assign t[87] = t[113] ^ x[28];
  assign t[88] = t[114] ^ x[32];
  assign t[89] = t[115] ^ x[31];
  assign t[8] = x[2] ? x[3] : t[12];
  assign t[90] = t[116] ^ x[35];
  assign t[91] = t[117] ^ x[34];
  assign t[92] = t[118] ^ x[38];
  assign t[93] = t[119] ^ x[37];
  assign t[94] = t[120] ^ x[41];
  assign t[95] = t[121] ^ x[40];
  assign t[96] = t[122] ^ x[44];
  assign t[97] = t[123] ^ x[43];
  assign t[98] = (x[6]);
  assign t[99] = (x[6]);
  assign t[9] = x[2] ? x[4] : t[13];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [414:0] x;
 output [149:0] y;

  R2ind0 R2ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[2], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[15], x[14], x[13], x[3]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[15], x[14], x[13], x[3]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[12], x[11], x[10], x[3]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[12], x[11], x[10], x[3]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[9], x[8], x[7], x[15], x[14], x[13], x[3]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[9], x[8], x[7], x[15], x[14], x[13], x[3]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[21], x[20], x[19], x[3]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[21], x[20], x[19], x[3]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[24], x[23], x[22], x[3]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[24], x[23], x[22], x[3]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[6], x[5], x[4], x[3]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[6], x[5], x[4], x[3]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[21], x[20], x[19], x[18], x[17], x[16], x[3]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[21], x[20], x[19], x[18], x[17], x[16], x[3]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[27], x[26], x[25], x[3]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[27], x[26], x[25], x[3]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[27], x[26], x[25], x[30], x[29], x[28], x[3]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[27], x[26], x[25], x[30], x[29], x[28], x[3]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[27], x[26], x[25], x[33], x[3], x[32], x[31]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[27], x[26], x[25], x[33], x[3], x[32], x[31]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[42], x[41], x[40], x[27], x[26], x[25], x[45], x[44], x[43], x[39], x[38], x[37], x[48], x[3], x[47], x[46]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[42], x[41], x[40], x[27], x[26], x[25], x[45], x[44], x[43], x[39], x[38], x[37], x[48], x[3], x[47], x[46]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[39], x[38], x[37], x[45], x[44], x[43], x[42], x[41], x[40], x[36], x[35], x[34], x[27], x[26], x[25], x[51], x[3], x[50], x[49]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[39], x[38], x[37], x[45], x[44], x[43], x[42], x[41], x[40], x[36], x[35], x[34], x[27], x[26], x[25], x[51], x[3], x[50], x[49]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[39], x[38], x[37], x[45], x[44], x[43], x[42], x[41], x[40], x[27], x[26], x[25], x[36], x[35], x[34], x[54], x[3], x[53], x[52]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[39], x[38], x[37], x[45], x[44], x[43], x[42], x[41], x[40], x[27], x[26], x[25], x[36], x[35], x[34], x[54], x[3], x[53], x[52]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[27], x[26], x[25], x[60], x[59], x[58], x[57], x[3], x[56], x[55]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[27], x[26], x[25], x[60], x[59], x[58], x[57], x[3], x[56], x[55]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[66], x[65], x[64], x[27], x[26], x[25], x[69], x[68], x[67], x[63], x[62], x[61], x[72], x[3], x[71], x[70]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[66], x[65], x[64], x[27], x[26], x[25], x[69], x[68], x[67], x[63], x[62], x[61], x[72], x[3], x[71], x[70]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[27], x[26], x[25], x[60], x[59], x[58], x[75], x[3], x[74], x[73]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[27], x[26], x[25], x[60], x[59], x[58], x[75], x[3], x[74], x[73]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[27], x[26], x[25], x[60], x[59], x[58], x[78], x[3], x[77], x[76]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[63], x[62], x[61], x[69], x[68], x[67], x[66], x[65], x[64], x[27], x[26], x[25], x[60], x[59], x[58], x[78], x[3], x[77], x[76]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[27], x[26], x[25], x[84], x[83], x[82], x[81], x[3], x[80], x[79]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[27], x[26], x[25], x[84], x[83], x[82], x[81], x[3], x[80], x[79]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[90], x[89], x[88], x[27], x[26], x[25], x[93], x[92], x[91], x[87], x[86], x[85], x[96], x[3], x[95], x[94]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[90], x[89], x[88], x[27], x[26], x[25], x[93], x[92], x[91], x[87], x[86], x[85], x[96], x[3], x[95], x[94]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[87], x[86], x[85], x[93], x[92], x[91], x[90], x[89], x[88], x[27], x[26], x[25], x[84], x[83], x[82], x[99], x[3], x[98], x[97]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[87], x[86], x[85], x[93], x[92], x[91], x[90], x[89], x[88], x[27], x[26], x[25], x[84], x[83], x[82], x[99], x[3], x[98], x[97]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[87], x[86], x[85], x[93], x[92], x[91], x[90], x[89], x[88], x[27], x[26], x[25], x[84], x[83], x[82], x[102], x[3], x[101], x[100]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[87], x[86], x[85], x[93], x[92], x[91], x[90], x[89], x[88], x[27], x[26], x[25], x[84], x[83], x[82], x[102], x[3], x[101], x[100]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[27], x[26], x[25], x[108], x[107], x[106], x[105], x[3], x[104], x[103]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[27], x[26], x[25], x[108], x[107], x[106], x[105], x[3], x[104], x[103]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[114], x[113], x[112], x[27], x[26], x[25], x[117], x[116], x[115], x[111], x[110], x[109], x[120], x[3], x[119], x[118]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[114], x[113], x[112], x[27], x[26], x[25], x[117], x[116], x[115], x[111], x[110], x[109], x[120], x[3], x[119], x[118]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[111], x[110], x[109], x[117], x[116], x[115], x[114], x[113], x[112], x[27], x[26], x[25], x[108], x[107], x[106], x[123], x[3], x[122], x[121]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[111], x[110], x[109], x[117], x[116], x[115], x[114], x[113], x[112], x[27], x[26], x[25], x[108], x[107], x[106], x[123], x[3], x[122], x[121]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[111], x[110], x[109], x[117], x[116], x[115], x[114], x[113], x[112], x[27], x[26], x[25], x[108], x[107], x[106], x[126], x[3], x[125], x[124]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[111], x[110], x[109], x[117], x[116], x[115], x[114], x[113], x[112], x[27], x[26], x[25], x[108], x[107], x[106], x[126], x[3], x[125], x[124]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[27], x[26], x[25], x[132], x[131], x[130], x[129], x[3], x[128], x[127]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[27], x[26], x[25], x[132], x[131], x[130], x[129], x[3], x[128], x[127]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[138], x[137], x[136], x[27], x[26], x[25], x[141], x[140], x[139], x[135], x[134], x[133], x[144], x[3], x[143], x[142]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[138], x[137], x[136], x[27], x[26], x[25], x[141], x[140], x[139], x[135], x[134], x[133], x[144], x[3], x[143], x[142]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[135], x[134], x[133], x[141], x[140], x[139], x[138], x[137], x[136], x[27], x[26], x[25], x[132], x[131], x[130], x[147], x[3], x[146], x[145]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[135], x[134], x[133], x[141], x[140], x[139], x[138], x[137], x[136], x[27], x[26], x[25], x[132], x[131], x[130], x[147], x[3], x[146], x[145]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[135], x[134], x[133], x[141], x[140], x[139], x[138], x[137], x[136], x[27], x[26], x[25], x[132], x[131], x[130], x[150], x[3], x[149], x[148]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[135], x[134], x[133], x[141], x[140], x[139], x[138], x[137], x[136], x[27], x[26], x[25], x[132], x[131], x[130], x[150], x[3], x[149], x[148]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[27], x[26], x[25], x[156], x[155], x[154], x[153], x[3], x[152], x[151]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[27], x[26], x[25], x[156], x[155], x[154], x[153], x[3], x[152], x[151]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[162], x[161], x[160], x[27], x[26], x[25], x[165], x[164], x[163], x[159], x[158], x[157], x[168], x[3], x[167], x[166]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[162], x[161], x[160], x[27], x[26], x[25], x[165], x[164], x[163], x[159], x[158], x[157], x[168], x[3], x[167], x[166]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[159], x[158], x[157], x[165], x[164], x[163], x[162], x[161], x[160], x[156], x[155], x[154], x[27], x[26], x[25], x[171], x[3], x[170], x[169]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[159], x[158], x[157], x[165], x[164], x[163], x[162], x[161], x[160], x[156], x[155], x[154], x[27], x[26], x[25], x[171], x[3], x[170], x[169]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[159], x[158], x[157], x[165], x[164], x[163], x[162], x[161], x[160], x[156], x[155], x[154], x[27], x[26], x[25], x[174], x[3], x[173], x[172]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[159], x[158], x[157], x[165], x[164], x[163], x[162], x[161], x[160], x[156], x[155], x[154], x[27], x[26], x[25], x[174], x[3], x[173], x[172]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[27], x[26], x[25], x[177], x[3], x[176], x[175]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[27], x[26], x[25], x[177], x[3], x[176], x[175]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[186], x[185], x[184], x[189], x[188], x[187], x[183], x[182], x[181], x[27], x[26], x[25], x[192], x[3], x[191], x[190]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[186], x[185], x[184], x[189], x[188], x[187], x[183], x[182], x[181], x[27], x[26], x[25], x[192], x[3], x[191], x[190]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[27], x[26], x[25], x[195], x[3], x[194], x[193]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[27], x[26], x[25], x[195], x[3], x[194], x[193]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[27], x[26], x[25], x[198], x[3], x[197], x[196]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[183], x[182], x[181], x[189], x[188], x[187], x[186], x[185], x[184], x[180], x[179], x[178], x[27], x[26], x[25], x[198], x[3], x[197], x[196]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[27], x[26], x[25], x[204], x[203], x[202], x[201], x[3], x[200], x[199]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[27], x[26], x[25], x[204], x[203], x[202], x[201], x[3], x[200], x[199]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[210], x[209], x[208], x[27], x[26], x[25], x[213], x[212], x[211], x[207], x[206], x[205], x[216], x[3], x[215], x[214]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[210], x[209], x[208], x[27], x[26], x[25], x[213], x[212], x[211], x[207], x[206], x[205], x[216], x[3], x[215], x[214]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[207], x[206], x[205], x[213], x[212], x[211], x[210], x[209], x[208], x[27], x[26], x[25], x[204], x[203], x[202], x[219], x[3], x[218], x[217]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[207], x[206], x[205], x[213], x[212], x[211], x[210], x[209], x[208], x[27], x[26], x[25], x[204], x[203], x[202], x[219], x[3], x[218], x[217]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[207], x[206], x[205], x[213], x[212], x[211], x[210], x[209], x[208], x[27], x[26], x[25], x[204], x[203], x[202], x[222], x[3], x[221], x[220]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[207], x[206], x[205], x[213], x[212], x[211], x[210], x[209], x[208], x[27], x[26], x[25], x[204], x[203], x[202], x[222], x[3], x[221], x[220]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[237], x[236], x[235], x[45], x[44], x[43], x[234], x[233], x[232], x[231], x[230], x[229], x[42], x[41], x[40], x[39], x[38], x[37], x[228], x[227], x[226], x[36], x[35], x[34], x[27], x[26], x[25], x[225], x[33], x[3], x[224], x[223]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[237], x[236], x[235], x[45], x[44], x[43], x[234], x[233], x[232], x[231], x[230], x[229], x[42], x[41], x[40], x[39], x[38], x[37], x[228], x[227], x[226], x[36], x[35], x[34], x[27], x[26], x[25], x[225], x[33], x[3], x[224], x[223]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[234], x[233], x[232], x[42], x[41], x[40], x[237], x[236], x[235], x[231], x[230], x[229], x[45], x[44], x[43], x[39], x[38], x[37], x[240], x[48], x[27], x[26], x[25], x[3], x[239], x[238]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[234], x[233], x[232], x[42], x[41], x[40], x[237], x[236], x[235], x[231], x[230], x[229], x[45], x[44], x[43], x[39], x[38], x[37], x[240], x[48], x[27], x[26], x[25], x[3], x[239], x[238]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[231], x[230], x[229], x[39], x[38], x[37], x[237], x[236], x[235], x[234], x[233], x[232], x[45], x[44], x[43], x[42], x[41], x[40], x[228], x[227], x[226], x[36], x[35], x[34], x[27], x[26], x[25], x[243], x[51], x[3], x[242], x[241]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[231], x[230], x[229], x[39], x[38], x[37], x[237], x[236], x[235], x[234], x[233], x[232], x[45], x[44], x[43], x[42], x[41], x[40], x[228], x[227], x[226], x[36], x[35], x[34], x[27], x[26], x[25], x[243], x[51], x[3], x[242], x[241]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[231], x[230], x[229], x[39], x[38], x[37], x[237], x[236], x[235], x[234], x[233], x[232], x[45], x[44], x[43], x[42], x[41], x[40], x[228], x[227], x[226], x[36], x[35], x[34], x[27], x[26], x[25], x[246], x[54], x[3], x[245], x[244]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[231], x[230], x[229], x[39], x[38], x[37], x[237], x[236], x[235], x[234], x[233], x[232], x[45], x[44], x[43], x[42], x[41], x[40], x[228], x[227], x[226], x[36], x[35], x[34], x[27], x[26], x[25], x[246], x[54], x[3], x[245], x[244]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[261], x[260], x[259], x[69], x[68], x[67], x[258], x[257], x[256], x[255], x[254], x[253], x[66], x[65], x[64], x[63], x[62], x[61], x[252], x[251], x[250], x[60], x[59], x[58], x[249], x[57], x[27], x[26], x[25], x[3], x[248], x[247]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[261], x[260], x[259], x[69], x[68], x[67], x[258], x[257], x[256], x[255], x[254], x[253], x[66], x[65], x[64], x[63], x[62], x[61], x[252], x[251], x[250], x[60], x[59], x[58], x[249], x[57], x[27], x[26], x[25], x[3], x[248], x[247]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[258], x[257], x[256], x[66], x[65], x[64], x[261], x[260], x[259], x[255], x[254], x[253], x[69], x[68], x[67], x[63], x[62], x[61], x[27], x[26], x[25], x[264], x[72], x[3], x[263], x[262]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[258], x[257], x[256], x[66], x[65], x[64], x[261], x[260], x[259], x[255], x[254], x[253], x[69], x[68], x[67], x[63], x[62], x[61], x[27], x[26], x[25], x[264], x[72], x[3], x[263], x[262]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[255], x[254], x[253], x[63], x[62], x[61], x[261], x[260], x[259], x[258], x[257], x[256], x[69], x[68], x[67], x[66], x[65], x[64], x[252], x[251], x[250], x[60], x[59], x[58], x[27], x[26], x[25], x[267], x[75], x[3], x[266], x[265]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[255], x[254], x[253], x[63], x[62], x[61], x[261], x[260], x[259], x[258], x[257], x[256], x[69], x[68], x[67], x[66], x[65], x[64], x[252], x[251], x[250], x[60], x[59], x[58], x[27], x[26], x[25], x[267], x[75], x[3], x[266], x[265]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[255], x[254], x[253], x[63], x[62], x[61], x[261], x[260], x[259], x[258], x[257], x[256], x[69], x[68], x[67], x[66], x[65], x[64], x[252], x[251], x[250], x[60], x[59], x[58], x[270], x[78], x[27], x[26], x[25], x[3], x[269], x[268]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[255], x[254], x[253], x[63], x[62], x[61], x[261], x[260], x[259], x[258], x[257], x[256], x[69], x[68], x[67], x[66], x[65], x[64], x[252], x[251], x[250], x[60], x[59], x[58], x[270], x[78], x[27], x[26], x[25], x[3], x[269], x[268]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[285], x[284], x[283], x[93], x[92], x[91], x[282], x[281], x[280], x[279], x[278], x[277], x[90], x[89], x[88], x[87], x[86], x[85], x[276], x[275], x[274], x[27], x[26], x[25], x[84], x[83], x[82], x[273], x[81], x[9], x[8], x[7], x[3], x[272], x[271]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[285], x[284], x[283], x[93], x[92], x[91], x[282], x[281], x[280], x[279], x[278], x[277], x[90], x[89], x[88], x[87], x[86], x[85], x[276], x[275], x[274], x[27], x[26], x[25], x[84], x[83], x[82], x[273], x[81], x[9], x[8], x[7], x[3], x[272], x[271]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[282], x[281], x[280], x[90], x[89], x[88], x[285], x[284], x[283], x[279], x[278], x[277], x[27], x[26], x[25], x[93], x[92], x[91], x[87], x[86], x[85], x[288], x[96], x[15], x[14], x[13], x[3], x[287], x[286]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[282], x[281], x[280], x[90], x[89], x[88], x[285], x[284], x[283], x[279], x[278], x[277], x[27], x[26], x[25], x[93], x[92], x[91], x[87], x[86], x[85], x[288], x[96], x[15], x[14], x[13], x[3], x[287], x[286]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[279], x[278], x[277], x[87], x[86], x[85], x[285], x[284], x[283], x[282], x[281], x[280], x[93], x[92], x[91], x[90], x[89], x[88], x[276], x[275], x[274], x[27], x[26], x[25], x[84], x[83], x[82], x[291], x[99], x[12], x[11], x[10], x[3], x[290], x[289]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[279], x[278], x[277], x[87], x[86], x[85], x[285], x[284], x[283], x[282], x[281], x[280], x[93], x[92], x[91], x[90], x[89], x[88], x[276], x[275], x[274], x[27], x[26], x[25], x[84], x[83], x[82], x[291], x[99], x[12], x[11], x[10], x[3], x[290], x[289]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[279], x[278], x[277], x[87], x[86], x[85], x[285], x[284], x[283], x[282], x[281], x[280], x[93], x[92], x[91], x[90], x[89], x[88], x[276], x[275], x[274], x[27], x[26], x[25], x[84], x[83], x[82], x[294], x[102], x[3], x[293], x[292]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[279], x[278], x[277], x[87], x[86], x[85], x[285], x[284], x[283], x[282], x[281], x[280], x[93], x[92], x[91], x[90], x[89], x[88], x[276], x[275], x[274], x[27], x[26], x[25], x[84], x[83], x[82], x[294], x[102], x[3], x[293], x[292]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[309], x[308], x[307], x[117], x[116], x[115], x[306], x[305], x[304], x[303], x[302], x[301], x[114], x[113], x[112], x[111], x[110], x[109], x[300], x[299], x[298], x[27], x[26], x[25], x[108], x[107], x[106], x[297], x[105], x[18], x[17], x[16], x[3], x[296], x[295]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[309], x[308], x[307], x[117], x[116], x[115], x[306], x[305], x[304], x[303], x[302], x[301], x[114], x[113], x[112], x[111], x[110], x[109], x[300], x[299], x[298], x[27], x[26], x[25], x[108], x[107], x[106], x[297], x[105], x[18], x[17], x[16], x[3], x[296], x[295]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[306], x[305], x[304], x[114], x[113], x[112], x[309], x[308], x[307], x[303], x[302], x[301], x[27], x[26], x[25], x[117], x[116], x[115], x[111], x[110], x[109], x[312], x[120], x[21], x[20], x[19], x[3], x[311], x[310]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[306], x[305], x[304], x[114], x[113], x[112], x[309], x[308], x[307], x[303], x[302], x[301], x[27], x[26], x[25], x[117], x[116], x[115], x[111], x[110], x[109], x[312], x[120], x[21], x[20], x[19], x[3], x[311], x[310]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[303], x[302], x[301], x[111], x[110], x[109], x[309], x[308], x[307], x[306], x[305], x[304], x[117], x[116], x[115], x[114], x[113], x[112], x[300], x[299], x[298], x[27], x[26], x[25], x[108], x[107], x[106], x[315], x[123], x[24], x[23], x[22], x[3], x[314], x[313]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[303], x[302], x[301], x[111], x[110], x[109], x[309], x[308], x[307], x[306], x[305], x[304], x[117], x[116], x[115], x[114], x[113], x[112], x[300], x[299], x[298], x[27], x[26], x[25], x[108], x[107], x[106], x[315], x[123], x[24], x[23], x[22], x[3], x[314], x[313]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[303], x[302], x[301], x[111], x[110], x[109], x[309], x[308], x[307], x[306], x[305], x[304], x[117], x[116], x[115], x[114], x[113], x[112], x[300], x[299], x[298], x[27], x[26], x[25], x[108], x[107], x[106], x[318], x[126], x[6], x[5], x[4], x[3], x[317], x[316]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[303], x[302], x[301], x[111], x[110], x[109], x[309], x[308], x[307], x[306], x[305], x[304], x[117], x[116], x[115], x[114], x[113], x[112], x[300], x[299], x[298], x[27], x[26], x[25], x[108], x[107], x[106], x[318], x[126], x[6], x[5], x[4], x[3], x[317], x[316]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[45], x[44], x[43], x[141], x[140], x[139], x[333], x[332], x[331], x[42], x[41], x[40], x[39], x[38], x[37], x[138], x[137], x[136], x[135], x[134], x[133], x[330], x[329], x[328], x[327], x[326], x[325], x[36], x[35], x[34], x[132], x[131], x[130], x[324], x[323], x[322], x[27], x[26], x[25], x[33], x[129], x[321], x[3], x[320], x[319]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[45], x[44], x[43], x[141], x[140], x[139], x[333], x[332], x[331], x[42], x[41], x[40], x[39], x[38], x[37], x[138], x[137], x[136], x[135], x[134], x[133], x[330], x[329], x[328], x[327], x[326], x[325], x[36], x[35], x[34], x[132], x[131], x[130], x[324], x[323], x[322], x[27], x[26], x[25], x[33], x[129], x[321], x[3], x[320], x[319]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[42], x[41], x[40], x[138], x[137], x[136], x[330], x[329], x[328], x[45], x[44], x[43], x[39], x[38], x[37], x[141], x[140], x[139], x[135], x[134], x[133], x[333], x[332], x[331], x[327], x[326], x[325], x[27], x[26], x[25], x[48], x[144], x[336], x[3], x[335], x[334]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[42], x[41], x[40], x[138], x[137], x[136], x[330], x[329], x[328], x[45], x[44], x[43], x[39], x[38], x[37], x[141], x[140], x[139], x[135], x[134], x[133], x[333], x[332], x[331], x[327], x[326], x[325], x[27], x[26], x[25], x[48], x[144], x[336], x[3], x[335], x[334]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[39], x[38], x[37], x[135], x[134], x[133], x[327], x[326], x[325], x[45], x[44], x[43], x[42], x[41], x[40], x[141], x[140], x[139], x[138], x[137], x[136], x[333], x[332], x[331], x[330], x[329], x[328], x[36], x[35], x[34], x[132], x[131], x[130], x[324], x[323], x[322], x[27], x[26], x[25], x[51], x[147], x[339], x[3], x[338], x[337]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[39], x[38], x[37], x[135], x[134], x[133], x[327], x[326], x[325], x[45], x[44], x[43], x[42], x[41], x[40], x[141], x[140], x[139], x[138], x[137], x[136], x[333], x[332], x[331], x[330], x[329], x[328], x[36], x[35], x[34], x[132], x[131], x[130], x[324], x[323], x[322], x[27], x[26], x[25], x[51], x[147], x[339], x[3], x[338], x[337]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[39], x[38], x[37], x[135], x[134], x[133], x[327], x[326], x[325], x[45], x[44], x[43], x[42], x[41], x[40], x[141], x[140], x[139], x[138], x[137], x[136], x[333], x[332], x[331], x[330], x[329], x[328], x[36], x[35], x[34], x[132], x[131], x[130], x[324], x[323], x[322], x[27], x[26], x[25], x[54], x[150], x[342], x[3], x[341], x[340]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[39], x[38], x[37], x[135], x[134], x[133], x[327], x[326], x[325], x[45], x[44], x[43], x[42], x[41], x[40], x[141], x[140], x[139], x[138], x[137], x[136], x[333], x[332], x[331], x[330], x[329], x[328], x[36], x[35], x[34], x[132], x[131], x[130], x[324], x[323], x[322], x[27], x[26], x[25], x[54], x[150], x[342], x[3], x[341], x[340]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[69], x[68], x[67], x[165], x[164], x[163], x[357], x[356], x[355], x[66], x[65], x[64], x[63], x[62], x[61], x[162], x[161], x[160], x[159], x[158], x[157], x[354], x[353], x[352], x[351], x[350], x[349], x[60], x[59], x[58], x[156], x[155], x[154], x[348], x[347], x[346], x[27], x[26], x[25], x[57], x[153], x[345], x[3], x[344], x[343]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[69], x[68], x[67], x[165], x[164], x[163], x[357], x[356], x[355], x[66], x[65], x[64], x[63], x[62], x[61], x[162], x[161], x[160], x[159], x[158], x[157], x[354], x[353], x[352], x[351], x[350], x[349], x[60], x[59], x[58], x[156], x[155], x[154], x[348], x[347], x[346], x[27], x[26], x[25], x[57], x[153], x[345], x[3], x[344], x[343]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[66], x[65], x[64], x[162], x[161], x[160], x[354], x[353], x[352], x[69], x[68], x[67], x[63], x[62], x[61], x[165], x[164], x[163], x[159], x[158], x[157], x[357], x[356], x[355], x[351], x[350], x[349], x[72], x[168], x[360], x[27], x[26], x[25], x[3], x[359], x[358]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[66], x[65], x[64], x[162], x[161], x[160], x[354], x[353], x[352], x[69], x[68], x[67], x[63], x[62], x[61], x[165], x[164], x[163], x[159], x[158], x[157], x[357], x[356], x[355], x[351], x[350], x[349], x[72], x[168], x[360], x[27], x[26], x[25], x[3], x[359], x[358]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[63], x[62], x[61], x[159], x[158], x[157], x[351], x[350], x[349], x[69], x[68], x[67], x[66], x[65], x[64], x[165], x[164], x[163], x[162], x[161], x[160], x[357], x[356], x[355], x[354], x[353], x[352], x[60], x[59], x[58], x[156], x[155], x[154], x[348], x[347], x[346], x[75], x[171], x[363], x[27], x[26], x[25], x[3], x[362], x[361]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[63], x[62], x[61], x[159], x[158], x[157], x[351], x[350], x[349], x[69], x[68], x[67], x[66], x[65], x[64], x[165], x[164], x[163], x[162], x[161], x[160], x[357], x[356], x[355], x[354], x[353], x[352], x[60], x[59], x[58], x[156], x[155], x[154], x[348], x[347], x[346], x[75], x[171], x[363], x[27], x[26], x[25], x[3], x[362], x[361]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[63], x[62], x[61], x[159], x[158], x[157], x[351], x[350], x[349], x[69], x[68], x[67], x[66], x[65], x[64], x[165], x[164], x[163], x[162], x[161], x[160], x[357], x[356], x[355], x[354], x[353], x[352], x[60], x[59], x[58], x[156], x[155], x[154], x[348], x[347], x[346], x[27], x[26], x[25], x[78], x[174], x[366], x[3], x[365], x[364]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[63], x[62], x[61], x[159], x[158], x[157], x[351], x[350], x[349], x[69], x[68], x[67], x[66], x[65], x[64], x[165], x[164], x[163], x[162], x[161], x[160], x[357], x[356], x[355], x[354], x[353], x[352], x[60], x[59], x[58], x[156], x[155], x[154], x[348], x[347], x[346], x[27], x[26], x[25], x[78], x[174], x[366], x[3], x[365], x[364]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[93], x[92], x[91], x[189], x[188], x[187], x[381], x[380], x[379], x[90], x[89], x[88], x[87], x[86], x[85], x[186], x[185], x[184], x[183], x[182], x[181], x[378], x[377], x[376], x[375], x[374], x[373], x[84], x[83], x[82], x[180], x[179], x[178], x[372], x[371], x[370], x[81], x[177], x[369], x[27], x[26], x[25], x[3], x[368], x[367]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[93], x[92], x[91], x[189], x[188], x[187], x[381], x[380], x[379], x[90], x[89], x[88], x[87], x[86], x[85], x[186], x[185], x[184], x[183], x[182], x[181], x[378], x[377], x[376], x[375], x[374], x[373], x[84], x[83], x[82], x[180], x[179], x[178], x[372], x[371], x[370], x[81], x[177], x[369], x[27], x[26], x[25], x[3], x[368], x[367]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[90], x[89], x[88], x[186], x[185], x[184], x[378], x[377], x[376], x[93], x[92], x[91], x[87], x[86], x[85], x[189], x[188], x[187], x[183], x[182], x[181], x[381], x[380], x[379], x[375], x[374], x[373], x[27], x[26], x[25], x[96], x[192], x[384], x[3], x[383], x[382]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[90], x[89], x[88], x[186], x[185], x[184], x[378], x[377], x[376], x[93], x[92], x[91], x[87], x[86], x[85], x[189], x[188], x[187], x[183], x[182], x[181], x[381], x[380], x[379], x[375], x[374], x[373], x[27], x[26], x[25], x[96], x[192], x[384], x[3], x[383], x[382]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[87], x[86], x[85], x[183], x[182], x[181], x[375], x[374], x[373], x[93], x[92], x[91], x[90], x[89], x[88], x[189], x[188], x[187], x[186], x[185], x[184], x[381], x[380], x[379], x[378], x[377], x[376], x[84], x[83], x[82], x[180], x[179], x[178], x[372], x[371], x[370], x[27], x[26], x[25], x[99], x[195], x[387], x[3], x[386], x[385]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[87], x[86], x[85], x[183], x[182], x[181], x[375], x[374], x[373], x[93], x[92], x[91], x[90], x[89], x[88], x[189], x[188], x[187], x[186], x[185], x[184], x[381], x[380], x[379], x[378], x[377], x[376], x[84], x[83], x[82], x[180], x[179], x[178], x[372], x[371], x[370], x[27], x[26], x[25], x[99], x[195], x[387], x[3], x[386], x[385]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[87], x[86], x[85], x[183], x[182], x[181], x[375], x[374], x[373], x[93], x[92], x[91], x[90], x[89], x[88], x[189], x[188], x[187], x[186], x[185], x[184], x[381], x[380], x[379], x[378], x[377], x[376], x[84], x[83], x[82], x[180], x[179], x[178], x[372], x[371], x[370], x[102], x[198], x[390], x[27], x[26], x[25], x[3], x[389], x[388]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[87], x[86], x[85], x[183], x[182], x[181], x[375], x[374], x[373], x[93], x[92], x[91], x[90], x[89], x[88], x[189], x[188], x[187], x[186], x[185], x[184], x[381], x[380], x[379], x[378], x[377], x[376], x[84], x[83], x[82], x[180], x[179], x[178], x[372], x[371], x[370], x[102], x[198], x[390], x[27], x[26], x[25], x[3], x[389], x[388]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[117], x[116], x[115], x[213], x[212], x[211], x[405], x[404], x[403], x[114], x[113], x[112], x[111], x[110], x[109], x[210], x[209], x[208], x[207], x[206], x[205], x[402], x[401], x[400], x[399], x[398], x[397], x[108], x[107], x[106], x[204], x[203], x[202], x[396], x[395], x[394], x[27], x[26], x[25], x[105], x[201], x[393], x[3], x[392], x[391]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[117], x[116], x[115], x[213], x[212], x[211], x[405], x[404], x[403], x[114], x[113], x[112], x[111], x[110], x[109], x[210], x[209], x[208], x[207], x[206], x[205], x[402], x[401], x[400], x[399], x[398], x[397], x[108], x[107], x[106], x[204], x[203], x[202], x[396], x[395], x[394], x[27], x[26], x[25], x[105], x[201], x[393], x[3], x[392], x[391]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[114], x[113], x[112], x[210], x[209], x[208], x[402], x[401], x[400], x[117], x[116], x[115], x[111], x[110], x[109], x[213], x[212], x[211], x[207], x[206], x[205], x[405], x[404], x[403], x[399], x[398], x[397], x[27], x[26], x[25], x[120], x[216], x[408], x[3], x[407], x[406]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[114], x[113], x[112], x[210], x[209], x[208], x[402], x[401], x[400], x[117], x[116], x[115], x[111], x[110], x[109], x[213], x[212], x[211], x[207], x[206], x[205], x[405], x[404], x[403], x[399], x[398], x[397], x[27], x[26], x[25], x[120], x[216], x[408], x[3], x[407], x[406]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[111], x[110], x[109], x[207], x[206], x[205], x[399], x[398], x[397], x[117], x[116], x[115], x[114], x[113], x[112], x[213], x[212], x[211], x[210], x[209], x[208], x[405], x[404], x[403], x[402], x[401], x[400], x[108], x[107], x[106], x[204], x[203], x[202], x[396], x[395], x[394], x[123], x[219], x[411], x[27], x[26], x[25], x[3], x[410], x[409]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[111], x[110], x[109], x[207], x[206], x[205], x[399], x[398], x[397], x[117], x[116], x[115], x[114], x[113], x[112], x[213], x[212], x[211], x[210], x[209], x[208], x[405], x[404], x[403], x[402], x[401], x[400], x[108], x[107], x[106], x[204], x[203], x[202], x[396], x[395], x[394], x[123], x[219], x[411], x[27], x[26], x[25], x[3], x[410], x[409]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[111], x[110], x[109], x[207], x[206], x[205], x[399], x[398], x[397], x[117], x[116], x[115], x[114], x[113], x[112], x[213], x[212], x[211], x[210], x[209], x[208], x[405], x[404], x[403], x[402], x[401], x[400], x[108], x[107], x[106], x[204], x[203], x[202], x[396], x[395], x[394], x[27], x[26], x[25], x[126], x[222], x[414], x[3], x[413], x[412]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[111], x[110], x[109], x[207], x[206], x[205], x[399], x[398], x[397], x[117], x[116], x[115], x[114], x[113], x[112], x[213], x[212], x[211], x[210], x[209], x[208], x[405], x[404], x[403], x[402], x[401], x[400], x[108], x[107], x[106], x[204], x[203], x[202], x[396], x[395], x[394], x[27], x[26], x[25], x[126], x[222], x[414], x[3], x[413], x[412]}), .y(y[149]));
endmodule

