////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module SkinnyTop in file /AGEMA/Designs/Skinny64_64_round-based/AGEMA/SkinnyTop.v */
/* clock gating is added to the circuit, the latency increased 2 time(s)  */

module SkinnyTop_HPC3_ClockGating_d3 (Plaintext_s0, Key_s0, clk, rst, Key_s1, Key_s2, Key_s3, Plaintext_s1, Plaintext_s2, Plaintext_s3, Fresh, Ciphertext_s0, done, Ciphertext_s1, Ciphertext_s2, Ciphertext_s3, Synch);
    input [63:0] Plaintext_s0 ;
    input [63:0] Key_s0 ;
    input clk ;
    input rst ;
    input [63:0] Key_s1 ;
    input [63:0] Key_s2 ;
    input [63:0] Key_s3 ;
    input [63:0] Plaintext_s1 ;
    input [63:0] Plaintext_s2 ;
    input [63:0] Plaintext_s3 ;
    input [767:0] Fresh ;
    output [63:0] Ciphertext_s0 ;
    output done ;
    output [63:0] Ciphertext_s1 ;
    output [63:0] Ciphertext_s2 ;
    output [63:0] Ciphertext_s3 ;
    output Synch ;
    wire SubCellInst_SboxInst_0_n3 ;
    wire SubCellInst_SboxInst_0_YY_0_ ;
    wire SubCellInst_SboxInst_0_YY_1_ ;
    wire SubCellInst_SboxInst_0_L3 ;
    wire SubCellInst_SboxInst_0_YY_3 ;
    wire SubCellInst_SboxInst_0_L2 ;
    wire SubCellInst_SboxInst_0_T3 ;
    wire SubCellInst_SboxInst_0_Q7 ;
    wire SubCellInst_SboxInst_0_L1 ;
    wire SubCellInst_SboxInst_0_Q6 ;
    wire SubCellInst_SboxInst_0_L0 ;
    wire SubCellInst_SboxInst_0_T2 ;
    wire SubCellInst_SboxInst_0_Q4 ;
    wire SubCellInst_SboxInst_0_T1 ;
    wire SubCellInst_SboxInst_0_Q2 ;
    wire SubCellInst_SboxInst_0_T0 ;
    wire SubCellInst_SboxInst_0_Q1 ;
    wire SubCellInst_SboxInst_0_Q0 ;
    wire SubCellInst_SboxInst_0_XX_1_ ;
    wire SubCellInst_SboxInst_0_XX_2_ ;
    wire SubCellInst_SboxInst_1_n3 ;
    wire SubCellInst_SboxInst_1_YY_0_ ;
    wire SubCellInst_SboxInst_1_YY_1_ ;
    wire SubCellInst_SboxInst_1_L3 ;
    wire SubCellInst_SboxInst_1_YY_3 ;
    wire SubCellInst_SboxInst_1_L2 ;
    wire SubCellInst_SboxInst_1_T3 ;
    wire SubCellInst_SboxInst_1_Q7 ;
    wire SubCellInst_SboxInst_1_L1 ;
    wire SubCellInst_SboxInst_1_Q6 ;
    wire SubCellInst_SboxInst_1_L0 ;
    wire SubCellInst_SboxInst_1_T2 ;
    wire SubCellInst_SboxInst_1_Q4 ;
    wire SubCellInst_SboxInst_1_T1 ;
    wire SubCellInst_SboxInst_1_Q2 ;
    wire SubCellInst_SboxInst_1_T0 ;
    wire SubCellInst_SboxInst_1_Q1 ;
    wire SubCellInst_SboxInst_1_Q0 ;
    wire SubCellInst_SboxInst_1_XX_1_ ;
    wire SubCellInst_SboxInst_1_XX_2_ ;
    wire SubCellInst_SboxInst_2_n3 ;
    wire SubCellInst_SboxInst_2_YY_0_ ;
    wire SubCellInst_SboxInst_2_YY_1_ ;
    wire SubCellInst_SboxInst_2_L3 ;
    wire SubCellInst_SboxInst_2_YY_3 ;
    wire SubCellInst_SboxInst_2_L2 ;
    wire SubCellInst_SboxInst_2_T3 ;
    wire SubCellInst_SboxInst_2_Q7 ;
    wire SubCellInst_SboxInst_2_L1 ;
    wire SubCellInst_SboxInst_2_Q6 ;
    wire SubCellInst_SboxInst_2_L0 ;
    wire SubCellInst_SboxInst_2_T2 ;
    wire SubCellInst_SboxInst_2_Q4 ;
    wire SubCellInst_SboxInst_2_T1 ;
    wire SubCellInst_SboxInst_2_Q2 ;
    wire SubCellInst_SboxInst_2_T0 ;
    wire SubCellInst_SboxInst_2_Q1 ;
    wire SubCellInst_SboxInst_2_Q0 ;
    wire SubCellInst_SboxInst_2_XX_1_ ;
    wire SubCellInst_SboxInst_2_XX_2_ ;
    wire SubCellInst_SboxInst_3_n3 ;
    wire SubCellInst_SboxInst_3_YY_0_ ;
    wire SubCellInst_SboxInst_3_YY_1_ ;
    wire SubCellInst_SboxInst_3_L3 ;
    wire SubCellInst_SboxInst_3_YY_3 ;
    wire SubCellInst_SboxInst_3_L2 ;
    wire SubCellInst_SboxInst_3_T3 ;
    wire SubCellInst_SboxInst_3_Q7 ;
    wire SubCellInst_SboxInst_3_L1 ;
    wire SubCellInst_SboxInst_3_Q6 ;
    wire SubCellInst_SboxInst_3_L0 ;
    wire SubCellInst_SboxInst_3_T2 ;
    wire SubCellInst_SboxInst_3_Q4 ;
    wire SubCellInst_SboxInst_3_T1 ;
    wire SubCellInst_SboxInst_3_Q2 ;
    wire SubCellInst_SboxInst_3_T0 ;
    wire SubCellInst_SboxInst_3_Q1 ;
    wire SubCellInst_SboxInst_3_Q0 ;
    wire SubCellInst_SboxInst_3_XX_1_ ;
    wire SubCellInst_SboxInst_3_XX_2_ ;
    wire SubCellInst_SboxInst_4_n3 ;
    wire SubCellInst_SboxInst_4_YY_0_ ;
    wire SubCellInst_SboxInst_4_YY_1_ ;
    wire SubCellInst_SboxInst_4_L3 ;
    wire SubCellInst_SboxInst_4_YY_3 ;
    wire SubCellInst_SboxInst_4_L2 ;
    wire SubCellInst_SboxInst_4_T3 ;
    wire SubCellInst_SboxInst_4_Q7 ;
    wire SubCellInst_SboxInst_4_L1 ;
    wire SubCellInst_SboxInst_4_Q6 ;
    wire SubCellInst_SboxInst_4_L0 ;
    wire SubCellInst_SboxInst_4_T2 ;
    wire SubCellInst_SboxInst_4_Q4 ;
    wire SubCellInst_SboxInst_4_T1 ;
    wire SubCellInst_SboxInst_4_Q2 ;
    wire SubCellInst_SboxInst_4_T0 ;
    wire SubCellInst_SboxInst_4_Q1 ;
    wire SubCellInst_SboxInst_4_Q0 ;
    wire SubCellInst_SboxInst_4_XX_1_ ;
    wire SubCellInst_SboxInst_4_XX_2_ ;
    wire SubCellInst_SboxInst_5_n3 ;
    wire SubCellInst_SboxInst_5_YY_0_ ;
    wire SubCellInst_SboxInst_5_YY_1_ ;
    wire SubCellInst_SboxInst_5_L3 ;
    wire SubCellInst_SboxInst_5_YY_3 ;
    wire SubCellInst_SboxInst_5_L2 ;
    wire SubCellInst_SboxInst_5_T3 ;
    wire SubCellInst_SboxInst_5_Q7 ;
    wire SubCellInst_SboxInst_5_L1 ;
    wire SubCellInst_SboxInst_5_Q6 ;
    wire SubCellInst_SboxInst_5_L0 ;
    wire SubCellInst_SboxInst_5_T2 ;
    wire SubCellInst_SboxInst_5_Q4 ;
    wire SubCellInst_SboxInst_5_T1 ;
    wire SubCellInst_SboxInst_5_Q2 ;
    wire SubCellInst_SboxInst_5_T0 ;
    wire SubCellInst_SboxInst_5_Q1 ;
    wire SubCellInst_SboxInst_5_Q0 ;
    wire SubCellInst_SboxInst_5_XX_1_ ;
    wire SubCellInst_SboxInst_5_XX_2_ ;
    wire SubCellInst_SboxInst_6_n3 ;
    wire SubCellInst_SboxInst_6_YY_0_ ;
    wire SubCellInst_SboxInst_6_YY_1_ ;
    wire SubCellInst_SboxInst_6_L3 ;
    wire SubCellInst_SboxInst_6_YY_3 ;
    wire SubCellInst_SboxInst_6_L2 ;
    wire SubCellInst_SboxInst_6_T3 ;
    wire SubCellInst_SboxInst_6_Q7 ;
    wire SubCellInst_SboxInst_6_L1 ;
    wire SubCellInst_SboxInst_6_Q6 ;
    wire SubCellInst_SboxInst_6_L0 ;
    wire SubCellInst_SboxInst_6_T2 ;
    wire SubCellInst_SboxInst_6_Q4 ;
    wire SubCellInst_SboxInst_6_T1 ;
    wire SubCellInst_SboxInst_6_Q2 ;
    wire SubCellInst_SboxInst_6_T0 ;
    wire SubCellInst_SboxInst_6_Q1 ;
    wire SubCellInst_SboxInst_6_Q0 ;
    wire SubCellInst_SboxInst_6_XX_1_ ;
    wire SubCellInst_SboxInst_6_XX_2_ ;
    wire SubCellInst_SboxInst_7_n3 ;
    wire SubCellInst_SboxInst_7_YY_0_ ;
    wire SubCellInst_SboxInst_7_YY_1_ ;
    wire SubCellInst_SboxInst_7_L3 ;
    wire SubCellInst_SboxInst_7_YY_3 ;
    wire SubCellInst_SboxInst_7_L2 ;
    wire SubCellInst_SboxInst_7_T3 ;
    wire SubCellInst_SboxInst_7_Q7 ;
    wire SubCellInst_SboxInst_7_L1 ;
    wire SubCellInst_SboxInst_7_Q6 ;
    wire SubCellInst_SboxInst_7_L0 ;
    wire SubCellInst_SboxInst_7_T2 ;
    wire SubCellInst_SboxInst_7_Q4 ;
    wire SubCellInst_SboxInst_7_T1 ;
    wire SubCellInst_SboxInst_7_Q2 ;
    wire SubCellInst_SboxInst_7_T0 ;
    wire SubCellInst_SboxInst_7_Q1 ;
    wire SubCellInst_SboxInst_7_Q0 ;
    wire SubCellInst_SboxInst_7_XX_1_ ;
    wire SubCellInst_SboxInst_7_XX_2_ ;
    wire SubCellInst_SboxInst_8_n3 ;
    wire SubCellInst_SboxInst_8_YY_0_ ;
    wire SubCellInst_SboxInst_8_YY_1_ ;
    wire SubCellInst_SboxInst_8_L3 ;
    wire SubCellInst_SboxInst_8_YY_3 ;
    wire SubCellInst_SboxInst_8_L2 ;
    wire SubCellInst_SboxInst_8_T3 ;
    wire SubCellInst_SboxInst_8_Q7 ;
    wire SubCellInst_SboxInst_8_L1 ;
    wire SubCellInst_SboxInst_8_Q6 ;
    wire SubCellInst_SboxInst_8_L0 ;
    wire SubCellInst_SboxInst_8_T2 ;
    wire SubCellInst_SboxInst_8_Q4 ;
    wire SubCellInst_SboxInst_8_T1 ;
    wire SubCellInst_SboxInst_8_Q2 ;
    wire SubCellInst_SboxInst_8_T0 ;
    wire SubCellInst_SboxInst_8_Q1 ;
    wire SubCellInst_SboxInst_8_Q0 ;
    wire SubCellInst_SboxInst_8_XX_1_ ;
    wire SubCellInst_SboxInst_8_XX_2_ ;
    wire SubCellInst_SboxInst_9_n3 ;
    wire SubCellInst_SboxInst_9_YY_0_ ;
    wire SubCellInst_SboxInst_9_YY_1_ ;
    wire SubCellInst_SboxInst_9_L3 ;
    wire SubCellInst_SboxInst_9_YY_3 ;
    wire SubCellInst_SboxInst_9_L2 ;
    wire SubCellInst_SboxInst_9_T3 ;
    wire SubCellInst_SboxInst_9_Q7 ;
    wire SubCellInst_SboxInst_9_L1 ;
    wire SubCellInst_SboxInst_9_Q6 ;
    wire SubCellInst_SboxInst_9_L0 ;
    wire SubCellInst_SboxInst_9_T2 ;
    wire SubCellInst_SboxInst_9_Q4 ;
    wire SubCellInst_SboxInst_9_T1 ;
    wire SubCellInst_SboxInst_9_Q2 ;
    wire SubCellInst_SboxInst_9_T0 ;
    wire SubCellInst_SboxInst_9_Q1 ;
    wire SubCellInst_SboxInst_9_Q0 ;
    wire SubCellInst_SboxInst_9_XX_1_ ;
    wire SubCellInst_SboxInst_9_XX_2_ ;
    wire SubCellInst_SboxInst_10_n3 ;
    wire SubCellInst_SboxInst_10_YY_0_ ;
    wire SubCellInst_SboxInst_10_YY_1_ ;
    wire SubCellInst_SboxInst_10_L3 ;
    wire SubCellInst_SboxInst_10_YY_3 ;
    wire SubCellInst_SboxInst_10_L2 ;
    wire SubCellInst_SboxInst_10_T3 ;
    wire SubCellInst_SboxInst_10_Q7 ;
    wire SubCellInst_SboxInst_10_L1 ;
    wire SubCellInst_SboxInst_10_Q6 ;
    wire SubCellInst_SboxInst_10_L0 ;
    wire SubCellInst_SboxInst_10_T2 ;
    wire SubCellInst_SboxInst_10_Q4 ;
    wire SubCellInst_SboxInst_10_T1 ;
    wire SubCellInst_SboxInst_10_Q2 ;
    wire SubCellInst_SboxInst_10_T0 ;
    wire SubCellInst_SboxInst_10_Q1 ;
    wire SubCellInst_SboxInst_10_Q0 ;
    wire SubCellInst_SboxInst_10_XX_1_ ;
    wire SubCellInst_SboxInst_10_XX_2_ ;
    wire SubCellInst_SboxInst_11_n3 ;
    wire SubCellInst_SboxInst_11_YY_0_ ;
    wire SubCellInst_SboxInst_11_YY_1_ ;
    wire SubCellInst_SboxInst_11_L3 ;
    wire SubCellInst_SboxInst_11_YY_3 ;
    wire SubCellInst_SboxInst_11_L2 ;
    wire SubCellInst_SboxInst_11_T3 ;
    wire SubCellInst_SboxInst_11_Q7 ;
    wire SubCellInst_SboxInst_11_L1 ;
    wire SubCellInst_SboxInst_11_Q6 ;
    wire SubCellInst_SboxInst_11_L0 ;
    wire SubCellInst_SboxInst_11_T2 ;
    wire SubCellInst_SboxInst_11_Q4 ;
    wire SubCellInst_SboxInst_11_T1 ;
    wire SubCellInst_SboxInst_11_Q2 ;
    wire SubCellInst_SboxInst_11_T0 ;
    wire SubCellInst_SboxInst_11_Q1 ;
    wire SubCellInst_SboxInst_11_Q0 ;
    wire SubCellInst_SboxInst_11_XX_1_ ;
    wire SubCellInst_SboxInst_11_XX_2_ ;
    wire SubCellInst_SboxInst_12_n3 ;
    wire SubCellInst_SboxInst_12_YY_0_ ;
    wire SubCellInst_SboxInst_12_YY_1_ ;
    wire SubCellInst_SboxInst_12_L3 ;
    wire SubCellInst_SboxInst_12_YY_3 ;
    wire SubCellInst_SboxInst_12_L2 ;
    wire SubCellInst_SboxInst_12_T3 ;
    wire SubCellInst_SboxInst_12_Q7 ;
    wire SubCellInst_SboxInst_12_L1 ;
    wire SubCellInst_SboxInst_12_Q6 ;
    wire SubCellInst_SboxInst_12_L0 ;
    wire SubCellInst_SboxInst_12_T2 ;
    wire SubCellInst_SboxInst_12_Q4 ;
    wire SubCellInst_SboxInst_12_T1 ;
    wire SubCellInst_SboxInst_12_Q2 ;
    wire SubCellInst_SboxInst_12_T0 ;
    wire SubCellInst_SboxInst_12_Q1 ;
    wire SubCellInst_SboxInst_12_Q0 ;
    wire SubCellInst_SboxInst_12_XX_1_ ;
    wire SubCellInst_SboxInst_12_XX_2_ ;
    wire SubCellInst_SboxInst_13_n3 ;
    wire SubCellInst_SboxInst_13_YY_0_ ;
    wire SubCellInst_SboxInst_13_YY_1_ ;
    wire SubCellInst_SboxInst_13_L3 ;
    wire SubCellInst_SboxInst_13_YY_3 ;
    wire SubCellInst_SboxInst_13_L2 ;
    wire SubCellInst_SboxInst_13_T3 ;
    wire SubCellInst_SboxInst_13_Q7 ;
    wire SubCellInst_SboxInst_13_L1 ;
    wire SubCellInst_SboxInst_13_Q6 ;
    wire SubCellInst_SboxInst_13_L0 ;
    wire SubCellInst_SboxInst_13_T2 ;
    wire SubCellInst_SboxInst_13_Q4 ;
    wire SubCellInst_SboxInst_13_T1 ;
    wire SubCellInst_SboxInst_13_Q2 ;
    wire SubCellInst_SboxInst_13_T0 ;
    wire SubCellInst_SboxInst_13_Q1 ;
    wire SubCellInst_SboxInst_13_Q0 ;
    wire SubCellInst_SboxInst_13_XX_1_ ;
    wire SubCellInst_SboxInst_13_XX_2_ ;
    wire SubCellInst_SboxInst_14_n3 ;
    wire SubCellInst_SboxInst_14_YY_0_ ;
    wire SubCellInst_SboxInst_14_YY_1_ ;
    wire SubCellInst_SboxInst_14_L3 ;
    wire SubCellInst_SboxInst_14_YY_3 ;
    wire SubCellInst_SboxInst_14_L2 ;
    wire SubCellInst_SboxInst_14_T3 ;
    wire SubCellInst_SboxInst_14_Q7 ;
    wire SubCellInst_SboxInst_14_L1 ;
    wire SubCellInst_SboxInst_14_Q6 ;
    wire SubCellInst_SboxInst_14_L0 ;
    wire SubCellInst_SboxInst_14_T2 ;
    wire SubCellInst_SboxInst_14_Q4 ;
    wire SubCellInst_SboxInst_14_T1 ;
    wire SubCellInst_SboxInst_14_Q2 ;
    wire SubCellInst_SboxInst_14_T0 ;
    wire SubCellInst_SboxInst_14_Q1 ;
    wire SubCellInst_SboxInst_14_Q0 ;
    wire SubCellInst_SboxInst_14_XX_1_ ;
    wire SubCellInst_SboxInst_14_XX_2_ ;
    wire SubCellInst_SboxInst_15_n3 ;
    wire SubCellInst_SboxInst_15_YY_0_ ;
    wire SubCellInst_SboxInst_15_YY_1_ ;
    wire SubCellInst_SboxInst_15_L3 ;
    wire SubCellInst_SboxInst_15_YY_3 ;
    wire SubCellInst_SboxInst_15_L2 ;
    wire SubCellInst_SboxInst_15_T3 ;
    wire SubCellInst_SboxInst_15_Q7 ;
    wire SubCellInst_SboxInst_15_L1 ;
    wire SubCellInst_SboxInst_15_Q6 ;
    wire SubCellInst_SboxInst_15_L0 ;
    wire SubCellInst_SboxInst_15_T2 ;
    wire SubCellInst_SboxInst_15_Q4 ;
    wire SubCellInst_SboxInst_15_T1 ;
    wire SubCellInst_SboxInst_15_Q2 ;
    wire SubCellInst_SboxInst_15_T0 ;
    wire SubCellInst_SboxInst_15_Q1 ;
    wire SubCellInst_SboxInst_15_Q0 ;
    wire SubCellInst_SboxInst_15_XX_1_ ;
    wire SubCellInst_SboxInst_15_XX_2_ ;
    wire AddConstXOR_AddConstXOR_XORInst_0_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_0_3_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_0_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_1_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_2_n1 ;
    wire AddConstXOR_AddConstXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_0_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_1_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_2_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_3_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_4_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_5_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_6_3_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_0_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_1_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_2_n1 ;
    wire AddRoundTweakeyXOR_XORInst_7_3_n1 ;
    wire MCInst_MCR0_XORInst_0_0_n2 ;
    wire MCInst_MCR0_XORInst_0_0_n1 ;
    wire MCInst_MCR0_XORInst_0_1_n2 ;
    wire MCInst_MCR0_XORInst_0_1_n1 ;
    wire MCInst_MCR0_XORInst_0_2_n2 ;
    wire MCInst_MCR0_XORInst_0_2_n1 ;
    wire MCInst_MCR0_XORInst_0_3_n2 ;
    wire MCInst_MCR0_XORInst_0_3_n1 ;
    wire MCInst_MCR0_XORInst_1_0_n2 ;
    wire MCInst_MCR0_XORInst_1_0_n1 ;
    wire MCInst_MCR0_XORInst_1_1_n2 ;
    wire MCInst_MCR0_XORInst_1_1_n1 ;
    wire MCInst_MCR0_XORInst_1_2_n2 ;
    wire MCInst_MCR0_XORInst_1_2_n1 ;
    wire MCInst_MCR0_XORInst_1_3_n2 ;
    wire MCInst_MCR0_XORInst_1_3_n1 ;
    wire MCInst_MCR0_XORInst_2_0_n2 ;
    wire MCInst_MCR0_XORInst_2_0_n1 ;
    wire MCInst_MCR0_XORInst_2_1_n2 ;
    wire MCInst_MCR0_XORInst_2_1_n1 ;
    wire MCInst_MCR0_XORInst_2_2_n2 ;
    wire MCInst_MCR0_XORInst_2_2_n1 ;
    wire MCInst_MCR0_XORInst_2_3_n2 ;
    wire MCInst_MCR0_XORInst_2_3_n1 ;
    wire MCInst_MCR0_XORInst_3_0_n2 ;
    wire MCInst_MCR0_XORInst_3_0_n1 ;
    wire MCInst_MCR0_XORInst_3_1_n2 ;
    wire MCInst_MCR0_XORInst_3_1_n1 ;
    wire MCInst_MCR0_XORInst_3_2_n2 ;
    wire MCInst_MCR0_XORInst_3_2_n1 ;
    wire MCInst_MCR0_XORInst_3_3_n2 ;
    wire MCInst_MCR0_XORInst_3_3_n1 ;
    wire MCInst_MCR2_XORInst_0_0_n1 ;
    wire MCInst_MCR2_XORInst_0_1_n1 ;
    wire MCInst_MCR2_XORInst_0_2_n1 ;
    wire MCInst_MCR2_XORInst_0_3_n1 ;
    wire MCInst_MCR2_XORInst_1_0_n1 ;
    wire MCInst_MCR2_XORInst_1_1_n1 ;
    wire MCInst_MCR2_XORInst_1_2_n1 ;
    wire MCInst_MCR2_XORInst_1_3_n1 ;
    wire MCInst_MCR2_XORInst_2_0_n1 ;
    wire MCInst_MCR2_XORInst_2_1_n1 ;
    wire MCInst_MCR2_XORInst_2_2_n1 ;
    wire MCInst_MCR2_XORInst_2_3_n1 ;
    wire MCInst_MCR2_XORInst_3_0_n1 ;
    wire MCInst_MCR2_XORInst_3_1_n1 ;
    wire MCInst_MCR2_XORInst_3_2_n1 ;
    wire MCInst_MCR2_XORInst_3_3_n1 ;
    wire MCInst_MCR3_XORInst_0_0_n1 ;
    wire MCInst_MCR3_XORInst_0_1_n1 ;
    wire MCInst_MCR3_XORInst_0_2_n1 ;
    wire MCInst_MCR3_XORInst_0_3_n1 ;
    wire MCInst_MCR3_XORInst_1_0_n1 ;
    wire MCInst_MCR3_XORInst_1_1_n1 ;
    wire MCInst_MCR3_XORInst_1_2_n1 ;
    wire MCInst_MCR3_XORInst_1_3_n1 ;
    wire MCInst_MCR3_XORInst_2_0_n1 ;
    wire MCInst_MCR3_XORInst_2_1_n1 ;
    wire MCInst_MCR3_XORInst_2_2_n1 ;
    wire MCInst_MCR3_XORInst_2_3_n1 ;
    wire MCInst_MCR3_XORInst_3_0_n1 ;
    wire MCInst_MCR3_XORInst_3_1_n1 ;
    wire MCInst_MCR3_XORInst_3_2_n1 ;
    wire MCInst_MCR3_XORInst_3_3_n1 ;
    wire FSMUpdateInst_StateUpdateInst_0_n4 ;
    wire FSMUpdateInst_StateUpdateInst_0_n3 ;
    wire FSMUpdateInst_StateUpdateInst_0_n2 ;
    wire FSMUpdateInst_StateUpdateInst_0_n1 ;
    wire FSMUpdateInst_StateUpdateInst_2_n4 ;
    wire FSMUpdateInst_StateUpdateInst_2_n3 ;
    wire FSMUpdateInst_StateUpdateInst_2_n2 ;
    wire FSMUpdateInst_StateUpdateInst_2_n1 ;
    wire FSMUpdateInst_StateUpdateInst_5_n4 ;
    wire FSMUpdateInst_StateUpdateInst_5_n3 ;
    wire FSMUpdateInst_StateUpdateInst_5_n2 ;
    wire FSMUpdateInst_StateUpdateInst_5_n1 ;
    wire FSMSignalsInst_doneInst_n5 ;
    wire FSMSignalsInst_doneInst_n4 ;
    wire FSMSignalsInst_doneInst_n3 ;
    wire FSMSignalsInst_doneInst_n2 ;
    wire FSMSignalsInst_doneInst_n1 ;
    wire [63:0] MCOutput ;
    wire [63:0] StateRegInput ;
    wire [63:29] SubCellOutput ;
    wire [5:1] FSM ;
    wire [63:32] AddRoundConstantOutput ;
    wire [47:0] ShiftRowsOutput ;
    wire [5:0] FSMUpdate ;
    wire [5:0] FSMSelected ;
    wire [63:0] TweakeyGeneration_StateRegInput ;
    wire [63:0] TweakeyGeneration_key_Feedback ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2494 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2512 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2530 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2548 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2566 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U1 ( .a ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR_i1_U1 ( .a ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .b ({Ciphertext_s3[3], Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}), .c ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_0_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR_i2_U1 ( .a ({Ciphertext_s3[0], Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}), .b ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}), .c ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR0_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, SubCellInst_SboxInst_0_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR1_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_0_XX_1_}), .c ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR3_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, SubCellInst_SboxInst_0_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR5_U1 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_0_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR6_U1 ( .a ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_Q1}), .b ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_0_Q6}), .c ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_0_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR8_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, SubCellInst_SboxInst_0_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U1 ( .a ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR_i1_U1 ( .a ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .b ({Ciphertext_s3[7], Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}), .c ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_1_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR_i2_U1 ( .a ({Ciphertext_s3[4], Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}), .b ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}), .c ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR0_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}), .c ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, SubCellInst_SboxInst_1_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR1_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_1_XX_1_}), .c ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_1_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR3_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, SubCellInst_SboxInst_1_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR5_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_1_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR6_U1 ( .a ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_1_Q1}), .b ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_1_Q6}), .c ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, SubCellInst_SboxInst_1_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR8_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .c ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, SubCellInst_SboxInst_1_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U1 ( .a ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR_i1_U1 ( .a ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .b ({Ciphertext_s3[11], Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}), .c ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_2_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR_i2_U1 ( .a ({Ciphertext_s3[8], Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}), .b ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}), .c ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR0_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}), .c ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, SubCellInst_SboxInst_2_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR1_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_2_XX_1_}), .c ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_2_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR3_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, SubCellInst_SboxInst_2_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR5_U1 ( .a ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_2_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR6_U1 ( .a ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_2_Q1}), .b ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_2_Q6}), .c ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, SubCellInst_SboxInst_2_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR8_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .c ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, SubCellInst_SboxInst_2_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U1 ( .a ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR_i1_U1 ( .a ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .b ({Ciphertext_s3[15], Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}), .c ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_3_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR_i2_U1 ( .a ({Ciphertext_s3[12], Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}), .b ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}), .c ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR0_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}), .c ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, SubCellInst_SboxInst_3_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR1_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_3_XX_1_}), .c ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_3_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR3_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, SubCellInst_SboxInst_3_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR5_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_3_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR6_U1 ( .a ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_3_Q1}), .b ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_3_Q6}), .c ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, SubCellInst_SboxInst_3_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR8_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .c ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, SubCellInst_SboxInst_3_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U1 ( .a ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR_i1_U1 ( .a ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .b ({Ciphertext_s3[19], Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}), .c ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_4_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR_i2_U1 ( .a ({Ciphertext_s3[16], Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}), .b ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}), .c ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR0_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}), .c ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, SubCellInst_SboxInst_4_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR1_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_4_XX_1_}), .c ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_4_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR3_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, SubCellInst_SboxInst_4_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR5_U1 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_4_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR6_U1 ( .a ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_4_Q1}), .b ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_4_Q6}), .c ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, SubCellInst_SboxInst_4_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR8_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, SubCellInst_SboxInst_4_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U1 ( .a ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR_i1_U1 ( .a ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .b ({Ciphertext_s3[23], Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}), .c ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_5_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR_i2_U1 ( .a ({Ciphertext_s3[20], Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}), .b ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}), .c ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR0_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}), .c ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, SubCellInst_SboxInst_5_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR1_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_5_XX_1_}), .c ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_5_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR3_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, SubCellInst_SboxInst_5_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR5_U1 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_5_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR6_U1 ( .a ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_5_Q1}), .b ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_5_Q6}), .c ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, SubCellInst_SboxInst_5_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR8_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .c ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, SubCellInst_SboxInst_5_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U1 ( .a ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR_i1_U1 ( .a ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .b ({Ciphertext_s3[27], Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}), .c ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_6_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR_i2_U1 ( .a ({Ciphertext_s3[24], Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}), .b ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}), .c ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR0_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}), .c ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, SubCellInst_SboxInst_6_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR1_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_6_XX_1_}), .c ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_6_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR3_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, SubCellInst_SboxInst_6_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR5_U1 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_6_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR6_U1 ( .a ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_6_Q1}), .b ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_6_Q6}), .c ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_6_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR8_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, SubCellInst_SboxInst_6_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U1 ( .a ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR_i1_U1 ( .a ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .b ({Ciphertext_s3[31], Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}), .c ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_7_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR_i2_U1 ( .a ({Ciphertext_s3[28], Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}), .b ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}), .c ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR0_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, SubCellInst_SboxInst_7_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR1_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_7_XX_1_}), .c ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_7_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR3_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, SubCellInst_SboxInst_7_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR5_U1 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_7_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR6_U1 ( .a ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_7_Q1}), .b ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_7_Q6}), .c ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, SubCellInst_SboxInst_7_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR8_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, SubCellInst_SboxInst_7_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U1 ( .a ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR_i1_U1 ( .a ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .b ({Ciphertext_s3[35], Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}), .c ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_8_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR_i2_U1 ( .a ({Ciphertext_s3[32], Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}), .b ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}), .c ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR0_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, SubCellInst_SboxInst_8_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR1_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_8_XX_1_}), .c ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_8_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR3_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, SubCellInst_SboxInst_8_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR5_U1 ( .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_8_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR6_U1 ( .a ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_8_Q1}), .b ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_8_Q6}), .c ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, SubCellInst_SboxInst_8_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR8_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, SubCellInst_SboxInst_8_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U1 ( .a ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR_i1_U1 ( .a ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .b ({Ciphertext_s3[39], Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}), .c ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_9_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR_i2_U1 ( .a ({Ciphertext_s3[36], Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}), .b ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}), .c ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR0_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, SubCellInst_SboxInst_9_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR1_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_9_XX_1_}), .c ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, SubCellInst_SboxInst_9_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR3_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, SubCellInst_SboxInst_9_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR5_U1 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_9_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR6_U1 ( .a ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, SubCellInst_SboxInst_9_Q1}), .b ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_9_Q6}), .c ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, SubCellInst_SboxInst_9_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR8_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, SubCellInst_SboxInst_9_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U1 ( .a ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR_i1_U1 ( .a ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .b ({Ciphertext_s3[43], Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}), .c ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_10_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR_i2_U1 ( .a ({Ciphertext_s3[40], Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}), .b ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}), .c ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR0_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, SubCellInst_SboxInst_10_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR1_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_10_XX_1_}), .c ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_10_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR3_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, SubCellInst_SboxInst_10_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR5_U1 ( .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, SubCellInst_SboxInst_10_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR6_U1 ( .a ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_10_Q1}), .b ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, SubCellInst_SboxInst_10_Q6}), .c ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR8_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, SubCellInst_SboxInst_10_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U1 ( .a ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR_i1_U1 ( .a ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .b ({Ciphertext_s3[47], Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}), .c ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_11_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR_i2_U1 ( .a ({Ciphertext_s3[44], Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}), .b ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}), .c ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR0_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, SubCellInst_SboxInst_11_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR1_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_11_XX_1_}), .c ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_11_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR3_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, SubCellInst_SboxInst_11_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR5_U1 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_11_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR6_U1 ( .a ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_11_Q1}), .b ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_11_Q6}), .c ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, SubCellInst_SboxInst_11_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR8_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, SubCellInst_SboxInst_11_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U1 ( .a ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR_i1_U1 ( .a ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .b ({Ciphertext_s3[51], Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}), .c ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_12_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR_i2_U1 ( .a ({Ciphertext_s3[48], Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}), .b ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}), .c ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR0_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, SubCellInst_SboxInst_12_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR1_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_12_XX_1_}), .c ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_12_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR3_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, SubCellInst_SboxInst_12_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR5_U1 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR6_U1 ( .a ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_12_Q1}), .b ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_Q6}), .c ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, SubCellInst_SboxInst_12_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR8_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, SubCellInst_SboxInst_12_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U1 ( .a ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR_i1_U1 ( .a ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .b ({Ciphertext_s3[55], Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}), .c ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_13_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR_i2_U1 ( .a ({Ciphertext_s3[52], Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}), .b ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}), .c ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR0_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, SubCellInst_SboxInst_13_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR1_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_13_XX_1_}), .c ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, SubCellInst_SboxInst_13_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR3_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, SubCellInst_SboxInst_13_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR5_U1 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_13_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR6_U1 ( .a ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, SubCellInst_SboxInst_13_Q1}), .b ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_13_Q6}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, SubCellInst_SboxInst_13_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR8_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, SubCellInst_SboxInst_13_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U1 ( .a ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR_i1_U1 ( .a ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .b ({Ciphertext_s3[59], Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}), .c ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_14_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR_i2_U1 ( .a ({Ciphertext_s3[56], Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}), .b ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}), .c ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR0_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, SubCellInst_SboxInst_14_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR1_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_14_XX_1_}), .c ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_14_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR3_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, SubCellInst_SboxInst_14_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR5_U1 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, SubCellInst_SboxInst_14_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR6_U1 ( .a ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_14_Q1}), .b ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, SubCellInst_SboxInst_14_Q6}), .c ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, SubCellInst_SboxInst_14_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR8_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, SubCellInst_SboxInst_14_L2}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U1 ( .a ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR_i1_U1 ( .a ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .b ({Ciphertext_s3[63], Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}), .c ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_15_XX_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR_i2_U1 ( .a ({Ciphertext_s3[60], Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}), .b ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}), .c ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR0_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, SubCellInst_SboxInst_15_Q0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR1_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_15_XX_1_}), .c ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, SubCellInst_SboxInst_15_Q1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR3_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, SubCellInst_SboxInst_15_Q4}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR5_U1 ( .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_15_Q6}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR6_U1 ( .a ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, SubCellInst_SboxInst_15_Q1}), .b ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_15_Q6}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, SubCellInst_SboxInst_15_L1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR8_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, SubCellInst_SboxInst_15_L2}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[0]}), .a ({Key_s3[0], Key_s2[0], Key_s1[0], Key_s0[0]}), .c ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, TweakeyGeneration_key_Feedback[1]}), .a ({Key_s3[1], Key_s2[1], Key_s1[1], Key_s0[1]}), .c ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, TweakeyGeneration_StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[2]}), .a ({Key_s3[2], Key_s2[2], Key_s1[2], Key_s0[2]}), .c ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, TweakeyGeneration_key_Feedback[3]}), .a ({Key_s3[3], Key_s2[3], Key_s1[3], Key_s0[3]}), .c ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, TweakeyGeneration_StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[4]}), .a ({Key_s3[4], Key_s2[4], Key_s1[4], Key_s0[4]}), .c ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, TweakeyGeneration_key_Feedback[5]}), .a ({Key_s3[5], Key_s2[5], Key_s1[5], Key_s0[5]}), .c ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, TweakeyGeneration_StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[6]}), .a ({Key_s3[6], Key_s2[6], Key_s1[6], Key_s0[6]}), .c ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, TweakeyGeneration_key_Feedback[7]}), .a ({Key_s3[7], Key_s2[7], Key_s1[7], Key_s0[7]}), .c ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, TweakeyGeneration_StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[8]}), .a ({Key_s3[8], Key_s2[8], Key_s1[8], Key_s0[8]}), .c ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, TweakeyGeneration_key_Feedback[9]}), .a ({Key_s3[9], Key_s2[9], Key_s1[9], Key_s0[9]}), .c ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, TweakeyGeneration_StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[10]}), .a ({Key_s3[10], Key_s2[10], Key_s1[10], Key_s0[10]}), .c ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, TweakeyGeneration_key_Feedback[11]}), .a ({Key_s3[11], Key_s2[11], Key_s1[11], Key_s0[11]}), .c ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, TweakeyGeneration_StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[12]}), .a ({Key_s3[12], Key_s2[12], Key_s1[12], Key_s0[12]}), .c ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, TweakeyGeneration_key_Feedback[13]}), .a ({Key_s3[13], Key_s2[13], Key_s1[13], Key_s0[13]}), .c ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, TweakeyGeneration_StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[14]}), .a ({Key_s3[14], Key_s2[14], Key_s1[14], Key_s0[14]}), .c ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, TweakeyGeneration_key_Feedback[15]}), .a ({Key_s3[15], Key_s2[15], Key_s1[15], Key_s0[15]}), .c ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, TweakeyGeneration_StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[16]}), .a ({Key_s3[16], Key_s2[16], Key_s1[16], Key_s0[16]}), .c ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, TweakeyGeneration_key_Feedback[17]}), .a ({Key_s3[17], Key_s2[17], Key_s1[17], Key_s0[17]}), .c ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, TweakeyGeneration_StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[18]}), .a ({Key_s3[18], Key_s2[18], Key_s1[18], Key_s0[18]}), .c ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, TweakeyGeneration_key_Feedback[19]}), .a ({Key_s3[19], Key_s2[19], Key_s1[19], Key_s0[19]}), .c ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, TweakeyGeneration_StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[20]}), .a ({Key_s3[20], Key_s2[20], Key_s1[20], Key_s0[20]}), .c ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, TweakeyGeneration_key_Feedback[21]}), .a ({Key_s3[21], Key_s2[21], Key_s1[21], Key_s0[21]}), .c ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, TweakeyGeneration_StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[22]}), .a ({Key_s3[22], Key_s2[22], Key_s1[22], Key_s0[22]}), .c ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, TweakeyGeneration_key_Feedback[23]}), .a ({Key_s3[23], Key_s2[23], Key_s1[23], Key_s0[23]}), .c ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, TweakeyGeneration_StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[24]}), .a ({Key_s3[24], Key_s2[24], Key_s1[24], Key_s0[24]}), .c ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, TweakeyGeneration_key_Feedback[25]}), .a ({Key_s3[25], Key_s2[25], Key_s1[25], Key_s0[25]}), .c ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, TweakeyGeneration_StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[26]}), .a ({Key_s3[26], Key_s2[26], Key_s1[26], Key_s0[26]}), .c ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, TweakeyGeneration_key_Feedback[27]}), .a ({Key_s3[27], Key_s2[27], Key_s1[27], Key_s0[27]}), .c ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, TweakeyGeneration_StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[28]}), .a ({Key_s3[28], Key_s2[28], Key_s1[28], Key_s0[28]}), .c ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, TweakeyGeneration_key_Feedback[29]}), .a ({Key_s3[29], Key_s2[29], Key_s1[29], Key_s0[29]}), .c ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, TweakeyGeneration_StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[30]}), .a ({Key_s3[30], Key_s2[30], Key_s1[30], Key_s0[30]}), .c ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, TweakeyGeneration_key_Feedback[31]}), .a ({Key_s3[31], Key_s2[31], Key_s1[31], Key_s0[31]}), .c ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, TweakeyGeneration_StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, TweakeyGeneration_key_Feedback[32]}), .a ({Key_s3[32], Key_s2[32], Key_s1[32], Key_s0[32]}), .c ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, TweakeyGeneration_StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, TweakeyGeneration_key_Feedback[33]}), .a ({Key_s3[33], Key_s2[33], Key_s1[33], Key_s0[33]}), .c ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, TweakeyGeneration_StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, TweakeyGeneration_key_Feedback[34]}), .a ({Key_s3[34], Key_s2[34], Key_s1[34], Key_s0[34]}), .c ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, TweakeyGeneration_StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, TweakeyGeneration_key_Feedback[35]}), .a ({Key_s3[35], Key_s2[35], Key_s1[35], Key_s0[35]}), .c ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, TweakeyGeneration_StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, TweakeyGeneration_key_Feedback[36]}), .a ({Key_s3[36], Key_s2[36], Key_s1[36], Key_s0[36]}), .c ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, TweakeyGeneration_StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, TweakeyGeneration_key_Feedback[37]}), .a ({Key_s3[37], Key_s2[37], Key_s1[37], Key_s0[37]}), .c ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, TweakeyGeneration_StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, TweakeyGeneration_key_Feedback[38]}), .a ({Key_s3[38], Key_s2[38], Key_s1[38], Key_s0[38]}), .c ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, TweakeyGeneration_StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, TweakeyGeneration_key_Feedback[39]}), .a ({Key_s3[39], Key_s2[39], Key_s1[39], Key_s0[39]}), .c ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, TweakeyGeneration_StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, TweakeyGeneration_key_Feedback[40]}), .a ({Key_s3[40], Key_s2[40], Key_s1[40], Key_s0[40]}), .c ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, TweakeyGeneration_StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, TweakeyGeneration_key_Feedback[41]}), .a ({Key_s3[41], Key_s2[41], Key_s1[41], Key_s0[41]}), .c ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, TweakeyGeneration_StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, TweakeyGeneration_key_Feedback[42]}), .a ({Key_s3[42], Key_s2[42], Key_s1[42], Key_s0[42]}), .c ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, TweakeyGeneration_StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, TweakeyGeneration_key_Feedback[43]}), .a ({Key_s3[43], Key_s2[43], Key_s1[43], Key_s0[43]}), .c ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, TweakeyGeneration_StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, TweakeyGeneration_key_Feedback[44]}), .a ({Key_s3[44], Key_s2[44], Key_s1[44], Key_s0[44]}), .c ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, TweakeyGeneration_StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, TweakeyGeneration_key_Feedback[45]}), .a ({Key_s3[45], Key_s2[45], Key_s1[45], Key_s0[45]}), .c ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, TweakeyGeneration_StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, TweakeyGeneration_key_Feedback[46]}), .a ({Key_s3[46], Key_s2[46], Key_s1[46], Key_s0[46]}), .c ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, TweakeyGeneration_StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, TweakeyGeneration_key_Feedback[47]}), .a ({Key_s3[47], Key_s2[47], Key_s1[47], Key_s0[47]}), .c ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, TweakeyGeneration_StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, TweakeyGeneration_key_Feedback[48]}), .a ({Key_s3[48], Key_s2[48], Key_s1[48], Key_s0[48]}), .c ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, TweakeyGeneration_StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, TweakeyGeneration_key_Feedback[49]}), .a ({Key_s3[49], Key_s2[49], Key_s1[49], Key_s0[49]}), .c ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, TweakeyGeneration_StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, TweakeyGeneration_key_Feedback[50]}), .a ({Key_s3[50], Key_s2[50], Key_s1[50], Key_s0[50]}), .c ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, TweakeyGeneration_StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, TweakeyGeneration_key_Feedback[51]}), .a ({Key_s3[51], Key_s2[51], Key_s1[51], Key_s0[51]}), .c ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, TweakeyGeneration_StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, TweakeyGeneration_key_Feedback[52]}), .a ({Key_s3[52], Key_s2[52], Key_s1[52], Key_s0[52]}), .c ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, TweakeyGeneration_StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, TweakeyGeneration_key_Feedback[53]}), .a ({Key_s3[53], Key_s2[53], Key_s1[53], Key_s0[53]}), .c ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, TweakeyGeneration_StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, TweakeyGeneration_key_Feedback[54]}), .a ({Key_s3[54], Key_s2[54], Key_s1[54], Key_s0[54]}), .c ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, TweakeyGeneration_StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, TweakeyGeneration_key_Feedback[55]}), .a ({Key_s3[55], Key_s2[55], Key_s1[55], Key_s0[55]}), .c ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, TweakeyGeneration_StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, TweakeyGeneration_key_Feedback[56]}), .a ({Key_s3[56], Key_s2[56], Key_s1[56], Key_s0[56]}), .c ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, TweakeyGeneration_StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, TweakeyGeneration_key_Feedback[57]}), .a ({Key_s3[57], Key_s2[57], Key_s1[57], Key_s0[57]}), .c ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, TweakeyGeneration_StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, TweakeyGeneration_key_Feedback[58]}), .a ({Key_s3[58], Key_s2[58], Key_s1[58], Key_s0[58]}), .c ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, TweakeyGeneration_StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, TweakeyGeneration_key_Feedback[59]}), .a ({Key_s3[59], Key_s2[59], Key_s1[59], Key_s0[59]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, TweakeyGeneration_StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, TweakeyGeneration_key_Feedback[60]}), .a ({Key_s3[60], Key_s2[60], Key_s1[60], Key_s0[60]}), .c ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, TweakeyGeneration_StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, TweakeyGeneration_key_Feedback[61]}), .a ({Key_s3[61], Key_s2[61], Key_s1[61], Key_s0[61]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, TweakeyGeneration_StateRegInput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, TweakeyGeneration_key_Feedback[62]}), .a ({Key_s3[62], Key_s2[62], Key_s1[62], Key_s0[62]}), .c ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, TweakeyGeneration_StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_KEYMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, TweakeyGeneration_key_Feedback[63]}), .a ({Key_s3[63], Key_s2[63], Key_s1[63], Key_s0[63]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, TweakeyGeneration_StateRegInput[63]}) ) ;
    MUX2_X1 FSMMUX_MUXInst_0_U1 ( .S (rst), .A (FSMUpdate[0]), .B (1'b1), .Z (FSMSelected[0]) ) ;
    MUX2_X1 FSMMUX_MUXInst_1_U1 ( .S (rst), .A (FSMUpdate[1]), .B (1'b0), .Z (FSMSelected[1]) ) ;
    MUX2_X1 FSMMUX_MUXInst_2_U1 ( .S (rst), .A (FSMUpdate[2]), .B (1'b0), .Z (FSMSelected[2]) ) ;
    MUX2_X1 FSMMUX_MUXInst_3_U1 ( .S (rst), .A (FSMUpdate[3]), .B (1'b0), .Z (FSMSelected[3]) ) ;
    MUX2_X1 FSMMUX_MUXInst_4_U1 ( .S (rst), .A (FSMUpdate[4]), .B (1'b0), .Z (FSMSelected[4]) ) ;
    MUX2_X1 FSMMUX_MUXInst_5_U1 ( .S (rst), .A (FSMUpdate[5]), .B (1'b0), .Z (FSMSelected[5]) ) ;
    MUX2_X1 FSMUpdateInst_StateUpdateInst_0_U5 ( .S (FSM[4]), .A (FSMUpdateInst_StateUpdateInst_0_n4), .B (FSM[5]), .Z (FSMUpdate[0]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U4 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_0_n3), .ZN (FSMUpdateInst_StateUpdateInst_0_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_0_U3 ( .A1 (FSMUpdateInst_StateUpdateInst_0_n2), .A2 (FSMUpdateInst_StateUpdateInst_0_n1), .ZN (FSMUpdateInst_StateUpdateInst_0_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_0_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_0_n1) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_0_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_0_n2) ) ;
    AND2_X1 FSMUpdateInst_StateUpdateInst_2_U5 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n4), .A2 (FSM[1]), .ZN (FSMUpdate[2]) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U4 ( .A1 (FSMUpdateInst_StateUpdateInst_2_n3), .A2 (FSM[5]), .ZN (FSMUpdateInst_StateUpdateInst_2_n4) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U3 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_2_n2), .ZN (FSMUpdateInst_StateUpdateInst_2_n3) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_2_U2 ( .A1 (FSMUpdate[1]), .A2 (FSMUpdateInst_StateUpdateInst_2_n1), .ZN (FSMUpdateInst_StateUpdateInst_2_n2) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_2_U1 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdate[4]), .ZN (FSMUpdateInst_StateUpdateInst_2_n1) ) ;
    OR2_X1 FSMUpdateInst_StateUpdateInst_5_U5 ( .A1 (FSM[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n4), .ZN (FSMUpdate[5]) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U4 ( .A1 (FSMUpdate[4]), .A2 (FSMUpdateInst_StateUpdateInst_5_n3), .ZN (FSMUpdateInst_StateUpdateInst_5_n4) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U3 ( .A1 (FSM[5]), .A2 (FSMUpdateInst_StateUpdateInst_5_n2), .ZN (FSMUpdateInst_StateUpdateInst_5_n3) ) ;
    NOR2_X1 FSMUpdateInst_StateUpdateInst_5_U2 ( .A1 (FSMUpdate[3]), .A2 (FSMUpdateInst_StateUpdateInst_5_n1), .ZN (FSMUpdateInst_StateUpdateInst_5_n2) ) ;
    NAND2_X1 FSMUpdateInst_StateUpdateInst_5_U1 ( .A1 (FSMUpdate[1]), .A2 (FSM[1]), .ZN (FSMUpdateInst_StateUpdateInst_5_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U6 ( .A1 (FSMSignalsInst_doneInst_n5), .A2 (FSMSignalsInst_doneInst_n4), .ZN (done) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U5 ( .A1 (FSM[4]), .A2 (FSM[5]), .ZN (FSMSignalsInst_doneInst_n4) ) ;
    NAND2_X1 FSMSignalsInst_doneInst_U4 ( .A1 (FSMSignalsInst_doneInst_n3), .A2 (FSMSignalsInst_doneInst_n2), .ZN (FSMSignalsInst_doneInst_n5) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U3 ( .A1 (FSMUpdate[4]), .A2 (FSMSignalsInst_doneInst_n1), .ZN (FSMSignalsInst_doneInst_n2) ) ;
    INV_X1 FSMSignalsInst_doneInst_U2 ( .A (FSMUpdate[1]), .ZN (FSMSignalsInst_doneInst_n1) ) ;
    NOR2_X1 FSMSignalsInst_doneInst_U1 ( .A1 (FSM[1]), .A2 (FSMUpdate[3]), .ZN (FSMSignalsInst_doneInst_n3) ) ;
    ClockGatingController #(3) ClockGatingInst ( .clk (clk), .rst (rst), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_2_U1 ( .s (rst), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, MCOutput[2]}), .a ({Plaintext_s3[2], Plaintext_s2[2], Plaintext_s1[2], Plaintext_s0[2]}), .c ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, StateRegInput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_3_U1 ( .s (rst), .b ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, MCOutput[3]}), .a ({Plaintext_s3[3], Plaintext_s2[3], Plaintext_s1[3], Plaintext_s0[3]}), .c ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, StateRegInput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_6_U1 ( .s (rst), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, MCOutput[6]}), .a ({Plaintext_s3[6], Plaintext_s2[6], Plaintext_s1[6], Plaintext_s0[6]}), .c ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, StateRegInput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_7_U1 ( .s (rst), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, MCOutput[7]}), .a ({Plaintext_s3[7], Plaintext_s2[7], Plaintext_s1[7], Plaintext_s0[7]}), .c ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, StateRegInput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_10_U1 ( .s (rst), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, MCOutput[10]}), .a ({Plaintext_s3[10], Plaintext_s2[10], Plaintext_s1[10], Plaintext_s0[10]}), .c ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, StateRegInput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_11_U1 ( .s (rst), .b ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, MCOutput[11]}), .a ({Plaintext_s3[11], Plaintext_s2[11], Plaintext_s1[11], Plaintext_s0[11]}), .c ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, StateRegInput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_14_U1 ( .s (rst), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, new_AGEMA_signal_3771, MCOutput[14]}), .a ({Plaintext_s3[14], Plaintext_s2[14], Plaintext_s1[14], Plaintext_s0[14]}), .c ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, new_AGEMA_signal_3798, StateRegInput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_15_U1 ( .s (rst), .b ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903, MCOutput[15]}), .a ({Plaintext_s3[15], Plaintext_s2[15], Plaintext_s1[15], Plaintext_s0[15]}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, new_AGEMA_signal_3927, StateRegInput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_18_U1 ( .s (rst), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, MCOutput[18]}), .a ({Plaintext_s3[18], Plaintext_s2[18], Plaintext_s1[18], Plaintext_s0[18]}), .c ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, StateRegInput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_19_U1 ( .s (rst), .b ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, MCOutput[19]}), .a ({Plaintext_s3[19], Plaintext_s2[19], Plaintext_s1[19], Plaintext_s0[19]}), .c ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, StateRegInput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_22_U1 ( .s (rst), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, MCOutput[22]}), .a ({Plaintext_s3[22], Plaintext_s2[22], Plaintext_s1[22], Plaintext_s0[22]}), .c ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, StateRegInput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_23_U1 ( .s (rst), .b ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, MCOutput[23]}), .a ({Plaintext_s3[23], Plaintext_s2[23], Plaintext_s1[23], Plaintext_s0[23]}), .c ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, StateRegInput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_26_U1 ( .s (rst), .b ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, new_AGEMA_signal_3741, MCOutput[26]}), .a ({Plaintext_s3[26], Plaintext_s2[26], Plaintext_s1[26], Plaintext_s0[26]}), .c ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, new_AGEMA_signal_3816, StateRegInput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_27_U1 ( .s (rst), .b ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, new_AGEMA_signal_3885, MCOutput[27]}), .a ({Plaintext_s3[27], Plaintext_s2[27], Plaintext_s1[27], Plaintext_s0[27]}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, new_AGEMA_signal_3945, StateRegInput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_30_U1 ( .s (rst), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, MCOutput[30]}), .a ({Plaintext_s3[30], Plaintext_s2[30], Plaintext_s1[30], Plaintext_s0[30]}), .c ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, StateRegInput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_31_U1 ( .s (rst), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, MCOutput[31]}), .a ({Plaintext_s3[31], Plaintext_s2[31], Plaintext_s1[31], Plaintext_s0[31]}), .c ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, StateRegInput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_34_U1 ( .s (rst), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}), .a ({Plaintext_s3[34], Plaintext_s2[34], Plaintext_s1[34], Plaintext_s0[34]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, StateRegInput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_35_U1 ( .s (rst), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}), .a ({Plaintext_s3[35], Plaintext_s2[35], Plaintext_s1[35], Plaintext_s0[35]}), .c ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, StateRegInput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_38_U1 ( .s (rst), .b ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}), .a ({Plaintext_s3[38], Plaintext_s2[38], Plaintext_s1[38], Plaintext_s0[38]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, StateRegInput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_39_U1 ( .s (rst), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}), .a ({Plaintext_s3[39], Plaintext_s2[39], Plaintext_s1[39], Plaintext_s0[39]}), .c ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, StateRegInput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_42_U1 ( .s (rst), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}), .a ({Plaintext_s3[42], Plaintext_s2[42], Plaintext_s1[42], Plaintext_s0[42]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, StateRegInput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_43_U1 ( .s (rst), .b ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}), .a ({Plaintext_s3[43], Plaintext_s2[43], Plaintext_s1[43], Plaintext_s0[43]}), .c ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, StateRegInput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_46_U1 ( .s (rst), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}), .a ({Plaintext_s3[46], Plaintext_s2[46], Plaintext_s1[46], Plaintext_s0[46]}), .c ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, StateRegInput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_47_U1 ( .s (rst), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}), .a ({Plaintext_s3[47], Plaintext_s2[47], Plaintext_s1[47], Plaintext_s0[47]}), .c ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, StateRegInput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_50_U1 ( .s (rst), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, MCOutput[50]}), .a ({Plaintext_s3[50], Plaintext_s2[50], Plaintext_s1[50], Plaintext_s0[50]}), .c ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, StateRegInput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_51_U1 ( .s (rst), .b ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, MCOutput[51]}), .a ({Plaintext_s3[51], Plaintext_s2[51], Plaintext_s1[51], Plaintext_s0[51]}), .c ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, StateRegInput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_54_U1 ( .s (rst), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, MCOutput[54]}), .a ({Plaintext_s3[54], Plaintext_s2[54], Plaintext_s1[54], Plaintext_s0[54]}), .c ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, StateRegInput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_55_U1 ( .s (rst), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, MCOutput[55]}), .a ({Plaintext_s3[55], Plaintext_s2[55], Plaintext_s1[55], Plaintext_s0[55]}), .c ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, StateRegInput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_58_U1 ( .s (rst), .b ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, MCOutput[58]}), .a ({Plaintext_s3[58], Plaintext_s2[58], Plaintext_s1[58], Plaintext_s0[58]}), .c ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, StateRegInput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_59_U1 ( .s (rst), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, MCOutput[59]}), .a ({Plaintext_s3[59], Plaintext_s2[59], Plaintext_s1[59], Plaintext_s0[59]}), .c ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, StateRegInput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_62_U1 ( .s (rst), .b ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, new_AGEMA_signal_3723, MCOutput[62]}), .a ({Plaintext_s3[62], Plaintext_s2[62], Plaintext_s1[62], Plaintext_s0[62]}), .c ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, new_AGEMA_signal_3852, StateRegInput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_63_U1 ( .s (rst), .b ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, new_AGEMA_signal_3873, MCOutput[63]}), .a ({Plaintext_s3[63], Plaintext_s2[63], Plaintext_s1[63], Plaintext_s0[63]}), .c ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, new_AGEMA_signal_3981, StateRegInput[63]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U3 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, ShiftRowsOutput[7]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_U2 ( .a ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, SubCellInst_SboxInst_0_YY_0_}), .b ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, ShiftRowsOutput[6]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_AND1_U1 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_2036, new_AGEMA_signal_2035, new_AGEMA_signal_2034, SubCellInst_SboxInst_0_Q1}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, SubCellInst_SboxInst_0_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR2_U1 ( .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, new_AGEMA_signal_2031, SubCellInst_SboxInst_0_Q0}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, SubCellInst_SboxInst_0_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_AND3_U1 ( .a ({new_AGEMA_signal_1169, new_AGEMA_signal_1168, new_AGEMA_signal_1167, SubCellInst_SboxInst_0_n3}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, new_AGEMA_signal_2037, SubCellInst_SboxInst_0_Q4}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR7_U1 ( .a ({new_AGEMA_signal_2324, new_AGEMA_signal_2323, new_AGEMA_signal_2322, SubCellInst_SboxInst_0_L1}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, SubCellInst_SboxInst_0_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR11_U1 ( .a ({new_AGEMA_signal_1181, new_AGEMA_signal_1180, new_AGEMA_signal_1179, SubCellInst_SboxInst_0_XX_2_}), .b ({new_AGEMA_signal_2318, new_AGEMA_signal_2317, new_AGEMA_signal_2316, SubCellInst_SboxInst_0_T0}), .c ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, SubCellInst_SboxInst_0_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR12_U1 ( .a ({new_AGEMA_signal_2468, new_AGEMA_signal_2467, new_AGEMA_signal_2466, SubCellInst_SboxInst_0_L3}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, SubCellInst_SboxInst_0_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR13_U1 ( .a ({new_AGEMA_signal_1175, new_AGEMA_signal_1174, new_AGEMA_signal_1173, SubCellInst_SboxInst_0_XX_1_}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, new_AGEMA_signal_2469, SubCellInst_SboxInst_0_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U3 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[11]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_U2 ( .a ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, SubCellInst_SboxInst_1_YY_0_}), .b ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, ShiftRowsOutput[10]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_AND1_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_2054, new_AGEMA_signal_2053, new_AGEMA_signal_2052, SubCellInst_SboxInst_1_Q1}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, SubCellInst_SboxInst_1_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR2_U1 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, new_AGEMA_signal_2049, SubCellInst_SboxInst_1_Q0}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, SubCellInst_SboxInst_1_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_AND3_U1 ( .a ({new_AGEMA_signal_1187, new_AGEMA_signal_1186, new_AGEMA_signal_1185, SubCellInst_SboxInst_1_n3}), .b ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, new_AGEMA_signal_2055, SubCellInst_SboxInst_1_Q4}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR7_U1 ( .a ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, new_AGEMA_signal_2331, SubCellInst_SboxInst_1_L1}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, SubCellInst_SboxInst_1_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR11_U1 ( .a ({new_AGEMA_signal_1199, new_AGEMA_signal_1198, new_AGEMA_signal_1197, SubCellInst_SboxInst_1_XX_2_}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, new_AGEMA_signal_2325, SubCellInst_SboxInst_1_T0}), .c ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, SubCellInst_SboxInst_1_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR12_U1 ( .a ({new_AGEMA_signal_2480, new_AGEMA_signal_2479, new_AGEMA_signal_2478, SubCellInst_SboxInst_1_L3}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, SubCellInst_SboxInst_1_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR13_U1 ( .a ({new_AGEMA_signal_1193, new_AGEMA_signal_1192, new_AGEMA_signal_1191, SubCellInst_SboxInst_1_XX_1_}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2483, new_AGEMA_signal_2482, new_AGEMA_signal_2481, SubCellInst_SboxInst_1_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U3 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, ShiftRowsOutput[15]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_U2 ( .a ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, SubCellInst_SboxInst_2_YY_0_}), .b ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, ShiftRowsOutput[14]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_AND1_U1 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_2072, new_AGEMA_signal_2071, new_AGEMA_signal_2070, SubCellInst_SboxInst_2_Q1}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_2_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR2_U1 ( .a ({new_AGEMA_signal_2069, new_AGEMA_signal_2068, new_AGEMA_signal_2067, SubCellInst_SboxInst_2_Q0}), .b ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, SubCellInst_SboxInst_2_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_AND3_U1 ( .a ({new_AGEMA_signal_1205, new_AGEMA_signal_1204, new_AGEMA_signal_1203, SubCellInst_SboxInst_2_n3}), .b ({new_AGEMA_signal_2075, new_AGEMA_signal_2074, new_AGEMA_signal_2073, SubCellInst_SboxInst_2_Q4}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR7_U1 ( .a ({new_AGEMA_signal_2342, new_AGEMA_signal_2341, new_AGEMA_signal_2340, SubCellInst_SboxInst_2_L1}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, SubCellInst_SboxInst_2_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR11_U1 ( .a ({new_AGEMA_signal_1217, new_AGEMA_signal_1216, new_AGEMA_signal_1215, SubCellInst_SboxInst_2_XX_2_}), .b ({new_AGEMA_signal_2336, new_AGEMA_signal_2335, new_AGEMA_signal_2334, SubCellInst_SboxInst_2_T0}), .c ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, SubCellInst_SboxInst_2_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR12_U1 ( .a ({new_AGEMA_signal_2492, new_AGEMA_signal_2491, new_AGEMA_signal_2490, SubCellInst_SboxInst_2_L3}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, SubCellInst_SboxInst_2_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR13_U1 ( .a ({new_AGEMA_signal_1211, new_AGEMA_signal_1210, new_AGEMA_signal_1209, SubCellInst_SboxInst_2_XX_1_}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2495, new_AGEMA_signal_2494, new_AGEMA_signal_2493, SubCellInst_SboxInst_2_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U3 ( .a ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, ShiftRowsOutput[3]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_U2 ( .a ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, SubCellInst_SboxInst_3_YY_0_}), .b ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, ShiftRowsOutput[2]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_AND1_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_2090, new_AGEMA_signal_2089, new_AGEMA_signal_2088, SubCellInst_SboxInst_3_Q1}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, SubCellInst_SboxInst_3_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR2_U1 ( .a ({new_AGEMA_signal_2087, new_AGEMA_signal_2086, new_AGEMA_signal_2085, SubCellInst_SboxInst_3_Q0}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, SubCellInst_SboxInst_3_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_AND3_U1 ( .a ({new_AGEMA_signal_1223, new_AGEMA_signal_1222, new_AGEMA_signal_1221, SubCellInst_SboxInst_3_n3}), .b ({new_AGEMA_signal_2093, new_AGEMA_signal_2092, new_AGEMA_signal_2091, SubCellInst_SboxInst_3_Q4}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR7_U1 ( .a ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, new_AGEMA_signal_2349, SubCellInst_SboxInst_3_L1}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, SubCellInst_SboxInst_3_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR11_U1 ( .a ({new_AGEMA_signal_1235, new_AGEMA_signal_1234, new_AGEMA_signal_1233, SubCellInst_SboxInst_3_XX_2_}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, new_AGEMA_signal_2343, SubCellInst_SboxInst_3_T0}), .c ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellInst_SboxInst_3_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR12_U1 ( .a ({new_AGEMA_signal_2504, new_AGEMA_signal_2503, new_AGEMA_signal_2502, SubCellInst_SboxInst_3_L3}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, SubCellInst_SboxInst_3_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR13_U1 ( .a ({new_AGEMA_signal_1229, new_AGEMA_signal_1228, new_AGEMA_signal_1227, SubCellInst_SboxInst_3_XX_1_}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2507, new_AGEMA_signal_2506, new_AGEMA_signal_2505, SubCellInst_SboxInst_3_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U3 ( .a ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_U2 ( .a ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, SubCellInst_SboxInst_4_YY_0_}), .b ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_AND1_U1 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_2108, new_AGEMA_signal_2107, new_AGEMA_signal_2106, SubCellInst_SboxInst_4_Q1}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, SubCellInst_SboxInst_4_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR2_U1 ( .a ({new_AGEMA_signal_2105, new_AGEMA_signal_2104, new_AGEMA_signal_2103, SubCellInst_SboxInst_4_Q0}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, SubCellInst_SboxInst_4_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_AND3_U1 ( .a ({new_AGEMA_signal_1241, new_AGEMA_signal_1240, new_AGEMA_signal_1239, SubCellInst_SboxInst_4_n3}), .b ({new_AGEMA_signal_2111, new_AGEMA_signal_2110, new_AGEMA_signal_2109, SubCellInst_SboxInst_4_Q4}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR7_U1 ( .a ({new_AGEMA_signal_2360, new_AGEMA_signal_2359, new_AGEMA_signal_2358, SubCellInst_SboxInst_4_L1}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, SubCellInst_SboxInst_4_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR11_U1 ( .a ({new_AGEMA_signal_1253, new_AGEMA_signal_1252, new_AGEMA_signal_1251, SubCellInst_SboxInst_4_XX_2_}), .b ({new_AGEMA_signal_2354, new_AGEMA_signal_2353, new_AGEMA_signal_2352, SubCellInst_SboxInst_4_T0}), .c ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, SubCellInst_SboxInst_4_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR12_U1 ( .a ({new_AGEMA_signal_2516, new_AGEMA_signal_2515, new_AGEMA_signal_2514, SubCellInst_SboxInst_4_L3}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, SubCellInst_SboxInst_4_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR13_U1 ( .a ({new_AGEMA_signal_1247, new_AGEMA_signal_1246, new_AGEMA_signal_1245, SubCellInst_SboxInst_4_XX_1_}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2519, new_AGEMA_signal_2518, new_AGEMA_signal_2517, SubCellInst_SboxInst_4_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U3 ( .a ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_U2 ( .a ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, SubCellInst_SboxInst_5_YY_0_}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_AND1_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_2126, new_AGEMA_signal_2125, new_AGEMA_signal_2124, SubCellInst_SboxInst_5_Q1}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, SubCellInst_SboxInst_5_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR2_U1 ( .a ({new_AGEMA_signal_2123, new_AGEMA_signal_2122, new_AGEMA_signal_2121, SubCellInst_SboxInst_5_Q0}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, SubCellInst_SboxInst_5_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_AND3_U1 ( .a ({new_AGEMA_signal_1259, new_AGEMA_signal_1258, new_AGEMA_signal_1257, SubCellInst_SboxInst_5_n3}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, new_AGEMA_signal_2127, SubCellInst_SboxInst_5_Q4}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR7_U1 ( .a ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, new_AGEMA_signal_2367, SubCellInst_SboxInst_5_L1}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, SubCellInst_SboxInst_5_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR11_U1 ( .a ({new_AGEMA_signal_1271, new_AGEMA_signal_1270, new_AGEMA_signal_1269, SubCellInst_SboxInst_5_XX_2_}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, new_AGEMA_signal_2361, SubCellInst_SboxInst_5_T0}), .c ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, SubCellInst_SboxInst_5_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR12_U1 ( .a ({new_AGEMA_signal_2528, new_AGEMA_signal_2527, new_AGEMA_signal_2526, SubCellInst_SboxInst_5_L3}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, SubCellInst_SboxInst_5_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR13_U1 ( .a ({new_AGEMA_signal_1265, new_AGEMA_signal_1264, new_AGEMA_signal_1263, SubCellInst_SboxInst_5_XX_1_}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2531, new_AGEMA_signal_2530, new_AGEMA_signal_2529, SubCellInst_SboxInst_5_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U3 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_U2 ( .a ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, SubCellInst_SboxInst_6_YY_0_}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_AND1_U1 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_2144, new_AGEMA_signal_2143, new_AGEMA_signal_2142, SubCellInst_SboxInst_6_Q1}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, SubCellInst_SboxInst_6_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR2_U1 ( .a ({new_AGEMA_signal_2141, new_AGEMA_signal_2140, new_AGEMA_signal_2139, SubCellInst_SboxInst_6_Q0}), .b ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, SubCellInst_SboxInst_6_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_AND3_U1 ( .a ({new_AGEMA_signal_1277, new_AGEMA_signal_1276, new_AGEMA_signal_1275, SubCellInst_SboxInst_6_n3}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, new_AGEMA_signal_2145, SubCellInst_SboxInst_6_Q4}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR7_U1 ( .a ({new_AGEMA_signal_2378, new_AGEMA_signal_2377, new_AGEMA_signal_2376, SubCellInst_SboxInst_6_L1}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, SubCellInst_SboxInst_6_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR11_U1 ( .a ({new_AGEMA_signal_1289, new_AGEMA_signal_1288, new_AGEMA_signal_1287, SubCellInst_SboxInst_6_XX_2_}), .b ({new_AGEMA_signal_2372, new_AGEMA_signal_2371, new_AGEMA_signal_2370, SubCellInst_SboxInst_6_T0}), .c ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, SubCellInst_SboxInst_6_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR12_U1 ( .a ({new_AGEMA_signal_2540, new_AGEMA_signal_2539, new_AGEMA_signal_2538, SubCellInst_SboxInst_6_L3}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, SubCellInst_SboxInst_6_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR13_U1 ( .a ({new_AGEMA_signal_1283, new_AGEMA_signal_1282, new_AGEMA_signal_1281, SubCellInst_SboxInst_6_XX_1_}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2543, new_AGEMA_signal_2542, new_AGEMA_signal_2541, SubCellInst_SboxInst_6_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U3 ( .a ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_U2 ( .a ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, SubCellInst_SboxInst_7_YY_0_}), .b ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_AND1_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_2162, new_AGEMA_signal_2161, new_AGEMA_signal_2160, SubCellInst_SboxInst_7_Q1}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, SubCellInst_SboxInst_7_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR2_U1 ( .a ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, new_AGEMA_signal_2157, SubCellInst_SboxInst_7_Q0}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, SubCellInst_SboxInst_7_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_AND3_U1 ( .a ({new_AGEMA_signal_1295, new_AGEMA_signal_1294, new_AGEMA_signal_1293, SubCellInst_SboxInst_7_n3}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, new_AGEMA_signal_2163, SubCellInst_SboxInst_7_Q4}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR7_U1 ( .a ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, new_AGEMA_signal_2385, SubCellInst_SboxInst_7_L1}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, SubCellInst_SboxInst_7_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR11_U1 ( .a ({new_AGEMA_signal_1307, new_AGEMA_signal_1306, new_AGEMA_signal_1305, SubCellInst_SboxInst_7_XX_2_}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, new_AGEMA_signal_2379, SubCellInst_SboxInst_7_T0}), .c ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, SubCellInst_SboxInst_7_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR12_U1 ( .a ({new_AGEMA_signal_2552, new_AGEMA_signal_2551, new_AGEMA_signal_2550, SubCellInst_SboxInst_7_L3}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, SubCellInst_SboxInst_7_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR13_U1 ( .a ({new_AGEMA_signal_1301, new_AGEMA_signal_1300, new_AGEMA_signal_1299, SubCellInst_SboxInst_7_XX_1_}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2555, new_AGEMA_signal_2554, new_AGEMA_signal_2553, SubCellInst_SboxInst_7_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U3 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, AddRoundConstantOutput[35]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_U2 ( .a ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, SubCellInst_SboxInst_8_YY_0_}), .b ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, AddRoundConstantOutput[34]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_AND1_U1 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_2180, new_AGEMA_signal_2179, new_AGEMA_signal_2178, SubCellInst_SboxInst_8_Q1}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_8_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR2_U1 ( .a ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, new_AGEMA_signal_2175, SubCellInst_SboxInst_8_Q0}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, SubCellInst_SboxInst_8_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_AND3_U1 ( .a ({new_AGEMA_signal_1313, new_AGEMA_signal_1312, new_AGEMA_signal_1311, SubCellInst_SboxInst_8_n3}), .b ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, new_AGEMA_signal_2181, SubCellInst_SboxInst_8_Q4}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR7_U1 ( .a ({new_AGEMA_signal_2396, new_AGEMA_signal_2395, new_AGEMA_signal_2394, SubCellInst_SboxInst_8_L1}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, SubCellInst_SboxInst_8_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR11_U1 ( .a ({new_AGEMA_signal_1325, new_AGEMA_signal_1324, new_AGEMA_signal_1323, SubCellInst_SboxInst_8_XX_2_}), .b ({new_AGEMA_signal_2390, new_AGEMA_signal_2389, new_AGEMA_signal_2388, SubCellInst_SboxInst_8_T0}), .c ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, SubCellInst_SboxInst_8_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR12_U1 ( .a ({new_AGEMA_signal_2564, new_AGEMA_signal_2563, new_AGEMA_signal_2562, SubCellInst_SboxInst_8_L3}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, SubCellInst_SboxInst_8_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR13_U1 ( .a ({new_AGEMA_signal_1319, new_AGEMA_signal_1318, new_AGEMA_signal_1317, SubCellInst_SboxInst_8_XX_1_}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2567, new_AGEMA_signal_2566, new_AGEMA_signal_2565, SubCellInst_SboxInst_8_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U3 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, AddRoundConstantOutput[39]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_U2 ( .a ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, SubCellInst_SboxInst_9_YY_0_}), .b ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, AddRoundConstantOutput[38]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_AND1_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_2198, new_AGEMA_signal_2197, new_AGEMA_signal_2196, SubCellInst_SboxInst_9_Q1}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, SubCellInst_SboxInst_9_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR2_U1 ( .a ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, new_AGEMA_signal_2193, SubCellInst_SboxInst_9_Q0}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, SubCellInst_SboxInst_9_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_AND3_U1 ( .a ({new_AGEMA_signal_1331, new_AGEMA_signal_1330, new_AGEMA_signal_1329, SubCellInst_SboxInst_9_n3}), .b ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, new_AGEMA_signal_2199, SubCellInst_SboxInst_9_Q4}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR7_U1 ( .a ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, new_AGEMA_signal_2403, SubCellInst_SboxInst_9_L1}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, SubCellInst_SboxInst_9_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR11_U1 ( .a ({new_AGEMA_signal_1343, new_AGEMA_signal_1342, new_AGEMA_signal_1341, SubCellInst_SboxInst_9_XX_2_}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, new_AGEMA_signal_2397, SubCellInst_SboxInst_9_T0}), .c ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, SubCellInst_SboxInst_9_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR12_U1 ( .a ({new_AGEMA_signal_2576, new_AGEMA_signal_2575, new_AGEMA_signal_2574, SubCellInst_SboxInst_9_L3}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, SubCellInst_SboxInst_9_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR13_U1 ( .a ({new_AGEMA_signal_1337, new_AGEMA_signal_1336, new_AGEMA_signal_1335, SubCellInst_SboxInst_9_XX_1_}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, new_AGEMA_signal_2577, SubCellInst_SboxInst_9_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U3 ( .a ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, AddRoundConstantOutput[43]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_U2 ( .a ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, SubCellInst_SboxInst_10_YY_0_}), .b ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, AddRoundConstantOutput[42]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_AND1_U1 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_2216, new_AGEMA_signal_2215, new_AGEMA_signal_2214, SubCellInst_SboxInst_10_Q1}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, SubCellInst_SboxInst_10_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR2_U1 ( .a ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, new_AGEMA_signal_2211, SubCellInst_SboxInst_10_Q0}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, SubCellInst_SboxInst_10_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_AND3_U1 ( .a ({new_AGEMA_signal_1349, new_AGEMA_signal_1348, new_AGEMA_signal_1347, SubCellInst_SboxInst_10_n3}), .b ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, new_AGEMA_signal_2217, SubCellInst_SboxInst_10_Q4}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR7_U1 ( .a ({new_AGEMA_signal_2414, new_AGEMA_signal_2413, new_AGEMA_signal_2412, SubCellInst_SboxInst_10_L1}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, SubCellInst_SboxInst_10_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR11_U1 ( .a ({new_AGEMA_signal_1361, new_AGEMA_signal_1360, new_AGEMA_signal_1359, SubCellInst_SboxInst_10_XX_2_}), .b ({new_AGEMA_signal_2408, new_AGEMA_signal_2407, new_AGEMA_signal_2406, SubCellInst_SboxInst_10_T0}), .c ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, SubCellInst_SboxInst_10_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR12_U1 ( .a ({new_AGEMA_signal_2588, new_AGEMA_signal_2587, new_AGEMA_signal_2586, SubCellInst_SboxInst_10_L3}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, SubCellInst_SboxInst_10_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR13_U1 ( .a ({new_AGEMA_signal_1355, new_AGEMA_signal_1354, new_AGEMA_signal_1353, SubCellInst_SboxInst_10_XX_1_}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, new_AGEMA_signal_2589, SubCellInst_SboxInst_10_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U3 ( .a ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, SubCellOutput[47]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_U2 ( .a ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, SubCellInst_SboxInst_11_YY_0_}), .b ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, SubCellOutput[46]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_AND1_U1 ( .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_2234, new_AGEMA_signal_2233, new_AGEMA_signal_2232, SubCellInst_SboxInst_11_Q1}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, SubCellInst_SboxInst_11_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR2_U1 ( .a ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, new_AGEMA_signal_2229, SubCellInst_SboxInst_11_Q0}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, SubCellInst_SboxInst_11_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_AND3_U1 ( .a ({new_AGEMA_signal_1367, new_AGEMA_signal_1366, new_AGEMA_signal_1365, SubCellInst_SboxInst_11_n3}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, new_AGEMA_signal_2235, SubCellInst_SboxInst_11_Q4}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR7_U1 ( .a ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, new_AGEMA_signal_2421, SubCellInst_SboxInst_11_L1}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, SubCellInst_SboxInst_11_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR11_U1 ( .a ({new_AGEMA_signal_1379, new_AGEMA_signal_1378, new_AGEMA_signal_1377, SubCellInst_SboxInst_11_XX_2_}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, new_AGEMA_signal_2415, SubCellInst_SboxInst_11_T0}), .c ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, SubCellInst_SboxInst_11_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR12_U1 ( .a ({new_AGEMA_signal_2600, new_AGEMA_signal_2599, new_AGEMA_signal_2598, SubCellInst_SboxInst_11_L3}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, SubCellInst_SboxInst_11_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR13_U1 ( .a ({new_AGEMA_signal_1373, new_AGEMA_signal_1372, new_AGEMA_signal_1371, SubCellInst_SboxInst_11_XX_1_}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, new_AGEMA_signal_2601, SubCellInst_SboxInst_11_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U3 ( .a ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, AddRoundConstantOutput[51]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_U2 ( .a ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, SubCellInst_SboxInst_12_YY_0_}), .b ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, AddRoundConstantOutput[50]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_AND1_U1 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_2252, new_AGEMA_signal_2251, new_AGEMA_signal_2250, SubCellInst_SboxInst_12_Q1}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_12_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR2_U1 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, new_AGEMA_signal_2247, SubCellInst_SboxInst_12_Q0}), .b ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, SubCellInst_SboxInst_12_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_AND3_U1 ( .a ({new_AGEMA_signal_1385, new_AGEMA_signal_1384, new_AGEMA_signal_1383, SubCellInst_SboxInst_12_n3}), .b ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, new_AGEMA_signal_2253, SubCellInst_SboxInst_12_Q4}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR7_U1 ( .a ({new_AGEMA_signal_2432, new_AGEMA_signal_2431, new_AGEMA_signal_2430, SubCellInst_SboxInst_12_L1}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, SubCellInst_SboxInst_12_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR11_U1 ( .a ({new_AGEMA_signal_1397, new_AGEMA_signal_1396, new_AGEMA_signal_1395, SubCellInst_SboxInst_12_XX_2_}), .b ({new_AGEMA_signal_2426, new_AGEMA_signal_2425, new_AGEMA_signal_2424, SubCellInst_SboxInst_12_T0}), .c ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, SubCellInst_SboxInst_12_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR12_U1 ( .a ({new_AGEMA_signal_2612, new_AGEMA_signal_2611, new_AGEMA_signal_2610, SubCellInst_SboxInst_12_L3}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, SubCellInst_SboxInst_12_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR13_U1 ( .a ({new_AGEMA_signal_1391, new_AGEMA_signal_1390, new_AGEMA_signal_1389, SubCellInst_SboxInst_12_XX_1_}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, new_AGEMA_signal_2613, SubCellInst_SboxInst_12_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U3 ( .a ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, AddRoundConstantOutput[55]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_U2 ( .a ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, SubCellInst_SboxInst_13_YY_0_}), .b ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, AddRoundConstantOutput[54]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_AND1_U1 ( .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_2270, new_AGEMA_signal_2269, new_AGEMA_signal_2268, SubCellInst_SboxInst_13_Q1}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, SubCellInst_SboxInst_13_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR2_U1 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, new_AGEMA_signal_2265, SubCellInst_SboxInst_13_Q0}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, SubCellInst_SboxInst_13_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_AND3_U1 ( .a ({new_AGEMA_signal_1403, new_AGEMA_signal_1402, new_AGEMA_signal_1401, SubCellInst_SboxInst_13_n3}), .b ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, new_AGEMA_signal_2271, SubCellInst_SboxInst_13_Q4}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR7_U1 ( .a ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, new_AGEMA_signal_2439, SubCellInst_SboxInst_13_L1}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, SubCellInst_SboxInst_13_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR11_U1 ( .a ({new_AGEMA_signal_1415, new_AGEMA_signal_1414, new_AGEMA_signal_1413, SubCellInst_SboxInst_13_XX_2_}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, new_AGEMA_signal_2433, SubCellInst_SboxInst_13_T0}), .c ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, SubCellInst_SboxInst_13_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR12_U1 ( .a ({new_AGEMA_signal_2624, new_AGEMA_signal_2623, new_AGEMA_signal_2622, SubCellInst_SboxInst_13_L3}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, SubCellInst_SboxInst_13_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR13_U1 ( .a ({new_AGEMA_signal_1409, new_AGEMA_signal_1408, new_AGEMA_signal_1407, SubCellInst_SboxInst_13_XX_1_}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, new_AGEMA_signal_2625, SubCellInst_SboxInst_13_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U3 ( .a ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, AddRoundConstantOutput[59]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_U2 ( .a ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, SubCellInst_SboxInst_14_YY_0_}), .b ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, AddRoundConstantOutput[58]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_AND1_U1 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_2288, new_AGEMA_signal_2287, new_AGEMA_signal_2286, SubCellInst_SboxInst_14_Q1}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, SubCellInst_SboxInst_14_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR2_U1 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, new_AGEMA_signal_2283, SubCellInst_SboxInst_14_Q0}), .b ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, SubCellInst_SboxInst_14_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_AND3_U1 ( .a ({new_AGEMA_signal_1421, new_AGEMA_signal_1420, new_AGEMA_signal_1419, SubCellInst_SboxInst_14_n3}), .b ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, new_AGEMA_signal_2289, SubCellInst_SboxInst_14_Q4}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR7_U1 ( .a ({new_AGEMA_signal_2450, new_AGEMA_signal_2449, new_AGEMA_signal_2448, SubCellInst_SboxInst_14_L1}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, SubCellInst_SboxInst_14_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR11_U1 ( .a ({new_AGEMA_signal_1433, new_AGEMA_signal_1432, new_AGEMA_signal_1431, SubCellInst_SboxInst_14_XX_2_}), .b ({new_AGEMA_signal_2444, new_AGEMA_signal_2443, new_AGEMA_signal_2442, SubCellInst_SboxInst_14_T0}), .c ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, SubCellInst_SboxInst_14_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR12_U1 ( .a ({new_AGEMA_signal_2636, new_AGEMA_signal_2635, new_AGEMA_signal_2634, SubCellInst_SboxInst_14_L3}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, SubCellInst_SboxInst_14_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR13_U1 ( .a ({new_AGEMA_signal_1427, new_AGEMA_signal_1426, new_AGEMA_signal_1425, SubCellInst_SboxInst_14_XX_1_}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, new_AGEMA_signal_2637, SubCellInst_SboxInst_14_YY_0_}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U3 ( .a ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, SubCellOutput[63]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_U2 ( .a ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, SubCellInst_SboxInst_15_YY_0_}), .b ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, SubCellOutput[62]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_AND1_U1 ( .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_2306, new_AGEMA_signal_2305, new_AGEMA_signal_2304, SubCellInst_SboxInst_15_Q1}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, SubCellInst_SboxInst_15_T0}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR2_U1 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, new_AGEMA_signal_2301, SubCellInst_SboxInst_15_Q0}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, SubCellInst_SboxInst_15_Q2}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_AND3_U1 ( .a ({new_AGEMA_signal_1439, new_AGEMA_signal_1438, new_AGEMA_signal_1437, SubCellInst_SboxInst_15_n3}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, new_AGEMA_signal_2307, SubCellInst_SboxInst_15_Q4}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR7_U1 ( .a ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, new_AGEMA_signal_2457, SubCellInst_SboxInst_15_L1}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, SubCellInst_SboxInst_15_Q7}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR11_U1 ( .a ({new_AGEMA_signal_1451, new_AGEMA_signal_1450, new_AGEMA_signal_1449, SubCellInst_SboxInst_15_XX_2_}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, new_AGEMA_signal_2451, SubCellInst_SboxInst_15_T0}), .c ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, SubCellInst_SboxInst_15_L3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR12_U1 ( .a ({new_AGEMA_signal_2648, new_AGEMA_signal_2647, new_AGEMA_signal_2646, SubCellInst_SboxInst_15_L3}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, SubCellInst_SboxInst_15_YY_1_}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR13_U1 ( .a ({new_AGEMA_signal_1445, new_AGEMA_signal_1444, new_AGEMA_signal_1443, SubCellInst_SboxInst_15_XX_1_}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, new_AGEMA_signal_2649, SubCellInst_SboxInst_15_YY_0_}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, AddConstXOR_AddConstXOR_XORInst_0_2_n1}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[3]}), .c ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, AddRoundConstantOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2834, new_AGEMA_signal_2833, new_AGEMA_signal_2832, SubCellOutput[62]}), .c ({new_AGEMA_signal_2942, new_AGEMA_signal_2941, new_AGEMA_signal_2940, AddConstXOR_AddConstXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, AddConstXOR_AddConstXOR_XORInst_0_3_n1}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[4]}), .c ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, AddRoundConstantOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2936, new_AGEMA_signal_2935, new_AGEMA_signal_2934, SubCellOutput[63]}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, new_AGEMA_signal_3075, AddConstXOR_AddConstXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, AddConstXOR_AddConstXOR_XORInst_1_2_n1}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, AddRoundConstantOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2786, new_AGEMA_signal_2785, new_AGEMA_signal_2784, SubCellOutput[46]}), .c ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, new_AGEMA_signal_2943, AddConstXOR_AddConstXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, AddConstXOR_AddConstXOR_XORInst_1_3_n1}), .b ({1'b0, 1'b0, 1'b0, 1'b0}), .c ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, AddRoundConstantOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2912, new_AGEMA_signal_2911, new_AGEMA_signal_2910, SubCellOutput[47]}), .c ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, new_AGEMA_signal_3081, AddConstXOR_AddConstXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, AddRoundTweakeyXOR_XORInst_0_2_n1}), .b ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[2]}), .c ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, ShiftRowsOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2750, new_AGEMA_signal_2749, new_AGEMA_signal_2748, AddRoundConstantOutput[34]}), .c ({new_AGEMA_signal_2948, new_AGEMA_signal_2947, new_AGEMA_signal_2946, AddRoundTweakeyXOR_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, AddRoundTweakeyXOR_XORInst_0_3_n1}), .b ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, TweakeyGeneration_key_Feedback[3]}), .c ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, ShiftRowsOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2894, new_AGEMA_signal_2893, new_AGEMA_signal_2892, AddRoundConstantOutput[35]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, new_AGEMA_signal_3087, AddRoundTweakeyXOR_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, AddRoundTweakeyXOR_XORInst_1_2_n1}), .b ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[6]}), .c ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, ShiftRowsOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2762, new_AGEMA_signal_2761, new_AGEMA_signal_2760, AddRoundConstantOutput[38]}), .c ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, new_AGEMA_signal_2949, AddRoundTweakeyXOR_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, AddRoundTweakeyXOR_XORInst_1_3_n1}), .b ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, TweakeyGeneration_key_Feedback[7]}), .c ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, ShiftRowsOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2900, new_AGEMA_signal_2899, new_AGEMA_signal_2898, AddRoundConstantOutput[39]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, new_AGEMA_signal_3093, AddRoundTweakeyXOR_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, AddRoundTweakeyXOR_XORInst_2_2_n1}), .b ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[10]}), .c ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, ShiftRowsOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2774, new_AGEMA_signal_2773, new_AGEMA_signal_2772, AddRoundConstantOutput[42]}), .c ({new_AGEMA_signal_2954, new_AGEMA_signal_2953, new_AGEMA_signal_2952, AddRoundTweakeyXOR_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, AddRoundTweakeyXOR_XORInst_2_3_n1}), .b ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, TweakeyGeneration_key_Feedback[11]}), .c ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, ShiftRowsOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2906, new_AGEMA_signal_2905, new_AGEMA_signal_2904, AddRoundConstantOutput[43]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, new_AGEMA_signal_3099, AddRoundTweakeyXOR_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, AddRoundTweakeyXOR_XORInst_3_2_n1}), .b ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[14]}), .c ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, ShiftRowsOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3080, new_AGEMA_signal_3079, new_AGEMA_signal_3078, AddRoundConstantOutput[46]}), .c ({new_AGEMA_signal_3230, new_AGEMA_signal_3229, new_AGEMA_signal_3228, AddRoundTweakeyXOR_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, AddRoundTweakeyXOR_XORInst_3_3_n1}), .b ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, TweakeyGeneration_key_Feedback[15]}), .c ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, ShiftRowsOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, new_AGEMA_signal_3207, AddRoundConstantOutput[47]}), .c ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, new_AGEMA_signal_3345, AddRoundTweakeyXOR_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_2_U2 ( .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, AddRoundTweakeyXOR_XORInst_4_2_n1}), .b ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[18]}), .c ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2798, new_AGEMA_signal_2797, new_AGEMA_signal_2796, AddRoundConstantOutput[50]}), .c ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, new_AGEMA_signal_2955, AddRoundTweakeyXOR_XORInst_4_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_3_U2 ( .a ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, AddRoundTweakeyXOR_XORInst_4_3_n1}), .b ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, TweakeyGeneration_key_Feedback[19]}), .c ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2918, new_AGEMA_signal_2917, new_AGEMA_signal_2916, AddRoundConstantOutput[51]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, new_AGEMA_signal_3105, AddRoundTweakeyXOR_XORInst_4_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_2_U2 ( .a ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, AddRoundTweakeyXOR_XORInst_5_2_n1}), .b ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[22]}), .c ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2810, new_AGEMA_signal_2809, new_AGEMA_signal_2808, AddRoundConstantOutput[54]}), .c ({new_AGEMA_signal_2960, new_AGEMA_signal_2959, new_AGEMA_signal_2958, AddRoundTweakeyXOR_XORInst_5_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_3_U2 ( .a ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, AddRoundTweakeyXOR_XORInst_5_3_n1}), .b ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, TweakeyGeneration_key_Feedback[23]}), .c ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2924, new_AGEMA_signal_2923, new_AGEMA_signal_2922, AddRoundConstantOutput[55]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, new_AGEMA_signal_3111, AddRoundTweakeyXOR_XORInst_5_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_2_U2 ( .a ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, AddRoundTweakeyXOR_XORInst_6_2_n1}), .b ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[26]}), .c ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2822, new_AGEMA_signal_2821, new_AGEMA_signal_2820, AddRoundConstantOutput[58]}), .c ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, new_AGEMA_signal_2961, AddRoundTweakeyXOR_XORInst_6_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_3_U2 ( .a ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, AddRoundTweakeyXOR_XORInst_6_3_n1}), .b ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, TweakeyGeneration_key_Feedback[27]}), .c ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_2930, new_AGEMA_signal_2929, new_AGEMA_signal_2928, AddRoundConstantOutput[59]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, new_AGEMA_signal_3117, AddRoundTweakeyXOR_XORInst_6_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_2_U2 ( .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, AddRoundTweakeyXOR_XORInst_7_2_n1}), .b ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[30]}), .c ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3074, new_AGEMA_signal_3073, new_AGEMA_signal_3072, AddRoundConstantOutput[62]}), .c ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, new_AGEMA_signal_3249, AddRoundTweakeyXOR_XORInst_7_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_3_U2 ( .a ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, AddRoundTweakeyXOR_XORInst_7_3_n1}), .b ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, TweakeyGeneration_key_Feedback[31]}), .c ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, new_AGEMA_signal_3201, AddRoundConstantOutput[63]}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, new_AGEMA_signal_3369, AddRoundTweakeyXOR_XORInst_7_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U3 ( .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, MCInst_MCR0_XORInst_0_2_n2}), .b ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCInst_MCR0_XORInst_0_2_n1}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, new_AGEMA_signal_3375, MCOutput[50]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}), .b ({new_AGEMA_signal_2690, new_AGEMA_signal_2689, new_AGEMA_signal_2688, ShiftRowsOutput[2]}), .c ({new_AGEMA_signal_2966, new_AGEMA_signal_2965, new_AGEMA_signal_2964, MCInst_MCR0_XORInst_0_2_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}), .c ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, new_AGEMA_signal_3255, MCInst_MCR0_XORInst_0_2_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U3 ( .a ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, MCInst_MCR0_XORInst_0_3_n2}), .b ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, MCInst_MCR0_XORInst_0_3_n1}), .c ({new_AGEMA_signal_3554, new_AGEMA_signal_3553, new_AGEMA_signal_3552, MCOutput[51]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}), .b ({new_AGEMA_signal_2864, new_AGEMA_signal_2863, new_AGEMA_signal_2862, ShiftRowsOutput[3]}), .c ({new_AGEMA_signal_3122, new_AGEMA_signal_3121, new_AGEMA_signal_3120, MCInst_MCR0_XORInst_0_3_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}), .c ({new_AGEMA_signal_3380, new_AGEMA_signal_3379, new_AGEMA_signal_3378, MCInst_MCR0_XORInst_0_3_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U3 ( .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, MCInst_MCR0_XORInst_1_2_n2}), .b ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, MCInst_MCR0_XORInst_1_2_n1}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, new_AGEMA_signal_3381, MCOutput[54]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}), .b ({new_AGEMA_signal_2654, new_AGEMA_signal_2653, new_AGEMA_signal_2652, ShiftRowsOutput[6]}), .c ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, new_AGEMA_signal_2967, MCInst_MCR0_XORInst_1_2_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}), .c ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, new_AGEMA_signal_3261, MCInst_MCR0_XORInst_1_2_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U3 ( .a ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, MCInst_MCR0_XORInst_1_3_n2}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, MCInst_MCR0_XORInst_1_3_n1}), .c ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, new_AGEMA_signal_3561, MCOutput[55]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}), .b ({new_AGEMA_signal_2846, new_AGEMA_signal_2845, new_AGEMA_signal_2844, ShiftRowsOutput[7]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, new_AGEMA_signal_3123, MCInst_MCR0_XORInst_1_3_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}), .c ({new_AGEMA_signal_3386, new_AGEMA_signal_3385, new_AGEMA_signal_3384, MCInst_MCR0_XORInst_1_3_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U3 ( .a ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, MCInst_MCR0_XORInst_2_2_n2}), .b ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCInst_MCR0_XORInst_2_2_n1}), .c ({new_AGEMA_signal_3392, new_AGEMA_signal_3391, new_AGEMA_signal_3390, MCOutput[58]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}), .b ({new_AGEMA_signal_2666, new_AGEMA_signal_2665, new_AGEMA_signal_2664, ShiftRowsOutput[10]}), .c ({new_AGEMA_signal_2972, new_AGEMA_signal_2971, new_AGEMA_signal_2970, MCInst_MCR0_XORInst_2_2_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}), .c ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, new_AGEMA_signal_3267, MCInst_MCR0_XORInst_2_2_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U3 ( .a ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, MCInst_MCR0_XORInst_2_3_n2}), .b ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, MCInst_MCR0_XORInst_2_3_n1}), .c ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, new_AGEMA_signal_3567, MCOutput[59]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}), .b ({new_AGEMA_signal_2852, new_AGEMA_signal_2851, new_AGEMA_signal_2850, ShiftRowsOutput[11]}), .c ({new_AGEMA_signal_3128, new_AGEMA_signal_3127, new_AGEMA_signal_3126, MCInst_MCR0_XORInst_2_3_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, new_AGEMA_signal_3393, MCInst_MCR0_XORInst_2_3_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U3 ( .a ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, MCInst_MCR0_XORInst_3_2_n2}), .b ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, MCInst_MCR0_XORInst_3_2_n1}), .c ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, new_AGEMA_signal_3723, MCOutput[62]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}), .b ({new_AGEMA_signal_2678, new_AGEMA_signal_2677, new_AGEMA_signal_2676, ShiftRowsOutput[14]}), .c ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, new_AGEMA_signal_2973, MCInst_MCR0_XORInst_3_2_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}), .c ({new_AGEMA_signal_3572, new_AGEMA_signal_3571, new_AGEMA_signal_3570, MCInst_MCR0_XORInst_3_2_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U3 ( .a ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726, MCInst_MCR0_XORInst_3_3_n2}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, MCInst_MCR0_XORInst_3_3_n1}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, new_AGEMA_signal_3873, MCOutput[63]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}), .b ({new_AGEMA_signal_2858, new_AGEMA_signal_2857, new_AGEMA_signal_2856, ShiftRowsOutput[15]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, new_AGEMA_signal_3129, MCInst_MCR0_XORInst_3_3_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}), .c ({new_AGEMA_signal_3728, new_AGEMA_signal_3727, new_AGEMA_signal_3726, MCInst_MCR0_XORInst_3_3_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, MCInst_MCR2_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, new_AGEMA_signal_3399, MCOutput[18]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3092, new_AGEMA_signal_3091, new_AGEMA_signal_3090, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, new_AGEMA_signal_3273, MCInst_MCR2_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, MCInst_MCR2_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_3578, new_AGEMA_signal_3577, new_AGEMA_signal_3576, MCOutput[19]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, new_AGEMA_signal_3219, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_3404, new_AGEMA_signal_3403, new_AGEMA_signal_3402, MCInst_MCR2_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, MCInst_MCR2_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, new_AGEMA_signal_3405, MCOutput[22]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3098, new_AGEMA_signal_3097, new_AGEMA_signal_3096, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_3278, new_AGEMA_signal_3277, new_AGEMA_signal_3276, MCInst_MCR2_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, MCInst_MCR2_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_3584, new_AGEMA_signal_3583, new_AGEMA_signal_3582, MCOutput[23]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, new_AGEMA_signal_3225, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_3410, new_AGEMA_signal_3409, new_AGEMA_signal_3408, MCInst_MCR2_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, MCInst_MCR2_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, new_AGEMA_signal_3741, MCOutput[26]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3344, new_AGEMA_signal_3343, new_AGEMA_signal_3342, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, new_AGEMA_signal_3585, MCInst_MCR2_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, new_AGEMA_signal_3744, MCInst_MCR2_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, new_AGEMA_signal_3885, MCOutput[27]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, new_AGEMA_signal_3531, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_3746, new_AGEMA_signal_3745, new_AGEMA_signal_3744, MCInst_MCR2_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, MCInst_MCR2_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, new_AGEMA_signal_3411, MCOutput[30]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3086, new_AGEMA_signal_3085, new_AGEMA_signal_3084, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, new_AGEMA_signal_3279, MCInst_MCR2_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, MCInst_MCR2_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, new_AGEMA_signal_3591, MCOutput[31]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, new_AGEMA_signal_3213, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_3416, new_AGEMA_signal_3415, new_AGEMA_signal_3414, MCInst_MCR2_XORInst_3_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_2_U2 ( .a ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, MCInst_MCR3_XORInst_0_2_n1}), .b ({new_AGEMA_signal_2726, new_AGEMA_signal_2725, new_AGEMA_signal_2724, ShiftRowsOutput[18]}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, new_AGEMA_signal_3417, MCOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3104, new_AGEMA_signal_3103, new_AGEMA_signal_3102, MCOutput[34]}), .c ({new_AGEMA_signal_3284, new_AGEMA_signal_3283, new_AGEMA_signal_3282, MCInst_MCR3_XORInst_0_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_3_U2 ( .a ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, MCInst_MCR3_XORInst_0_3_n1}), .b ({new_AGEMA_signal_2882, new_AGEMA_signal_2881, new_AGEMA_signal_2880, ShiftRowsOutput[19]}), .c ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, new_AGEMA_signal_3597, MCOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3236, new_AGEMA_signal_3235, new_AGEMA_signal_3234, MCOutput[35]}), .c ({new_AGEMA_signal_3422, new_AGEMA_signal_3421, new_AGEMA_signal_3420, MCInst_MCR3_XORInst_0_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_2_U2 ( .a ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, MCInst_MCR3_XORInst_1_2_n1}), .b ({new_AGEMA_signal_2738, new_AGEMA_signal_2737, new_AGEMA_signal_2736, ShiftRowsOutput[22]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, new_AGEMA_signal_3423, MCOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3110, new_AGEMA_signal_3109, new_AGEMA_signal_3108, MCOutput[38]}), .c ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, new_AGEMA_signal_3285, MCInst_MCR3_XORInst_1_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_3_U2 ( .a ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, MCInst_MCR3_XORInst_1_3_n1}), .b ({new_AGEMA_signal_2888, new_AGEMA_signal_2887, new_AGEMA_signal_2886, ShiftRowsOutput[23]}), .c ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, new_AGEMA_signal_3603, MCOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3242, new_AGEMA_signal_3241, new_AGEMA_signal_3240, MCOutput[39]}), .c ({new_AGEMA_signal_3428, new_AGEMA_signal_3427, new_AGEMA_signal_3426, MCInst_MCR3_XORInst_1_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_2_U2 ( .a ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, MCInst_MCR3_XORInst_2_2_n1}), .b ({new_AGEMA_signal_2702, new_AGEMA_signal_2701, new_AGEMA_signal_2700, ShiftRowsOutput[26]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, new_AGEMA_signal_3429, MCOutput[10]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3116, new_AGEMA_signal_3115, new_AGEMA_signal_3114, MCOutput[42]}), .c ({new_AGEMA_signal_3290, new_AGEMA_signal_3289, new_AGEMA_signal_3288, MCInst_MCR3_XORInst_2_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_3_U2 ( .a ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, MCInst_MCR3_XORInst_2_3_n1}), .b ({new_AGEMA_signal_2870, new_AGEMA_signal_2869, new_AGEMA_signal_2868, ShiftRowsOutput[27]}), .c ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, new_AGEMA_signal_3609, MCOutput[11]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3248, new_AGEMA_signal_3247, new_AGEMA_signal_3246, MCOutput[43]}), .c ({new_AGEMA_signal_3434, new_AGEMA_signal_3433, new_AGEMA_signal_3432, MCInst_MCR3_XORInst_2_3_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_2_U2 ( .a ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, MCInst_MCR3_XORInst_3_2_n1}), .b ({new_AGEMA_signal_2714, new_AGEMA_signal_2713, new_AGEMA_signal_2712, ShiftRowsOutput[30]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, new_AGEMA_signal_3771, MCOutput[14]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_2_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3368, new_AGEMA_signal_3367, new_AGEMA_signal_3366, MCOutput[46]}), .c ({new_AGEMA_signal_3614, new_AGEMA_signal_3613, new_AGEMA_signal_3612, MCInst_MCR3_XORInst_3_2_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_3_U2 ( .a ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, new_AGEMA_signal_3774, MCInst_MCR3_XORInst_3_3_n1}), .b ({new_AGEMA_signal_2876, new_AGEMA_signal_2875, new_AGEMA_signal_2874, ShiftRowsOutput[31]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, new_AGEMA_signal_3903, MCOutput[15]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_3_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3548, new_AGEMA_signal_3547, new_AGEMA_signal_3546, MCOutput[47]}), .c ({new_AGEMA_signal_3776, new_AGEMA_signal_3775, new_AGEMA_signal_3774, MCInst_MCR3_XORInst_3_3_n1}) ) ;

    /* cells in depth 2 */
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_0_U1 ( .s (rst), .b ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, new_AGEMA_signal_3753, MCOutput[0]}), .a ({Plaintext_s3[0], Plaintext_s2[0], Plaintext_s1[0], Plaintext_s0[0]}), .c ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, new_AGEMA_signal_3780, StateRegInput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_1_U1 ( .s (rst), .b ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891, MCOutput[1]}), .a ({Plaintext_s3[1], Plaintext_s2[1], Plaintext_s1[1], Plaintext_s0[1]}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, new_AGEMA_signal_3909, StateRegInput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_4_U1 ( .s (rst), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, new_AGEMA_signal_3759, MCOutput[4]}), .a ({Plaintext_s3[4], Plaintext_s2[4], Plaintext_s1[4], Plaintext_s0[4]}), .c ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, new_AGEMA_signal_3786, StateRegInput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_5_U1 ( .s (rst), .b ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, new_AGEMA_signal_3894, MCOutput[5]}), .a ({Plaintext_s3[5], Plaintext_s2[5], Plaintext_s1[5], Plaintext_s0[5]}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, new_AGEMA_signal_3915, StateRegInput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_8_U1 ( .s (rst), .b ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, new_AGEMA_signal_3765, MCOutput[8]}), .a ({Plaintext_s3[8], Plaintext_s2[8], Plaintext_s1[8], Plaintext_s0[8]}), .c ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, new_AGEMA_signal_3792, StateRegInput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_9_U1 ( .s (rst), .b ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, new_AGEMA_signal_3897, MCOutput[9]}), .a ({Plaintext_s3[9], Plaintext_s2[9], Plaintext_s1[9], Plaintext_s0[9]}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, new_AGEMA_signal_3921, StateRegInput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_12_U1 ( .s (rst), .b ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, new_AGEMA_signal_3996, MCOutput[12]}), .a ({Plaintext_s3[12], Plaintext_s2[12], Plaintext_s1[12], Plaintext_s0[12]}), .c ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, new_AGEMA_signal_4005, StateRegInput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_13_U1 ( .s (rst), .b ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026, MCOutput[13]}), .a ({Plaintext_s3[13], Plaintext_s2[13], Plaintext_s1[13], Plaintext_s0[13]}), .c ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, new_AGEMA_signal_4032, StateRegInput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_16_U1 ( .s (rst), .b ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, new_AGEMA_signal_3729, MCOutput[16]}), .a ({Plaintext_s3[16], Plaintext_s2[16], Plaintext_s1[16], Plaintext_s0[16]}), .c ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, new_AGEMA_signal_3804, StateRegInput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_17_U1 ( .s (rst), .b ({new_AGEMA_signal_3878, new_AGEMA_signal_3877, new_AGEMA_signal_3876, MCOutput[17]}), .a ({Plaintext_s3[17], Plaintext_s2[17], Plaintext_s1[17], Plaintext_s0[17]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, new_AGEMA_signal_3933, StateRegInput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_20_U1 ( .s (rst), .b ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735, MCOutput[20]}), .a ({Plaintext_s3[20], Plaintext_s2[20], Plaintext_s1[20], Plaintext_s0[20]}), .c ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, new_AGEMA_signal_3810, StateRegInput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_21_U1 ( .s (rst), .b ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, new_AGEMA_signal_3879, MCOutput[21]}), .a ({Plaintext_s3[21], Plaintext_s2[21], Plaintext_s1[21], Plaintext_s0[21]}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939, StateRegInput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_24_U1 ( .s (rst), .b ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, new_AGEMA_signal_3990, MCOutput[24]}), .a ({Plaintext_s3[24], Plaintext_s2[24], Plaintext_s1[24], Plaintext_s0[24]}), .c ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, new_AGEMA_signal_4011, StateRegInput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_25_U1 ( .s (rst), .b ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023, MCOutput[25]}), .a ({Plaintext_s3[25], Plaintext_s2[25], Plaintext_s1[25], Plaintext_s0[25]}), .c ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038, StateRegInput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_28_U1 ( .s (rst), .b ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747, MCOutput[28]}), .a ({Plaintext_s3[28], Plaintext_s2[28], Plaintext_s1[28], Plaintext_s0[28]}), .c ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822, StateRegInput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_29_U1 ( .s (rst), .b ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, new_AGEMA_signal_3888, MCOutput[29]}), .a ({Plaintext_s3[29], Plaintext_s2[29], Plaintext_s1[29], Plaintext_s0[29]}), .c ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, new_AGEMA_signal_3951, StateRegInput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_32_U1 ( .s (rst), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}), .a ({Plaintext_s3[32], Plaintext_s2[32], Plaintext_s1[32], Plaintext_s0[32]}), .c ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, StateRegInput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_33_U1 ( .s (rst), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}), .a ({Plaintext_s3[33], Plaintext_s2[33], Plaintext_s1[33], Plaintext_s0[33]}), .c ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, StateRegInput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_36_U1 ( .s (rst), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}), .a ({Plaintext_s3[36], Plaintext_s2[36], Plaintext_s1[36], Plaintext_s0[36]}), .c ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, StateRegInput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_37_U1 ( .s (rst), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}), .a ({Plaintext_s3[37], Plaintext_s2[37], Plaintext_s1[37], Plaintext_s0[37]}), .c ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, StateRegInput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_40_U1 ( .s (rst), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}), .a ({Plaintext_s3[40], Plaintext_s2[40], Plaintext_s1[40], Plaintext_s0[40]}), .c ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, StateRegInput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_41_U1 ( .s (rst), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}), .a ({Plaintext_s3[41], Plaintext_s2[41], Plaintext_s1[41], Plaintext_s0[41]}), .c ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, StateRegInput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_44_U1 ( .s (rst), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}), .a ({Plaintext_s3[44], Plaintext_s2[44], Plaintext_s1[44], Plaintext_s0[44]}), .c ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, new_AGEMA_signal_3828, StateRegInput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_45_U1 ( .s (rst), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}), .a ({Plaintext_s3[45], Plaintext_s2[45], Plaintext_s1[45], Plaintext_s0[45]}), .c ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, new_AGEMA_signal_3957, StateRegInput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_48_U1 ( .s (rst), .b ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, MCOutput[48]}), .a ({Plaintext_s3[48], Plaintext_s2[48], Plaintext_s1[48], Plaintext_s0[48]}), .c ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, new_AGEMA_signal_3834, StateRegInput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_49_U1 ( .s (rst), .b ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, new_AGEMA_signal_3861, MCOutput[49]}), .a ({Plaintext_s3[49], Plaintext_s2[49], Plaintext_s1[49], Plaintext_s0[49]}), .c ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, new_AGEMA_signal_3963, StateRegInput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_52_U1 ( .s (rst), .b ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, MCOutput[52]}), .a ({Plaintext_s3[52], Plaintext_s2[52], Plaintext_s1[52], Plaintext_s0[52]}), .c ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, new_AGEMA_signal_3840, StateRegInput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_53_U1 ( .s (rst), .b ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, new_AGEMA_signal_3864, MCOutput[53]}), .a ({Plaintext_s3[53], Plaintext_s2[53], Plaintext_s1[53], Plaintext_s0[53]}), .c ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, new_AGEMA_signal_3969, StateRegInput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_56_U1 ( .s (rst), .b ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, MCOutput[56]}), .a ({Plaintext_s3[56], Plaintext_s2[56], Plaintext_s1[56], Plaintext_s0[56]}), .c ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, new_AGEMA_signal_3846, StateRegInput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_57_U1 ( .s (rst), .b ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, new_AGEMA_signal_3867, MCOutput[57]}), .a ({Plaintext_s3[57], Plaintext_s2[57], Plaintext_s1[57], Plaintext_s0[57]}), .c ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975, StateRegInput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_60_U1 ( .s (rst), .b ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, new_AGEMA_signal_3984, MCOutput[60]}), .a ({Plaintext_s3[60], Plaintext_s2[60], Plaintext_s1[60], Plaintext_s0[60]}), .c ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, new_AGEMA_signal_4017, StateRegInput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) PlaintextMUX_MUXInst_61_U1 ( .s (rst), .b ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, new_AGEMA_signal_4020, MCOutput[61]}), .a ({Plaintext_s3[61], Plaintext_s2[61], Plaintext_s1[61], Plaintext_s0[61]}), .c ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, new_AGEMA_signal_4044, StateRegInput[61]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_AND2_U1 ( .a ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}), .b ({new_AGEMA_signal_2462, new_AGEMA_signal_2461, new_AGEMA_signal_2460, SubCellInst_SboxInst_0_Q2}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, SubCellInst_SboxInst_0_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR4_U1 ( .a ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, new_AGEMA_signal_2655, SubCellInst_SboxInst_0_T1}), .b ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, new_AGEMA_signal_2319, SubCellInst_SboxInst_0_T2}), .c ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, SubCellInst_SboxInst_0_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_AND4_U1 ( .a ({new_AGEMA_signal_2042, new_AGEMA_signal_2041, new_AGEMA_signal_2040, SubCellInst_SboxInst_0_Q6}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, new_AGEMA_signal_2463, SubCellInst_SboxInst_0_Q7}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, SubCellInst_SboxInst_0_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR9_U1 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, new_AGEMA_signal_2043, SubCellInst_SboxInst_0_L2}), .c ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, SubCellInst_SboxInst_0_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR10_U1 ( .a ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, new_AGEMA_signal_2847, SubCellInst_SboxInst_0_L0}), .b ({new_AGEMA_signal_2660, new_AGEMA_signal_2659, new_AGEMA_signal_2658, SubCellInst_SboxInst_0_T3}), .c ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, ShiftRowsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_0_XOR_o1_U1 ( .a ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, new_AGEMA_signal_2661, SubCellInst_SboxInst_0_YY_1_}), .b ({new_AGEMA_signal_2978, new_AGEMA_signal_2977, new_AGEMA_signal_2976, SubCellInst_SboxInst_0_YY_3}), .c ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, ShiftRowsOutput[5]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_AND2_U1 ( .a ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}), .b ({new_AGEMA_signal_2474, new_AGEMA_signal_2473, new_AGEMA_signal_2472, SubCellInst_SboxInst_1_Q2}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, SubCellInst_SboxInst_1_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR4_U1 ( .a ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, new_AGEMA_signal_2667, SubCellInst_SboxInst_1_T1}), .b ({new_AGEMA_signal_2330, new_AGEMA_signal_2329, new_AGEMA_signal_2328, SubCellInst_SboxInst_1_T2}), .c ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, SubCellInst_SboxInst_1_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_AND4_U1 ( .a ({new_AGEMA_signal_2060, new_AGEMA_signal_2059, new_AGEMA_signal_2058, SubCellInst_SboxInst_1_Q6}), .b ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, new_AGEMA_signal_2475, SubCellInst_SboxInst_1_Q7}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, SubCellInst_SboxInst_1_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR9_U1 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, new_AGEMA_signal_2061, SubCellInst_SboxInst_1_L2}), .c ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, SubCellInst_SboxInst_1_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR10_U1 ( .a ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, new_AGEMA_signal_2853, SubCellInst_SboxInst_1_L0}), .b ({new_AGEMA_signal_2672, new_AGEMA_signal_2671, new_AGEMA_signal_2670, SubCellInst_SboxInst_1_T3}), .c ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, ShiftRowsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_1_XOR_o1_U1 ( .a ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, new_AGEMA_signal_2673, SubCellInst_SboxInst_1_YY_1_}), .b ({new_AGEMA_signal_2984, new_AGEMA_signal_2983, new_AGEMA_signal_2982, SubCellInst_SboxInst_1_YY_3}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, ShiftRowsOutput[9]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_AND2_U1 ( .a ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}), .b ({new_AGEMA_signal_2486, new_AGEMA_signal_2485, new_AGEMA_signal_2484, SubCellInst_SboxInst_2_Q2}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, SubCellInst_SboxInst_2_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR4_U1 ( .a ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, new_AGEMA_signal_2679, SubCellInst_SboxInst_2_T1}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, new_AGEMA_signal_2337, SubCellInst_SboxInst_2_T2}), .c ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, SubCellInst_SboxInst_2_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_AND4_U1 ( .a ({new_AGEMA_signal_2078, new_AGEMA_signal_2077, new_AGEMA_signal_2076, SubCellInst_SboxInst_2_Q6}), .b ({new_AGEMA_signal_2489, new_AGEMA_signal_2488, new_AGEMA_signal_2487, SubCellInst_SboxInst_2_Q7}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, SubCellInst_SboxInst_2_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR9_U1 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_2081, new_AGEMA_signal_2080, new_AGEMA_signal_2079, SubCellInst_SboxInst_2_L2}), .c ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, SubCellInst_SboxInst_2_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR10_U1 ( .a ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, new_AGEMA_signal_2859, SubCellInst_SboxInst_2_L0}), .b ({new_AGEMA_signal_2684, new_AGEMA_signal_2683, new_AGEMA_signal_2682, SubCellInst_SboxInst_2_T3}), .c ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, ShiftRowsOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_2_XOR_o1_U1 ( .a ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, new_AGEMA_signal_2685, SubCellInst_SboxInst_2_YY_1_}), .b ({new_AGEMA_signal_2990, new_AGEMA_signal_2989, new_AGEMA_signal_2988, SubCellInst_SboxInst_2_YY_3}), .c ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, ShiftRowsOutput[13]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_AND2_U1 ( .a ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}), .b ({new_AGEMA_signal_2498, new_AGEMA_signal_2497, new_AGEMA_signal_2496, SubCellInst_SboxInst_3_Q2}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, SubCellInst_SboxInst_3_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR4_U1 ( .a ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, new_AGEMA_signal_2691, SubCellInst_SboxInst_3_T1}), .b ({new_AGEMA_signal_2348, new_AGEMA_signal_2347, new_AGEMA_signal_2346, SubCellInst_SboxInst_3_T2}), .c ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, SubCellInst_SboxInst_3_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_AND4_U1 ( .a ({new_AGEMA_signal_2096, new_AGEMA_signal_2095, new_AGEMA_signal_2094, SubCellInst_SboxInst_3_Q6}), .b ({new_AGEMA_signal_2501, new_AGEMA_signal_2500, new_AGEMA_signal_2499, SubCellInst_SboxInst_3_Q7}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, SubCellInst_SboxInst_3_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR9_U1 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_2099, new_AGEMA_signal_2098, new_AGEMA_signal_2097, SubCellInst_SboxInst_3_L2}), .c ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, SubCellInst_SboxInst_3_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR10_U1 ( .a ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, new_AGEMA_signal_2865, SubCellInst_SboxInst_3_L0}), .b ({new_AGEMA_signal_2696, new_AGEMA_signal_2695, new_AGEMA_signal_2694, SubCellInst_SboxInst_3_T3}), .c ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, ShiftRowsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_3_XOR_o1_U1 ( .a ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, new_AGEMA_signal_2697, SubCellInst_SboxInst_3_YY_1_}), .b ({new_AGEMA_signal_2996, new_AGEMA_signal_2995, new_AGEMA_signal_2994, SubCellInst_SboxInst_3_YY_3}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, ShiftRowsOutput[1]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_AND2_U1 ( .a ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}), .b ({new_AGEMA_signal_2510, new_AGEMA_signal_2509, new_AGEMA_signal_2508, SubCellInst_SboxInst_4_Q2}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, SubCellInst_SboxInst_4_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR4_U1 ( .a ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, new_AGEMA_signal_2703, SubCellInst_SboxInst_4_T1}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, new_AGEMA_signal_2355, SubCellInst_SboxInst_4_T2}), .c ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, SubCellInst_SboxInst_4_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_AND4_U1 ( .a ({new_AGEMA_signal_2114, new_AGEMA_signal_2113, new_AGEMA_signal_2112, SubCellInst_SboxInst_4_Q6}), .b ({new_AGEMA_signal_2513, new_AGEMA_signal_2512, new_AGEMA_signal_2511, SubCellInst_SboxInst_4_Q7}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, SubCellInst_SboxInst_4_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR9_U1 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, new_AGEMA_signal_2115, SubCellInst_SboxInst_4_L2}), .c ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, SubCellInst_SboxInst_4_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR10_U1 ( .a ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, new_AGEMA_signal_2871, SubCellInst_SboxInst_4_L0}), .b ({new_AGEMA_signal_2708, new_AGEMA_signal_2707, new_AGEMA_signal_2706, SubCellInst_SboxInst_4_T3}), .c ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_4_XOR_o1_U1 ( .a ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, new_AGEMA_signal_2709, SubCellInst_SboxInst_4_YY_1_}), .b ({new_AGEMA_signal_3002, new_AGEMA_signal_3001, new_AGEMA_signal_3000, SubCellInst_SboxInst_4_YY_3}), .c ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_AND2_U1 ( .a ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}), .b ({new_AGEMA_signal_2522, new_AGEMA_signal_2521, new_AGEMA_signal_2520, SubCellInst_SboxInst_5_Q2}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, SubCellInst_SboxInst_5_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR4_U1 ( .a ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, new_AGEMA_signal_2715, SubCellInst_SboxInst_5_T1}), .b ({new_AGEMA_signal_2366, new_AGEMA_signal_2365, new_AGEMA_signal_2364, SubCellInst_SboxInst_5_T2}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, SubCellInst_SboxInst_5_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_AND4_U1 ( .a ({new_AGEMA_signal_2132, new_AGEMA_signal_2131, new_AGEMA_signal_2130, SubCellInst_SboxInst_5_Q6}), .b ({new_AGEMA_signal_2525, new_AGEMA_signal_2524, new_AGEMA_signal_2523, SubCellInst_SboxInst_5_Q7}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, SubCellInst_SboxInst_5_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR9_U1 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_2135, new_AGEMA_signal_2134, new_AGEMA_signal_2133, SubCellInst_SboxInst_5_L2}), .c ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, SubCellInst_SboxInst_5_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR10_U1 ( .a ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, new_AGEMA_signal_2877, SubCellInst_SboxInst_5_L0}), .b ({new_AGEMA_signal_2720, new_AGEMA_signal_2719, new_AGEMA_signal_2718, SubCellInst_SboxInst_5_T3}), .c ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_5_XOR_o1_U1 ( .a ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, new_AGEMA_signal_2721, SubCellInst_SboxInst_5_YY_1_}), .b ({new_AGEMA_signal_3008, new_AGEMA_signal_3007, new_AGEMA_signal_3006, SubCellInst_SboxInst_5_YY_3}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_AND2_U1 ( .a ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}), .b ({new_AGEMA_signal_2534, new_AGEMA_signal_2533, new_AGEMA_signal_2532, SubCellInst_SboxInst_6_Q2}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, SubCellInst_SboxInst_6_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR4_U1 ( .a ({new_AGEMA_signal_2729, new_AGEMA_signal_2728, new_AGEMA_signal_2727, SubCellInst_SboxInst_6_T1}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, new_AGEMA_signal_2373, SubCellInst_SboxInst_6_T2}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, SubCellInst_SboxInst_6_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_AND4_U1 ( .a ({new_AGEMA_signal_2150, new_AGEMA_signal_2149, new_AGEMA_signal_2148, SubCellInst_SboxInst_6_Q6}), .b ({new_AGEMA_signal_2537, new_AGEMA_signal_2536, new_AGEMA_signal_2535, SubCellInst_SboxInst_6_Q7}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, SubCellInst_SboxInst_6_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR9_U1 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, new_AGEMA_signal_2151, SubCellInst_SboxInst_6_L2}), .c ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, SubCellInst_SboxInst_6_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR10_U1 ( .a ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, new_AGEMA_signal_2883, SubCellInst_SboxInst_6_L0}), .b ({new_AGEMA_signal_2732, new_AGEMA_signal_2731, new_AGEMA_signal_2730, SubCellInst_SboxInst_6_T3}), .c ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_6_XOR_o1_U1 ( .a ({new_AGEMA_signal_2735, new_AGEMA_signal_2734, new_AGEMA_signal_2733, SubCellInst_SboxInst_6_YY_1_}), .b ({new_AGEMA_signal_3014, new_AGEMA_signal_3013, new_AGEMA_signal_3012, SubCellInst_SboxInst_6_YY_3}), .c ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_AND2_U1 ( .a ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}), .b ({new_AGEMA_signal_2546, new_AGEMA_signal_2545, new_AGEMA_signal_2544, SubCellInst_SboxInst_7_Q2}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, SubCellInst_SboxInst_7_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR4_U1 ( .a ({new_AGEMA_signal_2741, new_AGEMA_signal_2740, new_AGEMA_signal_2739, SubCellInst_SboxInst_7_T1}), .b ({new_AGEMA_signal_2384, new_AGEMA_signal_2383, new_AGEMA_signal_2382, SubCellInst_SboxInst_7_T2}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, SubCellInst_SboxInst_7_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_AND4_U1 ( .a ({new_AGEMA_signal_2168, new_AGEMA_signal_2167, new_AGEMA_signal_2166, SubCellInst_SboxInst_7_Q6}), .b ({new_AGEMA_signal_2549, new_AGEMA_signal_2548, new_AGEMA_signal_2547, SubCellInst_SboxInst_7_Q7}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, SubCellInst_SboxInst_7_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR9_U1 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, new_AGEMA_signal_2169, SubCellInst_SboxInst_7_L2}), .c ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, SubCellInst_SboxInst_7_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR10_U1 ( .a ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, new_AGEMA_signal_2889, SubCellInst_SboxInst_7_L0}), .b ({new_AGEMA_signal_2744, new_AGEMA_signal_2743, new_AGEMA_signal_2742, SubCellInst_SboxInst_7_T3}), .c ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_7_XOR_o1_U1 ( .a ({new_AGEMA_signal_2747, new_AGEMA_signal_2746, new_AGEMA_signal_2745, SubCellInst_SboxInst_7_YY_1_}), .b ({new_AGEMA_signal_3020, new_AGEMA_signal_3019, new_AGEMA_signal_3018, SubCellInst_SboxInst_7_YY_3}), .c ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, SubCellOutput[29]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_AND2_U1 ( .a ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}), .b ({new_AGEMA_signal_2558, new_AGEMA_signal_2557, new_AGEMA_signal_2556, SubCellInst_SboxInst_8_Q2}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, SubCellInst_SboxInst_8_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR4_U1 ( .a ({new_AGEMA_signal_2753, new_AGEMA_signal_2752, new_AGEMA_signal_2751, SubCellInst_SboxInst_8_T1}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, new_AGEMA_signal_2391, SubCellInst_SboxInst_8_T2}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, SubCellInst_SboxInst_8_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_AND4_U1 ( .a ({new_AGEMA_signal_2186, new_AGEMA_signal_2185, new_AGEMA_signal_2184, SubCellInst_SboxInst_8_Q6}), .b ({new_AGEMA_signal_2561, new_AGEMA_signal_2560, new_AGEMA_signal_2559, SubCellInst_SboxInst_8_Q7}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, SubCellInst_SboxInst_8_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR9_U1 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, new_AGEMA_signal_2187, SubCellInst_SboxInst_8_L2}), .c ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, SubCellInst_SboxInst_8_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR10_U1 ( .a ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, new_AGEMA_signal_2895, SubCellInst_SboxInst_8_L0}), .b ({new_AGEMA_signal_2756, new_AGEMA_signal_2755, new_AGEMA_signal_2754, SubCellInst_SboxInst_8_T3}), .c ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, AddRoundConstantOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_8_XOR_o1_U1 ( .a ({new_AGEMA_signal_2759, new_AGEMA_signal_2758, new_AGEMA_signal_2757, SubCellInst_SboxInst_8_YY_1_}), .b ({new_AGEMA_signal_3026, new_AGEMA_signal_3025, new_AGEMA_signal_3024, SubCellInst_SboxInst_8_YY_3}), .c ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, AddRoundConstantOutput[33]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_AND2_U1 ( .a ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}), .b ({new_AGEMA_signal_2570, new_AGEMA_signal_2569, new_AGEMA_signal_2568, SubCellInst_SboxInst_9_Q2}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, SubCellInst_SboxInst_9_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR4_U1 ( .a ({new_AGEMA_signal_2765, new_AGEMA_signal_2764, new_AGEMA_signal_2763, SubCellInst_SboxInst_9_T1}), .b ({new_AGEMA_signal_2402, new_AGEMA_signal_2401, new_AGEMA_signal_2400, SubCellInst_SboxInst_9_T2}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, SubCellInst_SboxInst_9_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_AND4_U1 ( .a ({new_AGEMA_signal_2204, new_AGEMA_signal_2203, new_AGEMA_signal_2202, SubCellInst_SboxInst_9_Q6}), .b ({new_AGEMA_signal_2573, new_AGEMA_signal_2572, new_AGEMA_signal_2571, SubCellInst_SboxInst_9_Q7}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, SubCellInst_SboxInst_9_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR9_U1 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, new_AGEMA_signal_2205, SubCellInst_SboxInst_9_L2}), .c ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, SubCellInst_SboxInst_9_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR10_U1 ( .a ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, new_AGEMA_signal_2901, SubCellInst_SboxInst_9_L0}), .b ({new_AGEMA_signal_2768, new_AGEMA_signal_2767, new_AGEMA_signal_2766, SubCellInst_SboxInst_9_T3}), .c ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, AddRoundConstantOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_9_XOR_o1_U1 ( .a ({new_AGEMA_signal_2771, new_AGEMA_signal_2770, new_AGEMA_signal_2769, SubCellInst_SboxInst_9_YY_1_}), .b ({new_AGEMA_signal_3032, new_AGEMA_signal_3031, new_AGEMA_signal_3030, SubCellInst_SboxInst_9_YY_3}), .c ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, AddRoundConstantOutput[37]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_AND2_U1 ( .a ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}), .b ({new_AGEMA_signal_2582, new_AGEMA_signal_2581, new_AGEMA_signal_2580, SubCellInst_SboxInst_10_Q2}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, SubCellInst_SboxInst_10_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR4_U1 ( .a ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, new_AGEMA_signal_2775, SubCellInst_SboxInst_10_T1}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, new_AGEMA_signal_2409, SubCellInst_SboxInst_10_T2}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, SubCellInst_SboxInst_10_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_AND4_U1 ( .a ({new_AGEMA_signal_2222, new_AGEMA_signal_2221, new_AGEMA_signal_2220, SubCellInst_SboxInst_10_Q6}), .b ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, new_AGEMA_signal_2583, SubCellInst_SboxInst_10_Q7}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, SubCellInst_SboxInst_10_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR9_U1 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, new_AGEMA_signal_2223, SubCellInst_SboxInst_10_L2}), .c ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, SubCellInst_SboxInst_10_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR10_U1 ( .a ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, new_AGEMA_signal_2907, SubCellInst_SboxInst_10_L0}), .b ({new_AGEMA_signal_2780, new_AGEMA_signal_2779, new_AGEMA_signal_2778, SubCellInst_SboxInst_10_T3}), .c ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, AddRoundConstantOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_10_XOR_o1_U1 ( .a ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, new_AGEMA_signal_2781, SubCellInst_SboxInst_10_YY_1_}), .b ({new_AGEMA_signal_3038, new_AGEMA_signal_3037, new_AGEMA_signal_3036, SubCellInst_SboxInst_10_YY_3}), .c ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, AddRoundConstantOutput[41]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_AND2_U1 ( .a ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}), .b ({new_AGEMA_signal_2594, new_AGEMA_signal_2593, new_AGEMA_signal_2592, SubCellInst_SboxInst_11_Q2}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, SubCellInst_SboxInst_11_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR4_U1 ( .a ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, new_AGEMA_signal_2787, SubCellInst_SboxInst_11_T1}), .b ({new_AGEMA_signal_2420, new_AGEMA_signal_2419, new_AGEMA_signal_2418, SubCellInst_SboxInst_11_T2}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, SubCellInst_SboxInst_11_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_AND4_U1 ( .a ({new_AGEMA_signal_2240, new_AGEMA_signal_2239, new_AGEMA_signal_2238, SubCellInst_SboxInst_11_Q6}), .b ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, new_AGEMA_signal_2595, SubCellInst_SboxInst_11_Q7}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, SubCellInst_SboxInst_11_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR9_U1 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, new_AGEMA_signal_2241, SubCellInst_SboxInst_11_L2}), .c ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, SubCellInst_SboxInst_11_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR10_U1 ( .a ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, new_AGEMA_signal_2913, SubCellInst_SboxInst_11_L0}), .b ({new_AGEMA_signal_2792, new_AGEMA_signal_2791, new_AGEMA_signal_2790, SubCellInst_SboxInst_11_T3}), .c ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, SubCellOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_11_XOR_o1_U1 ( .a ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, new_AGEMA_signal_2793, SubCellInst_SboxInst_11_YY_1_}), .b ({new_AGEMA_signal_3044, new_AGEMA_signal_3043, new_AGEMA_signal_3042, SubCellInst_SboxInst_11_YY_3}), .c ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, SubCellOutput[45]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_AND2_U1 ( .a ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}), .b ({new_AGEMA_signal_2606, new_AGEMA_signal_2605, new_AGEMA_signal_2604, SubCellInst_SboxInst_12_Q2}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, SubCellInst_SboxInst_12_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR4_U1 ( .a ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, new_AGEMA_signal_2799, SubCellInst_SboxInst_12_T1}), .b ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, new_AGEMA_signal_2427, SubCellInst_SboxInst_12_T2}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, SubCellInst_SboxInst_12_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_AND4_U1 ( .a ({new_AGEMA_signal_2258, new_AGEMA_signal_2257, new_AGEMA_signal_2256, SubCellInst_SboxInst_12_Q6}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, new_AGEMA_signal_2607, SubCellInst_SboxInst_12_Q7}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, SubCellInst_SboxInst_12_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR9_U1 ( .a ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, new_AGEMA_signal_2259, SubCellInst_SboxInst_12_L2}), .c ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, SubCellInst_SboxInst_12_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR10_U1 ( .a ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, new_AGEMA_signal_2919, SubCellInst_SboxInst_12_L0}), .b ({new_AGEMA_signal_2804, new_AGEMA_signal_2803, new_AGEMA_signal_2802, SubCellInst_SboxInst_12_T3}), .c ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, AddRoundConstantOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_12_XOR_o1_U1 ( .a ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, new_AGEMA_signal_2805, SubCellInst_SboxInst_12_YY_1_}), .b ({new_AGEMA_signal_3050, new_AGEMA_signal_3049, new_AGEMA_signal_3048, SubCellInst_SboxInst_12_YY_3}), .c ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, AddRoundConstantOutput[49]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_AND2_U1 ( .a ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}), .b ({new_AGEMA_signal_2618, new_AGEMA_signal_2617, new_AGEMA_signal_2616, SubCellInst_SboxInst_13_Q2}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, SubCellInst_SboxInst_13_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR4_U1 ( .a ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, new_AGEMA_signal_2811, SubCellInst_SboxInst_13_T1}), .b ({new_AGEMA_signal_2438, new_AGEMA_signal_2437, new_AGEMA_signal_2436, SubCellInst_SboxInst_13_T2}), .c ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, SubCellInst_SboxInst_13_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_AND4_U1 ( .a ({new_AGEMA_signal_2276, new_AGEMA_signal_2275, new_AGEMA_signal_2274, SubCellInst_SboxInst_13_Q6}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, new_AGEMA_signal_2619, SubCellInst_SboxInst_13_Q7}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, SubCellInst_SboxInst_13_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR9_U1 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, new_AGEMA_signal_2277, SubCellInst_SboxInst_13_L2}), .c ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, SubCellInst_SboxInst_13_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR10_U1 ( .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, new_AGEMA_signal_2925, SubCellInst_SboxInst_13_L0}), .b ({new_AGEMA_signal_2816, new_AGEMA_signal_2815, new_AGEMA_signal_2814, SubCellInst_SboxInst_13_T3}), .c ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, AddRoundConstantOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_13_XOR_o1_U1 ( .a ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, new_AGEMA_signal_2817, SubCellInst_SboxInst_13_YY_1_}), .b ({new_AGEMA_signal_3056, new_AGEMA_signal_3055, new_AGEMA_signal_3054, SubCellInst_SboxInst_13_YY_3}), .c ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, AddRoundConstantOutput[53]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_AND2_U1 ( .a ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}), .b ({new_AGEMA_signal_2630, new_AGEMA_signal_2629, new_AGEMA_signal_2628, SubCellInst_SboxInst_14_Q2}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, SubCellInst_SboxInst_14_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR4_U1 ( .a ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, new_AGEMA_signal_2823, SubCellInst_SboxInst_14_T1}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, new_AGEMA_signal_2445, SubCellInst_SboxInst_14_T2}), .c ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, SubCellInst_SboxInst_14_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_AND4_U1 ( .a ({new_AGEMA_signal_2294, new_AGEMA_signal_2293, new_AGEMA_signal_2292, SubCellInst_SboxInst_14_Q6}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, new_AGEMA_signal_2631, SubCellInst_SboxInst_14_Q7}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, SubCellInst_SboxInst_14_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR9_U1 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, new_AGEMA_signal_2295, SubCellInst_SboxInst_14_L2}), .c ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, SubCellInst_SboxInst_14_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR10_U1 ( .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, new_AGEMA_signal_2931, SubCellInst_SboxInst_14_L0}), .b ({new_AGEMA_signal_2828, new_AGEMA_signal_2827, new_AGEMA_signal_2826, SubCellInst_SboxInst_14_T3}), .c ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, AddRoundConstantOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_14_XOR_o1_U1 ( .a ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, new_AGEMA_signal_2829, SubCellInst_SboxInst_14_YY_1_}), .b ({new_AGEMA_signal_3062, new_AGEMA_signal_3061, new_AGEMA_signal_3060, SubCellInst_SboxInst_14_YY_3}), .c ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, AddRoundConstantOutput[57]}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_AND2_U1 ( .a ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}), .b ({new_AGEMA_signal_2642, new_AGEMA_signal_2641, new_AGEMA_signal_2640, SubCellInst_SboxInst_15_Q2}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, SubCellInst_SboxInst_15_T1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR4_U1 ( .a ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, new_AGEMA_signal_2835, SubCellInst_SboxInst_15_T1}), .b ({new_AGEMA_signal_2456, new_AGEMA_signal_2455, new_AGEMA_signal_2454, SubCellInst_SboxInst_15_T2}), .c ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, SubCellInst_SboxInst_15_L0}) ) ;
    and_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_AND4_U1 ( .a ({new_AGEMA_signal_2312, new_AGEMA_signal_2311, new_AGEMA_signal_2310, SubCellInst_SboxInst_15_Q6}), .b ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, new_AGEMA_signal_2643, SubCellInst_SboxInst_15_Q7}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, SubCellInst_SboxInst_15_T3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR9_U1 ( .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, new_AGEMA_signal_2313, SubCellInst_SboxInst_15_L2}), .c ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, SubCellInst_SboxInst_15_YY_3}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR10_U1 ( .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, new_AGEMA_signal_2937, SubCellInst_SboxInst_15_L0}), .b ({new_AGEMA_signal_2840, new_AGEMA_signal_2839, new_AGEMA_signal_2838, SubCellInst_SboxInst_15_T3}), .c ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, SubCellOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) SubCellInst_SboxInst_15_XOR_o1_U1 ( .a ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, new_AGEMA_signal_2841, SubCellInst_SboxInst_15_YY_1_}), .b ({new_AGEMA_signal_3068, new_AGEMA_signal_3067, new_AGEMA_signal_3066, SubCellInst_SboxInst_15_YY_3}), .c ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, SubCellOutput[61]}) ) ;
    not_masked #(.security_order(3), .pipeline(0)) AddConstXOR_U2 ( .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, new_AGEMA_signal_3171, SubCellOutput[29]}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, AddConstXOR_AddConstXOR_XORInst_0_0_n1}), .b ({1'b0, 1'b0, 1'b0, FSMUpdate[1]}), .c ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, AddRoundConstantOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, new_AGEMA_signal_3069, SubCellOutput[60]}), .c ({new_AGEMA_signal_3200, new_AGEMA_signal_3199, new_AGEMA_signal_3198, AddConstXOR_AddConstXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, AddConstXOR_AddConstXOR_XORInst_0_1_n1}), .b ({1'b0, 1'b0, 1'b0, FSM[1]}), .c ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, AddRoundConstantOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, new_AGEMA_signal_3195, SubCellOutput[61]}), .c ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, new_AGEMA_signal_3315, AddConstXOR_AddConstXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, AddConstXOR_AddConstXOR_XORInst_1_0_n1}), .b ({1'b0, 1'b0, 1'b0, FSM[4]}), .c ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, AddRoundConstantOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, new_AGEMA_signal_3045, SubCellOutput[44]}), .c ({new_AGEMA_signal_3206, new_AGEMA_signal_3205, new_AGEMA_signal_3204, AddConstXOR_AddConstXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, AddConstXOR_AddConstXOR_XORInst_1_1_n1}), .b ({1'b0, 1'b0, 1'b0, FSM[5]}), .c ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, AddRoundConstantOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddConstXOR_AddConstXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, new_AGEMA_signal_3183, SubCellOutput[45]}), .c ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, new_AGEMA_signal_3321, AddConstXOR_AddConstXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, AddRoundTweakeyXOR_XORInst_0_0_n1}), .b ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[0]}), .c ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, ShiftRowsOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, new_AGEMA_signal_3027, AddRoundConstantOutput[32]}), .c ({new_AGEMA_signal_3212, new_AGEMA_signal_3211, new_AGEMA_signal_3210, AddRoundTweakeyXOR_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, AddRoundTweakeyXOR_XORInst_0_1_n1}), .b ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, TweakeyGeneration_key_Feedback[1]}), .c ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, ShiftRowsOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3176, new_AGEMA_signal_3175, new_AGEMA_signal_3174, AddRoundConstantOutput[33]}), .c ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, new_AGEMA_signal_3327, AddRoundTweakeyXOR_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, AddRoundTweakeyXOR_XORInst_1_0_n1}), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[4]}), .c ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, ShiftRowsOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, new_AGEMA_signal_3033, AddRoundConstantOutput[36]}), .c ({new_AGEMA_signal_3218, new_AGEMA_signal_3217, new_AGEMA_signal_3216, AddRoundTweakeyXOR_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, AddRoundTweakeyXOR_XORInst_1_1_n1}), .b ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, TweakeyGeneration_key_Feedback[5]}), .c ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, ShiftRowsOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, new_AGEMA_signal_3177, AddRoundConstantOutput[37]}), .c ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, new_AGEMA_signal_3333, AddRoundTweakeyXOR_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, AddRoundTweakeyXOR_XORInst_2_0_n1}), .b ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[8]}), .c ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, ShiftRowsOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, new_AGEMA_signal_3039, AddRoundConstantOutput[40]}), .c ({new_AGEMA_signal_3224, new_AGEMA_signal_3223, new_AGEMA_signal_3222, AddRoundTweakeyXOR_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, AddRoundTweakeyXOR_XORInst_2_1_n1}), .b ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, TweakeyGeneration_key_Feedback[9]}), .c ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, ShiftRowsOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3182, new_AGEMA_signal_3181, new_AGEMA_signal_3180, AddRoundConstantOutput[41]}), .c ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, new_AGEMA_signal_3339, AddRoundTweakeyXOR_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, AddRoundTweakeyXOR_XORInst_3_0_n1}), .b ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[12]}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, ShiftRowsOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3320, new_AGEMA_signal_3319, new_AGEMA_signal_3318, AddRoundConstantOutput[44]}), .c ({new_AGEMA_signal_3530, new_AGEMA_signal_3529, new_AGEMA_signal_3528, AddRoundTweakeyXOR_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, AddRoundTweakeyXOR_XORInst_3_1_n1}), .b ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, TweakeyGeneration_key_Feedback[13]}), .c ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, new_AGEMA_signal_3855, ShiftRowsOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3518, new_AGEMA_signal_3517, new_AGEMA_signal_3516, AddRoundConstantOutput[45]}), .c ({new_AGEMA_signal_3698, new_AGEMA_signal_3697, new_AGEMA_signal_3696, AddRoundTweakeyXOR_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_0_U2 ( .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, AddRoundTweakeyXOR_XORInst_4_0_n1}), .b ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[16]}), .c ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, new_AGEMA_signal_3051, AddRoundConstantOutput[48]}), .c ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, new_AGEMA_signal_3231, AddRoundTweakeyXOR_XORInst_4_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_1_U2 ( .a ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, AddRoundTweakeyXOR_XORInst_4_1_n1}), .b ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, TweakeyGeneration_key_Feedback[17]}), .c ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_4_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3188, new_AGEMA_signal_3187, new_AGEMA_signal_3186, AddRoundConstantOutput[49]}), .c ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, new_AGEMA_signal_3351, AddRoundTweakeyXOR_XORInst_4_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_0_U2 ( .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, AddRoundTweakeyXOR_XORInst_5_0_n1}), .b ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[20]}), .c ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, new_AGEMA_signal_3057, AddRoundConstantOutput[52]}), .c ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, new_AGEMA_signal_3237, AddRoundTweakeyXOR_XORInst_5_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_1_U2 ( .a ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, AddRoundTweakeyXOR_XORInst_5_1_n1}), .b ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, TweakeyGeneration_key_Feedback[21]}), .c ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_5_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, new_AGEMA_signal_3189, AddRoundConstantOutput[53]}), .c ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, new_AGEMA_signal_3357, AddRoundTweakeyXOR_XORInst_5_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_0_U2 ( .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, AddRoundTweakeyXOR_XORInst_6_0_n1}), .b ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[24]}), .c ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, new_AGEMA_signal_3063, AddRoundConstantOutput[56]}), .c ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, new_AGEMA_signal_3243, AddRoundTweakeyXOR_XORInst_6_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_1_U2 ( .a ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, AddRoundTweakeyXOR_XORInst_6_1_n1}), .b ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, TweakeyGeneration_key_Feedback[25]}), .c ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_6_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3194, new_AGEMA_signal_3193, new_AGEMA_signal_3192, AddRoundConstantOutput[57]}), .c ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, new_AGEMA_signal_3363, AddRoundTweakeyXOR_XORInst_6_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_0_U2 ( .a ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, AddRoundTweakeyXOR_XORInst_7_0_n1}), .b ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[28]}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3314, new_AGEMA_signal_3313, new_AGEMA_signal_3312, AddRoundConstantOutput[60]}), .c ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, new_AGEMA_signal_3543, AddRoundTweakeyXOR_XORInst_7_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_1_U2 ( .a ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, AddRoundTweakeyXOR_XORInst_7_1_n1}), .b ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, TweakeyGeneration_key_Feedback[29]}), .c ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) AddRoundTweakeyXOR_XORInst_7_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, new_AGEMA_signal_3513, AddRoundConstantOutput[61]}), .c ({new_AGEMA_signal_3704, new_AGEMA_signal_3703, new_AGEMA_signal_3702, AddRoundTweakeyXOR_XORInst_7_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U3 ( .a ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, MCInst_MCR0_XORInst_0_0_n2}), .b ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, MCInst_MCR0_XORInst_0_0_n1}), .c ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, new_AGEMA_signal_3705, MCOutput[48]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}), .b ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, new_AGEMA_signal_2997, ShiftRowsOutput[0]}), .c ({new_AGEMA_signal_3254, new_AGEMA_signal_3253, new_AGEMA_signal_3252, MCInst_MCR0_XORInst_0_0_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}), .c ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, new_AGEMA_signal_3549, MCInst_MCR0_XORInst_0_0_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U3 ( .a ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, MCInst_MCR0_XORInst_0_1_n2}), .b ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, MCInst_MCR0_XORInst_0_1_n1}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, new_AGEMA_signal_3861, MCOutput[49]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}), .b ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, new_AGEMA_signal_3159, ShiftRowsOutput[1]}), .c ({new_AGEMA_signal_3374, new_AGEMA_signal_3373, new_AGEMA_signal_3372, MCInst_MCR0_XORInst_0_1_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}), .c ({new_AGEMA_signal_3710, new_AGEMA_signal_3709, new_AGEMA_signal_3708, MCInst_MCR0_XORInst_0_1_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U3 ( .a ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, MCInst_MCR0_XORInst_1_0_n2}), .b ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, MCInst_MCR0_XORInst_1_0_n1}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, new_AGEMA_signal_3711, MCOutput[52]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, new_AGEMA_signal_2979, ShiftRowsOutput[4]}), .c ({new_AGEMA_signal_3260, new_AGEMA_signal_3259, new_AGEMA_signal_3258, MCInst_MCR0_XORInst_1_0_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}), .c ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, new_AGEMA_signal_3555, MCInst_MCR0_XORInst_1_0_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U3 ( .a ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, MCInst_MCR0_XORInst_1_1_n2}), .b ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, MCInst_MCR0_XORInst_1_1_n1}), .c ({new_AGEMA_signal_3866, new_AGEMA_signal_3865, new_AGEMA_signal_3864, MCOutput[53]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}), .b ({new_AGEMA_signal_3152, new_AGEMA_signal_3151, new_AGEMA_signal_3150, ShiftRowsOutput[5]}), .c ({new_AGEMA_signal_3560, new_AGEMA_signal_3559, new_AGEMA_signal_3558, MCInst_MCR0_XORInst_1_1_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}), .c ({new_AGEMA_signal_3716, new_AGEMA_signal_3715, new_AGEMA_signal_3714, MCInst_MCR0_XORInst_1_1_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U3 ( .a ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, MCInst_MCR0_XORInst_2_0_n2}), .b ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, MCInst_MCR0_XORInst_2_0_n1}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, new_AGEMA_signal_3717, MCOutput[56]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, new_AGEMA_signal_2985, ShiftRowsOutput[8]}), .c ({new_AGEMA_signal_3266, new_AGEMA_signal_3265, new_AGEMA_signal_3264, MCInst_MCR0_XORInst_2_0_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}), .c ({new_AGEMA_signal_3566, new_AGEMA_signal_3565, new_AGEMA_signal_3564, MCInst_MCR0_XORInst_2_0_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U3 ( .a ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, MCInst_MCR0_XORInst_2_1_n2}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, MCInst_MCR0_XORInst_2_1_n1}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, new_AGEMA_signal_3867, MCOutput[57]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, new_AGEMA_signal_3153, ShiftRowsOutput[9]}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, new_AGEMA_signal_3387, MCInst_MCR0_XORInst_2_1_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}), .c ({new_AGEMA_signal_3722, new_AGEMA_signal_3721, new_AGEMA_signal_3720, MCInst_MCR0_XORInst_2_1_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U3 ( .a ({new_AGEMA_signal_3872, new_AGEMA_signal_3871, new_AGEMA_signal_3870, MCInst_MCR0_XORInst_3_0_n2}), .b ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, MCInst_MCR0_XORInst_3_0_n1}), .c ({new_AGEMA_signal_3986, new_AGEMA_signal_3985, new_AGEMA_signal_3984, MCOutput[60]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}), .b ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, new_AGEMA_signal_2991, ShiftRowsOutput[12]}), .c ({new_AGEMA_signal_3272, new_AGEMA_signal_3271, new_AGEMA_signal_3270, MCInst_MCR0_XORInst_3_0_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}), .c ({new_AGEMA_signal_3872, new_AGEMA_signal_3871, new_AGEMA_signal_3870, MCInst_MCR0_XORInst_3_0_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U3 ( .a ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, new_AGEMA_signal_3987, MCInst_MCR0_XORInst_3_1_n2}), .b ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, MCInst_MCR0_XORInst_3_1_n1}), .c ({new_AGEMA_signal_4022, new_AGEMA_signal_4021, new_AGEMA_signal_4020, MCOutput[61]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}), .b ({new_AGEMA_signal_3158, new_AGEMA_signal_3157, new_AGEMA_signal_3156, ShiftRowsOutput[13]}), .c ({new_AGEMA_signal_3398, new_AGEMA_signal_3397, new_AGEMA_signal_3396, MCInst_MCR0_XORInst_3_1_n1}) ) ;
    xor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR0_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}), .c ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, new_AGEMA_signal_3987, MCInst_MCR0_XORInst_3_1_n2}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, MCInst_MCR2_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, new_AGEMA_signal_3729, MCOutput[16]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3332, new_AGEMA_signal_3331, new_AGEMA_signal_3330, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, new_AGEMA_signal_3573, MCInst_MCR2_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, new_AGEMA_signal_3732, MCInst_MCR2_XORInst_0_1_n1}), .b ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_3878, new_AGEMA_signal_3877, new_AGEMA_signal_3876, MCOutput[17]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3524, new_AGEMA_signal_3523, new_AGEMA_signal_3522, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_3734, new_AGEMA_signal_3733, new_AGEMA_signal_3732, MCInst_MCR2_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, MCInst_MCR2_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, new_AGEMA_signal_3735, MCOutput[20]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3338, new_AGEMA_signal_3337, new_AGEMA_signal_3336, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, new_AGEMA_signal_3579, MCInst_MCR2_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738, MCInst_MCR2_XORInst_1_1_n1}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, new_AGEMA_signal_3879, MCOutput[21]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, new_AGEMA_signal_3525, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_3740, new_AGEMA_signal_3739, new_AGEMA_signal_3738, MCInst_MCR2_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, new_AGEMA_signal_3882, MCInst_MCR2_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_3992, new_AGEMA_signal_3991, new_AGEMA_signal_3990, MCOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, new_AGEMA_signal_3693, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_3884, new_AGEMA_signal_3883, new_AGEMA_signal_3882, MCInst_MCR2_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, new_AGEMA_signal_3993, MCInst_MCR2_XORInst_2_1_n1}), .b ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, new_AGEMA_signal_4023, MCOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, new_AGEMA_signal_3855, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, new_AGEMA_signal_3993, MCInst_MCR2_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, MCInst_MCR2_XORInst_3_0_n1}), .b ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, new_AGEMA_signal_3747, MCOutput[28]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3326, new_AGEMA_signal_3325, new_AGEMA_signal_3324, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_3590, new_AGEMA_signal_3589, new_AGEMA_signal_3588, MCInst_MCR2_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750, MCInst_MCR2_XORInst_3_1_n1}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_3890, new_AGEMA_signal_3889, new_AGEMA_signal_3888, MCOutput[29]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR2_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, new_AGEMA_signal_3519, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_3752, new_AGEMA_signal_3751, new_AGEMA_signal_3750, MCInst_MCR2_XORInst_3_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_0_U2 ( .a ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, MCInst_MCR3_XORInst_0_0_n1}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, new_AGEMA_signal_3015, ShiftRowsOutput[16]}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, new_AGEMA_signal_3753, MCOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3350, new_AGEMA_signal_3349, new_AGEMA_signal_3348, MCOutput[32]}), .c ({new_AGEMA_signal_3596, new_AGEMA_signal_3595, new_AGEMA_signal_3594, MCInst_MCR3_XORInst_0_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_1_U2 ( .a ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, new_AGEMA_signal_3756, MCInst_MCR3_XORInst_0_1_n1}), .b ({new_AGEMA_signal_3170, new_AGEMA_signal_3169, new_AGEMA_signal_3168, ShiftRowsOutput[17]}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, new_AGEMA_signal_3891, MCOutput[1]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_0_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3536, new_AGEMA_signal_3535, new_AGEMA_signal_3534, MCOutput[33]}), .c ({new_AGEMA_signal_3758, new_AGEMA_signal_3757, new_AGEMA_signal_3756, MCInst_MCR3_XORInst_0_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_0_U2 ( .a ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, MCInst_MCR3_XORInst_1_0_n1}), .b ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, new_AGEMA_signal_3021, ShiftRowsOutput[20]}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, new_AGEMA_signal_3759, MCOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3356, new_AGEMA_signal_3355, new_AGEMA_signal_3354, MCOutput[36]}), .c ({new_AGEMA_signal_3602, new_AGEMA_signal_3601, new_AGEMA_signal_3600, MCInst_MCR3_XORInst_1_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_1_U2 ( .a ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, new_AGEMA_signal_3762, MCInst_MCR3_XORInst_1_1_n1}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, new_AGEMA_signal_3309, ShiftRowsOutput[21]}), .c ({new_AGEMA_signal_3896, new_AGEMA_signal_3895, new_AGEMA_signal_3894, MCOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_1_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, new_AGEMA_signal_3537, MCOutput[37]}), .c ({new_AGEMA_signal_3764, new_AGEMA_signal_3763, new_AGEMA_signal_3762, MCInst_MCR3_XORInst_1_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_0_U2 ( .a ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, MCInst_MCR3_XORInst_2_0_n1}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, new_AGEMA_signal_3003, ShiftRowsOutput[24]}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, new_AGEMA_signal_3765, MCOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3362, new_AGEMA_signal_3361, new_AGEMA_signal_3360, MCOutput[40]}), .c ({new_AGEMA_signal_3608, new_AGEMA_signal_3607, new_AGEMA_signal_3606, MCInst_MCR3_XORInst_2_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_1_U2 ( .a ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, new_AGEMA_signal_3768, MCInst_MCR3_XORInst_2_1_n1}), .b ({new_AGEMA_signal_3164, new_AGEMA_signal_3163, new_AGEMA_signal_3162, ShiftRowsOutput[25]}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, new_AGEMA_signal_3897, MCOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_2_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3542, new_AGEMA_signal_3541, new_AGEMA_signal_3540, MCOutput[41]}), .c ({new_AGEMA_signal_3770, new_AGEMA_signal_3769, new_AGEMA_signal_3768, MCInst_MCR3_XORInst_2_1_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_0_U2 ( .a ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, new_AGEMA_signal_3900, MCInst_MCR3_XORInst_3_0_n1}), .b ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, new_AGEMA_signal_3009, ShiftRowsOutput[28]}), .c ({new_AGEMA_signal_3998, new_AGEMA_signal_3997, new_AGEMA_signal_3996, MCOutput[12]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_0_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, new_AGEMA_signal_3699, MCOutput[44]}), .c ({new_AGEMA_signal_3902, new_AGEMA_signal_3901, new_AGEMA_signal_3900, MCInst_MCR3_XORInst_3_0_n1}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_1_U2 ( .a ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, new_AGEMA_signal_3999, MCInst_MCR3_XORInst_3_1_n1}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, new_AGEMA_signal_3165, ShiftRowsOutput[29]}), .c ({new_AGEMA_signal_4028, new_AGEMA_signal_4027, new_AGEMA_signal_4026, MCOutput[13]}) ) ;
    xnor_HPC3 #(.security_order(3), .pipeline(0)) MCInst_MCR3_XORInst_3_1_U1 ( .a ({1'b0, 1'b0, 1'b0, 1'b0}), .b ({new_AGEMA_signal_3860, new_AGEMA_signal_3859, new_AGEMA_signal_3858, MCOutput[45]}), .c ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, new_AGEMA_signal_3999, MCInst_MCR3_XORInst_3_1_n1}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, new_AGEMA_signal_3981, StateRegInput[63]}), .Q ({Ciphertext_s3[63], Ciphertext_s2[63], Ciphertext_s1[63], Ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3854, new_AGEMA_signal_3853, new_AGEMA_signal_3852, StateRegInput[62]}), .Q ({Ciphertext_s3[62], Ciphertext_s2[62], Ciphertext_s1[62], Ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4046, new_AGEMA_signal_4045, new_AGEMA_signal_4044, StateRegInput[61]}), .Q ({Ciphertext_s3[61], Ciphertext_s2[61], Ciphertext_s1[61], Ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, new_AGEMA_signal_4017, StateRegInput[60]}), .Q ({Ciphertext_s3[60], Ciphertext_s2[60], Ciphertext_s1[60], Ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3692, new_AGEMA_signal_3691, new_AGEMA_signal_3690, StateRegInput[59]}), .Q ({Ciphertext_s3[59], Ciphertext_s2[59], Ciphertext_s1[59], Ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3512, new_AGEMA_signal_3511, new_AGEMA_signal_3510, StateRegInput[58]}), .Q ({Ciphertext_s3[58], Ciphertext_s2[58], Ciphertext_s1[58], Ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, new_AGEMA_signal_3975, StateRegInput[57]}), .Q ({Ciphertext_s3[57], Ciphertext_s2[57], Ciphertext_s1[57], Ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3848, new_AGEMA_signal_3847, new_AGEMA_signal_3846, StateRegInput[56]}), .Q ({Ciphertext_s3[56], Ciphertext_s2[56], Ciphertext_s1[56], Ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3686, new_AGEMA_signal_3685, new_AGEMA_signal_3684, StateRegInput[55]}), .Q ({Ciphertext_s3[55], Ciphertext_s2[55], Ciphertext_s1[55], Ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3506, new_AGEMA_signal_3505, new_AGEMA_signal_3504, StateRegInput[54]}), .Q ({Ciphertext_s3[54], Ciphertext_s2[54], Ciphertext_s1[54], Ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, new_AGEMA_signal_3969, StateRegInput[53]}), .Q ({Ciphertext_s3[53], Ciphertext_s2[53], Ciphertext_s1[53], Ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3842, new_AGEMA_signal_3841, new_AGEMA_signal_3840, StateRegInput[52]}), .Q ({Ciphertext_s3[52], Ciphertext_s2[52], Ciphertext_s1[52], Ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3680, new_AGEMA_signal_3679, new_AGEMA_signal_3678, StateRegInput[51]}), .Q ({Ciphertext_s3[51], Ciphertext_s2[51], Ciphertext_s1[51], Ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3500, new_AGEMA_signal_3499, new_AGEMA_signal_3498, StateRegInput[50]}), .Q ({Ciphertext_s3[50], Ciphertext_s2[50], Ciphertext_s1[50], Ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, new_AGEMA_signal_3963, StateRegInput[49]}), .Q ({Ciphertext_s3[49], Ciphertext_s2[49], Ciphertext_s1[49], Ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3836, new_AGEMA_signal_3835, new_AGEMA_signal_3834, StateRegInput[48]}), .Q ({Ciphertext_s3[48], Ciphertext_s2[48], Ciphertext_s1[48], Ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3674, new_AGEMA_signal_3673, new_AGEMA_signal_3672, StateRegInput[47]}), .Q ({Ciphertext_s3[47], Ciphertext_s2[47], Ciphertext_s1[47], Ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3494, new_AGEMA_signal_3493, new_AGEMA_signal_3492, StateRegInput[46]}), .Q ({Ciphertext_s3[46], Ciphertext_s2[46], Ciphertext_s1[46], Ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, new_AGEMA_signal_3957, StateRegInput[45]}), .Q ({Ciphertext_s3[45], Ciphertext_s2[45], Ciphertext_s1[45], Ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3830, new_AGEMA_signal_3829, new_AGEMA_signal_3828, StateRegInput[44]}), .Q ({Ciphertext_s3[44], Ciphertext_s2[44], Ciphertext_s1[44], Ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3308, new_AGEMA_signal_3307, new_AGEMA_signal_3306, StateRegInput[43]}), .Q ({Ciphertext_s3[43], Ciphertext_s2[43], Ciphertext_s1[43], Ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, new_AGEMA_signal_3147, StateRegInput[42]}), .Q ({Ciphertext_s3[42], Ciphertext_s2[42], Ciphertext_s1[42], Ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3668, new_AGEMA_signal_3667, new_AGEMA_signal_3666, StateRegInput[41]}), .Q ({Ciphertext_s3[41], Ciphertext_s2[41], Ciphertext_s1[41], Ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3488, new_AGEMA_signal_3487, new_AGEMA_signal_3486, StateRegInput[40]}), .Q ({Ciphertext_s3[40], Ciphertext_s2[40], Ciphertext_s1[40], Ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3302, new_AGEMA_signal_3301, new_AGEMA_signal_3300, StateRegInput[39]}), .Q ({Ciphertext_s3[39], Ciphertext_s2[39], Ciphertext_s1[39], Ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, new_AGEMA_signal_3141, StateRegInput[38]}), .Q ({Ciphertext_s3[38], Ciphertext_s2[38], Ciphertext_s1[38], Ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3662, new_AGEMA_signal_3661, new_AGEMA_signal_3660, StateRegInput[37]}), .Q ({Ciphertext_s3[37], Ciphertext_s2[37], Ciphertext_s1[37], Ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3482, new_AGEMA_signal_3481, new_AGEMA_signal_3480, StateRegInput[36]}), .Q ({Ciphertext_s3[36], Ciphertext_s2[36], Ciphertext_s1[36], Ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3296, new_AGEMA_signal_3295, new_AGEMA_signal_3294, StateRegInput[35]}), .Q ({Ciphertext_s3[35], Ciphertext_s2[35], Ciphertext_s1[35], Ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, new_AGEMA_signal_3135, StateRegInput[34]}), .Q ({Ciphertext_s3[34], Ciphertext_s2[34], Ciphertext_s1[34], Ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3656, new_AGEMA_signal_3655, new_AGEMA_signal_3654, StateRegInput[33]}), .Q ({Ciphertext_s3[33], Ciphertext_s2[33], Ciphertext_s1[33], Ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3476, new_AGEMA_signal_3475, new_AGEMA_signal_3474, StateRegInput[32]}), .Q ({Ciphertext_s3[32], Ciphertext_s2[32], Ciphertext_s1[32], Ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3650, new_AGEMA_signal_3649, new_AGEMA_signal_3648, StateRegInput[31]}), .Q ({Ciphertext_s3[31], Ciphertext_s2[31], Ciphertext_s1[31], Ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3470, new_AGEMA_signal_3469, new_AGEMA_signal_3468, StateRegInput[30]}), .Q ({Ciphertext_s3[30], Ciphertext_s2[30], Ciphertext_s1[30], Ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, new_AGEMA_signal_3951, StateRegInput[29]}), .Q ({Ciphertext_s3[29], Ciphertext_s2[29], Ciphertext_s1[29], Ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3824, new_AGEMA_signal_3823, new_AGEMA_signal_3822, StateRegInput[28]}), .Q ({Ciphertext_s3[28], Ciphertext_s2[28], Ciphertext_s1[28], Ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, new_AGEMA_signal_3945, StateRegInput[27]}), .Q ({Ciphertext_s3[27], Ciphertext_s2[27], Ciphertext_s1[27], Ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3818, new_AGEMA_signal_3817, new_AGEMA_signal_3816, StateRegInput[26]}), .Q ({Ciphertext_s3[26], Ciphertext_s2[26], Ciphertext_s1[26], Ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4040, new_AGEMA_signal_4039, new_AGEMA_signal_4038, StateRegInput[25]}), .Q ({Ciphertext_s3[25], Ciphertext_s2[25], Ciphertext_s1[25], Ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, new_AGEMA_signal_4011, StateRegInput[24]}), .Q ({Ciphertext_s3[24], Ciphertext_s2[24], Ciphertext_s1[24], Ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3644, new_AGEMA_signal_3643, new_AGEMA_signal_3642, StateRegInput[23]}), .Q ({Ciphertext_s3[23], Ciphertext_s2[23], Ciphertext_s1[23], Ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3464, new_AGEMA_signal_3463, new_AGEMA_signal_3462, StateRegInput[22]}), .Q ({Ciphertext_s3[22], Ciphertext_s2[22], Ciphertext_s1[22], Ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, new_AGEMA_signal_3939, StateRegInput[21]}), .Q ({Ciphertext_s3[21], Ciphertext_s2[21], Ciphertext_s1[21], Ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3812, new_AGEMA_signal_3811, new_AGEMA_signal_3810, StateRegInput[20]}), .Q ({Ciphertext_s3[20], Ciphertext_s2[20], Ciphertext_s1[20], Ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3638, new_AGEMA_signal_3637, new_AGEMA_signal_3636, StateRegInput[19]}), .Q ({Ciphertext_s3[19], Ciphertext_s2[19], Ciphertext_s1[19], Ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3458, new_AGEMA_signal_3457, new_AGEMA_signal_3456, StateRegInput[18]}), .Q ({Ciphertext_s3[18], Ciphertext_s2[18], Ciphertext_s1[18], Ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, new_AGEMA_signal_3933, StateRegInput[17]}), .Q ({Ciphertext_s3[17], Ciphertext_s2[17], Ciphertext_s1[17], Ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3806, new_AGEMA_signal_3805, new_AGEMA_signal_3804, StateRegInput[16]}), .Q ({Ciphertext_s3[16], Ciphertext_s2[16], Ciphertext_s1[16], Ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, new_AGEMA_signal_3927, StateRegInput[15]}), .Q ({Ciphertext_s3[15], Ciphertext_s2[15], Ciphertext_s1[15], Ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3800, new_AGEMA_signal_3799, new_AGEMA_signal_3798, StateRegInput[14]}), .Q ({Ciphertext_s3[14], Ciphertext_s2[14], Ciphertext_s1[14], Ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4034, new_AGEMA_signal_4033, new_AGEMA_signal_4032, StateRegInput[13]}), .Q ({Ciphertext_s3[13], Ciphertext_s2[13], Ciphertext_s1[13], Ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, new_AGEMA_signal_4005, StateRegInput[12]}), .Q ({Ciphertext_s3[12], Ciphertext_s2[12], Ciphertext_s1[12], Ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3632, new_AGEMA_signal_3631, new_AGEMA_signal_3630, StateRegInput[11]}), .Q ({Ciphertext_s3[11], Ciphertext_s2[11], Ciphertext_s1[11], Ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3452, new_AGEMA_signal_3451, new_AGEMA_signal_3450, StateRegInput[10]}), .Q ({Ciphertext_s3[10], Ciphertext_s2[10], Ciphertext_s1[10], Ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, new_AGEMA_signal_3921, StateRegInput[9]}), .Q ({Ciphertext_s3[9], Ciphertext_s2[9], Ciphertext_s1[9], Ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3794, new_AGEMA_signal_3793, new_AGEMA_signal_3792, StateRegInput[8]}), .Q ({Ciphertext_s3[8], Ciphertext_s2[8], Ciphertext_s1[8], Ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3626, new_AGEMA_signal_3625, new_AGEMA_signal_3624, StateRegInput[7]}), .Q ({Ciphertext_s3[7], Ciphertext_s2[7], Ciphertext_s1[7], Ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3446, new_AGEMA_signal_3445, new_AGEMA_signal_3444, StateRegInput[6]}), .Q ({Ciphertext_s3[6], Ciphertext_s2[6], Ciphertext_s1[6], Ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, new_AGEMA_signal_3915, StateRegInput[5]}), .Q ({Ciphertext_s3[5], Ciphertext_s2[5], Ciphertext_s1[5], Ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3788, new_AGEMA_signal_3787, new_AGEMA_signal_3786, StateRegInput[4]}), .Q ({Ciphertext_s3[4], Ciphertext_s2[4], Ciphertext_s1[4], Ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3620, new_AGEMA_signal_3619, new_AGEMA_signal_3618, StateRegInput[3]}), .Q ({Ciphertext_s3[3], Ciphertext_s2[3], Ciphertext_s1[3], Ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3440, new_AGEMA_signal_3439, new_AGEMA_signal_3438, StateRegInput[2]}), .Q ({Ciphertext_s3[2], Ciphertext_s2[2], Ciphertext_s1[2], Ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, new_AGEMA_signal_3909, StateRegInput[1]}), .Q ({Ciphertext_s3[1], Ciphertext_s2[1], Ciphertext_s1[1], Ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_3782, new_AGEMA_signal_3781, new_AGEMA_signal_3780, StateRegInput[0]}), .Q ({Ciphertext_s3[0], Ciphertext_s2[0], Ciphertext_s1[0], Ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_63__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, new_AGEMA_signal_2025, TweakeyGeneration_StateRegInput[63]}), .Q ({new_AGEMA_signal_1733, new_AGEMA_signal_1732, new_AGEMA_signal_1731, TweakeyGeneration_key_Feedback[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_62__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2018, new_AGEMA_signal_2017, new_AGEMA_signal_2016, TweakeyGeneration_StateRegInput[62]}), .Q ({new_AGEMA_signal_1724, new_AGEMA_signal_1723, new_AGEMA_signal_1722, TweakeyGeneration_key_Feedback[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_61__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, new_AGEMA_signal_2007, TweakeyGeneration_StateRegInput[61]}), .Q ({new_AGEMA_signal_1715, new_AGEMA_signal_1714, new_AGEMA_signal_1713, TweakeyGeneration_key_Feedback[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_60__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_2000, new_AGEMA_signal_1999, new_AGEMA_signal_1998, TweakeyGeneration_StateRegInput[60]}), .Q ({new_AGEMA_signal_1706, new_AGEMA_signal_1705, new_AGEMA_signal_1704, TweakeyGeneration_key_Feedback[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_59__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, new_AGEMA_signal_1989, TweakeyGeneration_StateRegInput[59]}), .Q ({new_AGEMA_signal_1697, new_AGEMA_signal_1696, new_AGEMA_signal_1695, TweakeyGeneration_key_Feedback[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_58__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1982, new_AGEMA_signal_1981, new_AGEMA_signal_1980, TweakeyGeneration_StateRegInput[58]}), .Q ({new_AGEMA_signal_1688, new_AGEMA_signal_1687, new_AGEMA_signal_1686, TweakeyGeneration_key_Feedback[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_57__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1973, new_AGEMA_signal_1972, new_AGEMA_signal_1971, TweakeyGeneration_StateRegInput[57]}), .Q ({new_AGEMA_signal_1679, new_AGEMA_signal_1678, new_AGEMA_signal_1677, TweakeyGeneration_key_Feedback[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_56__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1964, new_AGEMA_signal_1963, new_AGEMA_signal_1962, TweakeyGeneration_StateRegInput[56]}), .Q ({new_AGEMA_signal_1670, new_AGEMA_signal_1669, new_AGEMA_signal_1668, TweakeyGeneration_key_Feedback[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_55__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1955, new_AGEMA_signal_1954, new_AGEMA_signal_1953, TweakeyGeneration_StateRegInput[55]}), .Q ({new_AGEMA_signal_1661, new_AGEMA_signal_1660, new_AGEMA_signal_1659, TweakeyGeneration_key_Feedback[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_54__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1946, new_AGEMA_signal_1945, new_AGEMA_signal_1944, TweakeyGeneration_StateRegInput[54]}), .Q ({new_AGEMA_signal_1652, new_AGEMA_signal_1651, new_AGEMA_signal_1650, TweakeyGeneration_key_Feedback[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_53__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1937, new_AGEMA_signal_1936, new_AGEMA_signal_1935, TweakeyGeneration_StateRegInput[53]}), .Q ({new_AGEMA_signal_1643, new_AGEMA_signal_1642, new_AGEMA_signal_1641, TweakeyGeneration_key_Feedback[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_52__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1928, new_AGEMA_signal_1927, new_AGEMA_signal_1926, TweakeyGeneration_StateRegInput[52]}), .Q ({new_AGEMA_signal_1634, new_AGEMA_signal_1633, new_AGEMA_signal_1632, TweakeyGeneration_key_Feedback[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_51__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1919, new_AGEMA_signal_1918, new_AGEMA_signal_1917, TweakeyGeneration_StateRegInput[51]}), .Q ({new_AGEMA_signal_1625, new_AGEMA_signal_1624, new_AGEMA_signal_1623, TweakeyGeneration_key_Feedback[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_50__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1910, new_AGEMA_signal_1909, new_AGEMA_signal_1908, TweakeyGeneration_StateRegInput[50]}), .Q ({new_AGEMA_signal_1616, new_AGEMA_signal_1615, new_AGEMA_signal_1614, TweakeyGeneration_key_Feedback[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_49__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1901, new_AGEMA_signal_1900, new_AGEMA_signal_1899, TweakeyGeneration_StateRegInput[49]}), .Q ({new_AGEMA_signal_1607, new_AGEMA_signal_1606, new_AGEMA_signal_1605, TweakeyGeneration_key_Feedback[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_48__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1892, new_AGEMA_signal_1891, new_AGEMA_signal_1890, TweakeyGeneration_StateRegInput[48]}), .Q ({new_AGEMA_signal_1598, new_AGEMA_signal_1597, new_AGEMA_signal_1596, TweakeyGeneration_key_Feedback[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_47__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1883, new_AGEMA_signal_1882, new_AGEMA_signal_1881, TweakeyGeneration_StateRegInput[47]}), .Q ({new_AGEMA_signal_1589, new_AGEMA_signal_1588, new_AGEMA_signal_1587, TweakeyGeneration_key_Feedback[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_46__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1874, new_AGEMA_signal_1873, new_AGEMA_signal_1872, TweakeyGeneration_StateRegInput[46]}), .Q ({new_AGEMA_signal_1580, new_AGEMA_signal_1579, new_AGEMA_signal_1578, TweakeyGeneration_key_Feedback[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_45__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1865, new_AGEMA_signal_1864, new_AGEMA_signal_1863, TweakeyGeneration_StateRegInput[45]}), .Q ({new_AGEMA_signal_1571, new_AGEMA_signal_1570, new_AGEMA_signal_1569, TweakeyGeneration_key_Feedback[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_44__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1856, new_AGEMA_signal_1855, new_AGEMA_signal_1854, TweakeyGeneration_StateRegInput[44]}), .Q ({new_AGEMA_signal_1562, new_AGEMA_signal_1561, new_AGEMA_signal_1560, TweakeyGeneration_key_Feedback[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_43__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1847, new_AGEMA_signal_1846, new_AGEMA_signal_1845, TweakeyGeneration_StateRegInput[43]}), .Q ({new_AGEMA_signal_1553, new_AGEMA_signal_1552, new_AGEMA_signal_1551, TweakeyGeneration_key_Feedback[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_42__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1838, new_AGEMA_signal_1837, new_AGEMA_signal_1836, TweakeyGeneration_StateRegInput[42]}), .Q ({new_AGEMA_signal_1544, new_AGEMA_signal_1543, new_AGEMA_signal_1542, TweakeyGeneration_key_Feedback[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_41__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1829, new_AGEMA_signal_1828, new_AGEMA_signal_1827, TweakeyGeneration_StateRegInput[41]}), .Q ({new_AGEMA_signal_1535, new_AGEMA_signal_1534, new_AGEMA_signal_1533, TweakeyGeneration_key_Feedback[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_40__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1820, new_AGEMA_signal_1819, new_AGEMA_signal_1818, TweakeyGeneration_StateRegInput[40]}), .Q ({new_AGEMA_signal_1526, new_AGEMA_signal_1525, new_AGEMA_signal_1524, TweakeyGeneration_key_Feedback[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_39__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1811, new_AGEMA_signal_1810, new_AGEMA_signal_1809, TweakeyGeneration_StateRegInput[39]}), .Q ({new_AGEMA_signal_1517, new_AGEMA_signal_1516, new_AGEMA_signal_1515, TweakeyGeneration_key_Feedback[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_38__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1802, new_AGEMA_signal_1801, new_AGEMA_signal_1800, TweakeyGeneration_StateRegInput[38]}), .Q ({new_AGEMA_signal_1508, new_AGEMA_signal_1507, new_AGEMA_signal_1506, TweakeyGeneration_key_Feedback[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_37__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1793, new_AGEMA_signal_1792, new_AGEMA_signal_1791, TweakeyGeneration_StateRegInput[37]}), .Q ({new_AGEMA_signal_1499, new_AGEMA_signal_1498, new_AGEMA_signal_1497, TweakeyGeneration_key_Feedback[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_36__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1784, new_AGEMA_signal_1783, new_AGEMA_signal_1782, TweakeyGeneration_StateRegInput[36]}), .Q ({new_AGEMA_signal_1490, new_AGEMA_signal_1489, new_AGEMA_signal_1488, TweakeyGeneration_key_Feedback[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_35__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1775, new_AGEMA_signal_1774, new_AGEMA_signal_1773, TweakeyGeneration_StateRegInput[35]}), .Q ({new_AGEMA_signal_1481, new_AGEMA_signal_1480, new_AGEMA_signal_1479, TweakeyGeneration_key_Feedback[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_34__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1766, new_AGEMA_signal_1765, new_AGEMA_signal_1764, TweakeyGeneration_StateRegInput[34]}), .Q ({new_AGEMA_signal_1472, new_AGEMA_signal_1471, new_AGEMA_signal_1470, TweakeyGeneration_key_Feedback[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_33__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1757, new_AGEMA_signal_1756, new_AGEMA_signal_1755, TweakeyGeneration_StateRegInput[33]}), .Q ({new_AGEMA_signal_1463, new_AGEMA_signal_1462, new_AGEMA_signal_1461, TweakeyGeneration_key_Feedback[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_32__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1748, new_AGEMA_signal_1747, new_AGEMA_signal_1746, TweakeyGeneration_StateRegInput[32]}), .Q ({new_AGEMA_signal_1454, new_AGEMA_signal_1453, new_AGEMA_signal_1452, TweakeyGeneration_key_Feedback[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_31__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1739, new_AGEMA_signal_1738, new_AGEMA_signal_1737, TweakeyGeneration_StateRegInput[31]}), .Q ({new_AGEMA_signal_1949, new_AGEMA_signal_1948, new_AGEMA_signal_1947, TweakeyGeneration_key_Feedback[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_30__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1730, new_AGEMA_signal_1729, new_AGEMA_signal_1728, TweakeyGeneration_StateRegInput[30]}), .Q ({new_AGEMA_signal_1940, new_AGEMA_signal_1939, new_AGEMA_signal_1938, TweakeyGeneration_key_Feedback[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_29__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1721, new_AGEMA_signal_1720, new_AGEMA_signal_1719, TweakeyGeneration_StateRegInput[29]}), .Q ({new_AGEMA_signal_1931, new_AGEMA_signal_1930, new_AGEMA_signal_1929, TweakeyGeneration_key_Feedback[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_28__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1712, new_AGEMA_signal_1711, new_AGEMA_signal_1710, TweakeyGeneration_StateRegInput[28]}), .Q ({new_AGEMA_signal_1922, new_AGEMA_signal_1921, new_AGEMA_signal_1920, TweakeyGeneration_key_Feedback[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_27__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1703, new_AGEMA_signal_1702, new_AGEMA_signal_1701, TweakeyGeneration_StateRegInput[27]}), .Q ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, new_AGEMA_signal_2019, TweakeyGeneration_key_Feedback[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_26__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1694, new_AGEMA_signal_1693, new_AGEMA_signal_1692, TweakeyGeneration_StateRegInput[26]}), .Q ({new_AGEMA_signal_2012, new_AGEMA_signal_2011, new_AGEMA_signal_2010, TweakeyGeneration_key_Feedback[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_25__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1685, new_AGEMA_signal_1684, new_AGEMA_signal_1683, TweakeyGeneration_StateRegInput[25]}), .Q ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, new_AGEMA_signal_2001, TweakeyGeneration_key_Feedback[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_24__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1676, new_AGEMA_signal_1675, new_AGEMA_signal_1674, TweakeyGeneration_StateRegInput[24]}), .Q ({new_AGEMA_signal_1994, new_AGEMA_signal_1993, new_AGEMA_signal_1992, TweakeyGeneration_key_Feedback[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_23__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1667, new_AGEMA_signal_1666, new_AGEMA_signal_1665, TweakeyGeneration_StateRegInput[23]}), .Q ({new_AGEMA_signal_1877, new_AGEMA_signal_1876, new_AGEMA_signal_1875, TweakeyGeneration_key_Feedback[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_22__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1658, new_AGEMA_signal_1657, new_AGEMA_signal_1656, TweakeyGeneration_StateRegInput[22]}), .Q ({new_AGEMA_signal_1868, new_AGEMA_signal_1867, new_AGEMA_signal_1866, TweakeyGeneration_key_Feedback[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_21__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1649, new_AGEMA_signal_1648, new_AGEMA_signal_1647, TweakeyGeneration_StateRegInput[21]}), .Q ({new_AGEMA_signal_1859, new_AGEMA_signal_1858, new_AGEMA_signal_1857, TweakeyGeneration_key_Feedback[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_20__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1640, new_AGEMA_signal_1639, new_AGEMA_signal_1638, TweakeyGeneration_StateRegInput[20]}), .Q ({new_AGEMA_signal_1850, new_AGEMA_signal_1849, new_AGEMA_signal_1848, TweakeyGeneration_key_Feedback[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_19__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1631, new_AGEMA_signal_1630, new_AGEMA_signal_1629, TweakeyGeneration_StateRegInput[19]}), .Q ({new_AGEMA_signal_1769, new_AGEMA_signal_1768, new_AGEMA_signal_1767, TweakeyGeneration_key_Feedback[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_18__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1622, new_AGEMA_signal_1621, new_AGEMA_signal_1620, TweakeyGeneration_StateRegInput[18]}), .Q ({new_AGEMA_signal_1760, new_AGEMA_signal_1759, new_AGEMA_signal_1758, TweakeyGeneration_key_Feedback[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_17__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1613, new_AGEMA_signal_1612, new_AGEMA_signal_1611, TweakeyGeneration_StateRegInput[17]}), .Q ({new_AGEMA_signal_1751, new_AGEMA_signal_1750, new_AGEMA_signal_1749, TweakeyGeneration_key_Feedback[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_16__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1604, new_AGEMA_signal_1603, new_AGEMA_signal_1602, TweakeyGeneration_StateRegInput[16]}), .Q ({new_AGEMA_signal_1742, new_AGEMA_signal_1741, new_AGEMA_signal_1740, TweakeyGeneration_key_Feedback[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_15__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1595, new_AGEMA_signal_1594, new_AGEMA_signal_1593, TweakeyGeneration_StateRegInput[15]}), .Q ({new_AGEMA_signal_1805, new_AGEMA_signal_1804, new_AGEMA_signal_1803, TweakeyGeneration_key_Feedback[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_14__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1586, new_AGEMA_signal_1585, new_AGEMA_signal_1584, TweakeyGeneration_StateRegInput[14]}), .Q ({new_AGEMA_signal_1796, new_AGEMA_signal_1795, new_AGEMA_signal_1794, TweakeyGeneration_key_Feedback[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_13__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1577, new_AGEMA_signal_1576, new_AGEMA_signal_1575, TweakeyGeneration_StateRegInput[13]}), .Q ({new_AGEMA_signal_1787, new_AGEMA_signal_1786, new_AGEMA_signal_1785, TweakeyGeneration_key_Feedback[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_12__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1568, new_AGEMA_signal_1567, new_AGEMA_signal_1566, TweakeyGeneration_StateRegInput[12]}), .Q ({new_AGEMA_signal_1778, new_AGEMA_signal_1777, new_AGEMA_signal_1776, TweakeyGeneration_key_Feedback[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_11__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1559, new_AGEMA_signal_1558, new_AGEMA_signal_1557, TweakeyGeneration_StateRegInput[11]}), .Q ({new_AGEMA_signal_1913, new_AGEMA_signal_1912, new_AGEMA_signal_1911, TweakeyGeneration_key_Feedback[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_10__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1550, new_AGEMA_signal_1549, new_AGEMA_signal_1548, TweakeyGeneration_StateRegInput[10]}), .Q ({new_AGEMA_signal_1904, new_AGEMA_signal_1903, new_AGEMA_signal_1902, TweakeyGeneration_key_Feedback[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_9__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1541, new_AGEMA_signal_1540, new_AGEMA_signal_1539, TweakeyGeneration_StateRegInput[9]}), .Q ({new_AGEMA_signal_1895, new_AGEMA_signal_1894, new_AGEMA_signal_1893, TweakeyGeneration_key_Feedback[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_8__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1532, new_AGEMA_signal_1531, new_AGEMA_signal_1530, TweakeyGeneration_StateRegInput[8]}), .Q ({new_AGEMA_signal_1886, new_AGEMA_signal_1885, new_AGEMA_signal_1884, TweakeyGeneration_key_Feedback[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_7__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1523, new_AGEMA_signal_1522, new_AGEMA_signal_1521, TweakeyGeneration_StateRegInput[7]}), .Q ({new_AGEMA_signal_1841, new_AGEMA_signal_1840, new_AGEMA_signal_1839, TweakeyGeneration_key_Feedback[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_6__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1514, new_AGEMA_signal_1513, new_AGEMA_signal_1512, TweakeyGeneration_StateRegInput[6]}), .Q ({new_AGEMA_signal_1832, new_AGEMA_signal_1831, new_AGEMA_signal_1830, TweakeyGeneration_key_Feedback[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_5__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1505, new_AGEMA_signal_1504, new_AGEMA_signal_1503, TweakeyGeneration_StateRegInput[5]}), .Q ({new_AGEMA_signal_1823, new_AGEMA_signal_1822, new_AGEMA_signal_1821, TweakeyGeneration_key_Feedback[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_4__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1496, new_AGEMA_signal_1495, new_AGEMA_signal_1494, TweakeyGeneration_StateRegInput[4]}), .Q ({new_AGEMA_signal_1814, new_AGEMA_signal_1813, new_AGEMA_signal_1812, TweakeyGeneration_key_Feedback[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_3__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1487, new_AGEMA_signal_1486, new_AGEMA_signal_1485, TweakeyGeneration_StateRegInput[3]}), .Q ({new_AGEMA_signal_1985, new_AGEMA_signal_1984, new_AGEMA_signal_1983, TweakeyGeneration_key_Feedback[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_2__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1478, new_AGEMA_signal_1477, new_AGEMA_signal_1476, TweakeyGeneration_StateRegInput[2]}), .Q ({new_AGEMA_signal_1976, new_AGEMA_signal_1975, new_AGEMA_signal_1974, TweakeyGeneration_key_Feedback[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_1__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1469, new_AGEMA_signal_1468, new_AGEMA_signal_1467, TweakeyGeneration_StateRegInput[1]}), .Q ({new_AGEMA_signal_1967, new_AGEMA_signal_1966, new_AGEMA_signal_1965, TweakeyGeneration_key_Feedback[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) TweakeyGeneration_StateReg_s_current_state_reg_0__FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_1460, new_AGEMA_signal_1459, new_AGEMA_signal_1458, TweakeyGeneration_StateRegInput[0]}), .Q ({new_AGEMA_signal_1958, new_AGEMA_signal_1957, new_AGEMA_signal_1956, TweakeyGeneration_key_Feedback[56]}) ) ;
    DFF_X1 FSMReg_s_current_state_reg_5__FF_FF ( .CK (clk_gated), .D (FSMSelected[5]), .Q (FSM[5]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_4__FF_FF ( .CK (clk_gated), .D (FSMSelected[4]), .Q (FSM[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_3__FF_FF ( .CK (clk_gated), .D (FSMSelected[3]), .Q (FSMUpdate[4]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_2__FF_FF ( .CK (clk_gated), .D (FSMSelected[2]), .Q (FSMUpdate[3]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_1__FF_FF ( .CK (clk_gated), .D (FSMSelected[1]), .Q (FSM[1]), .QN () ) ;
    DFF_X1 FSMReg_s_current_state_reg_0__FF_FF ( .CK (clk_gated), .D (FSMSelected[0]), .Q (FSMUpdate[1]), .QN () ) ;
endmodule
